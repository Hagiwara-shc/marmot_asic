magic
tech sky130A
magscale 1 2
timestamp 1653258511
<< metal1 >>
rect 300118 700680 300124 700732
rect 300176 700720 300182 700732
rect 356698 700720 356704 700732
rect 300176 700692 356704 700720
rect 300176 700680 300182 700692
rect 356698 700680 356704 700692
rect 356756 700680 356762 700732
rect 283834 700612 283840 700664
rect 283892 700652 283898 700664
rect 344278 700652 344284 700664
rect 283892 700624 344284 700652
rect 283892 700612 283898 700624
rect 344278 700612 344284 700624
rect 344336 700612 344342 700664
rect 348786 700612 348792 700664
rect 348844 700652 348850 700664
rect 396718 700652 396724 700664
rect 348844 700624 396724 700652
rect 348844 700612 348850 700624
rect 396718 700612 396724 700624
rect 396776 700612 396782 700664
rect 332502 700544 332508 700596
rect 332560 700584 332566 700596
rect 404998 700584 405004 700596
rect 332560 700556 405004 700584
rect 332560 700544 332566 700556
rect 404998 700544 405004 700556
rect 405056 700544 405062 700596
rect 170306 700476 170312 700528
rect 170364 700516 170370 700528
rect 177298 700516 177304 700528
rect 170364 700488 177304 700516
rect 170364 700476 170370 700488
rect 177298 700476 177304 700488
rect 177356 700476 177362 700528
rect 267642 700476 267648 700528
rect 267700 700516 267706 700528
rect 351178 700516 351184 700528
rect 267700 700488 351184 700516
rect 267700 700476 267706 700488
rect 351178 700476 351184 700488
rect 351236 700476 351242 700528
rect 137830 700408 137836 700460
rect 137888 700448 137894 700460
rect 184198 700448 184204 700460
rect 137888 700420 184204 700448
rect 137888 700408 137894 700420
rect 184198 700408 184204 700420
rect 184256 700408 184262 700460
rect 235166 700408 235172 700460
rect 235224 700448 235230 700460
rect 358078 700448 358084 700460
rect 235224 700420 358084 700448
rect 235224 700408 235230 700420
rect 358078 700408 358084 700420
rect 358136 700408 358142 700460
rect 408402 700408 408408 700460
rect 408460 700448 408466 700460
rect 429838 700448 429844 700460
rect 408460 700420 429844 700448
rect 408460 700408 408466 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 72970 700340 72976 700392
rect 73028 700380 73034 700392
rect 186958 700380 186964 700392
rect 73028 700352 186964 700380
rect 73028 700340 73034 700352
rect 186958 700340 186964 700352
rect 187016 700340 187022 700392
rect 218974 700340 218980 700392
rect 219032 700380 219038 700392
rect 348418 700380 348424 700392
rect 219032 700352 348424 700380
rect 219032 700340 219038 700352
rect 348418 700340 348424 700352
rect 348476 700340 348482 700392
rect 409782 700340 409788 700392
rect 409840 700380 409846 700392
rect 462314 700380 462320 700392
rect 409840 700352 462320 700380
rect 409840 700340 409846 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 527174 700340 527180 700392
rect 527232 700380 527238 700392
rect 546678 700380 546684 700392
rect 527232 700352 546684 700380
rect 527232 700340 527238 700352
rect 546678 700340 546684 700352
rect 546736 700340 546742 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 188338 700312 188344 700324
rect 8168 700284 188344 700312
rect 8168 700272 8174 700284
rect 188338 700272 188344 700284
rect 188396 700272 188402 700324
rect 202782 700272 202788 700324
rect 202840 700312 202846 700324
rect 353938 700312 353944 700324
rect 202840 700284 353944 700312
rect 202840 700272 202846 700284
rect 353938 700272 353944 700284
rect 353996 700272 354002 700324
rect 364978 700272 364984 700324
rect 365036 700312 365042 700324
rect 393958 700312 393964 700324
rect 365036 700284 393964 700312
rect 365036 700272 365042 700284
rect 393958 700272 393964 700284
rect 394016 700272 394022 700324
rect 408310 700272 408316 700324
rect 408368 700312 408374 700324
rect 478506 700312 478512 700324
rect 408368 700284 478512 700312
rect 408368 700272 408374 700284
rect 478506 700272 478512 700284
rect 478564 700272 478570 700324
rect 494790 700272 494796 700324
rect 494848 700312 494854 700324
rect 546770 700312 546776 700324
rect 494848 700284 546776 700312
rect 494848 700272 494854 700284
rect 546770 700272 546776 700284
rect 546828 700272 546834 700324
rect 548518 700272 548524 700324
rect 548576 700312 548582 700324
rect 559650 700312 559656 700324
rect 548576 700284 559656 700312
rect 548576 700272 548582 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 409690 699660 409696 699712
rect 409748 699700 409754 699712
rect 413646 699700 413652 699712
rect 409748 699672 413652 699700
rect 409748 699660 409754 699672
rect 413646 699660 413652 699672
rect 413704 699660 413710 699712
rect 543458 699660 543464 699712
rect 543516 699700 543522 699712
rect 547874 699700 547880 699712
rect 543516 699672 547880 699700
rect 543516 699660 543522 699672
rect 547874 699660 547880 699672
rect 547932 699660 547938 699712
rect 105446 698912 105452 698964
rect 105504 698952 105510 698964
rect 407758 698952 407764 698964
rect 105504 698924 407764 698952
rect 105504 698912 105510 698924
rect 407758 698912 407764 698924
rect 407816 698912 407822 698964
rect 577498 696940 577504 696992
rect 577556 696980 577562 696992
rect 580442 696980 580448 696992
rect 577556 696952 580448 696980
rect 577556 696940 577562 696952
rect 580442 696940 580448 696952
rect 580500 696940 580506 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 178770 683176 178776 683188
rect 3476 683148 178776 683176
rect 3476 683136 3482 683148
rect 178770 683136 178776 683148
rect 178828 683136 178834 683188
rect 28718 674976 28724 675028
rect 28776 675016 28782 675028
rect 28776 674988 35894 675016
rect 28776 674976 28782 674988
rect 28626 674908 28632 674960
rect 28684 674948 28690 674960
rect 34514 674948 34520 674960
rect 28684 674920 34520 674948
rect 28684 674908 28690 674920
rect 34514 674908 34520 674920
rect 34572 674908 34578 674960
rect 35866 674948 35894 674988
rect 46198 674948 46204 674960
rect 35866 674920 46204 674948
rect 46198 674908 46204 674920
rect 46256 674908 46262 674960
rect 28810 674840 28816 674892
rect 28868 674880 28874 674892
rect 46934 674880 46940 674892
rect 28868 674852 46940 674880
rect 28868 674840 28874 674852
rect 46934 674840 46940 674852
rect 46992 674840 46998 674892
rect 570598 670692 570604 670744
rect 570656 670732 570662 670744
rect 580166 670732 580172 670744
rect 570656 670704 580172 670732
rect 570656 670692 570662 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 340138 660288 340144 660340
rect 340196 660328 340202 660340
rect 488902 660328 488908 660340
rect 340196 660300 488908 660328
rect 340196 660288 340202 660300
rect 488902 660288 488908 660300
rect 488960 660288 488966 660340
rect 246298 659676 246304 659728
rect 246356 659716 246362 659728
rect 337102 659716 337108 659728
rect 246356 659688 337108 659716
rect 246356 659676 246362 659688
rect 337102 659676 337108 659688
rect 337160 659676 337166 659728
rect 408218 659676 408224 659728
rect 408276 659716 408282 659728
rect 499850 659716 499856 659728
rect 408276 659688 499856 659716
rect 408276 659676 408282 659688
rect 499850 659676 499856 659688
rect 499908 659676 499914 659728
rect 560938 643084 560944 643136
rect 560996 643124 561002 643136
rect 580166 643124 580172 643136
rect 560996 643096 580172 643124
rect 560996 643084 561002 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2958 618264 2964 618316
rect 3016 618304 3022 618316
rect 21358 618304 21364 618316
rect 3016 618276 21364 618304
rect 3016 618264 3022 618276
rect 21358 618264 21364 618276
rect 21416 618264 21422 618316
rect 567838 616836 567844 616888
rect 567896 616876 567902 616888
rect 580166 616876 580172 616888
rect 567896 616848 580172 616876
rect 567896 616836 567902 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 339402 612008 339408 612060
rect 339460 612048 339466 612060
rect 407114 612048 407120 612060
rect 339460 612020 407120 612048
rect 339460 612008 339466 612020
rect 407114 612008 407120 612020
rect 407172 612008 407178 612060
rect 339402 610580 339408 610632
rect 339460 610620 339466 610632
rect 407114 610620 407120 610632
rect 339460 610592 407120 610620
rect 339460 610580 339466 610592
rect 407114 610580 407120 610592
rect 407172 610580 407178 610632
rect 338298 608608 338304 608660
rect 338356 608648 338362 608660
rect 407114 608648 407120 608660
rect 338356 608620 407120 608648
rect 338356 608608 338362 608620
rect 407114 608608 407120 608620
rect 407172 608608 407178 608660
rect 338114 607180 338120 607232
rect 338172 607220 338178 607232
rect 407114 607220 407120 607232
rect 338172 607192 407120 607220
rect 338172 607180 338178 607192
rect 407114 607180 407120 607192
rect 407172 607180 407178 607232
rect 338390 605820 338396 605872
rect 338448 605860 338454 605872
rect 407114 605860 407120 605872
rect 338448 605832 407120 605860
rect 338448 605820 338454 605832
rect 407114 605820 407120 605832
rect 407172 605820 407178 605872
rect 338206 604460 338212 604512
rect 338264 604500 338270 604512
rect 339402 604500 339408 604512
rect 338264 604472 339408 604500
rect 338264 604460 338270 604472
rect 339402 604460 339408 604472
rect 339460 604500 339466 604512
rect 407114 604500 407120 604512
rect 339460 604472 407120 604500
rect 339460 604460 339466 604472
rect 407114 604460 407120 604472
rect 407172 604460 407178 604512
rect 339218 603712 339224 603764
rect 339276 603752 339282 603764
rect 407114 603752 407120 603764
rect 339276 603724 407120 603752
rect 339276 603712 339282 603724
rect 407114 603712 407120 603724
rect 407172 603712 407178 603764
rect 574738 590656 574744 590708
rect 574796 590696 574802 590708
rect 580166 590696 580172 590708
rect 574796 590668 580172 590696
rect 574796 590656 574802 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 99190 587392 99196 587444
rect 99248 587432 99254 587444
rect 170858 587432 170864 587444
rect 99248 587404 170864 587432
rect 99248 587392 99254 587404
rect 170858 587392 170864 587404
rect 170916 587392 170922 587444
rect 149514 587324 149520 587376
rect 149572 587364 149578 587376
rect 171594 587364 171600 587376
rect 149572 587336 171600 587364
rect 149572 587324 149578 587336
rect 171594 587324 171600 587336
rect 171652 587324 171658 587376
rect 143442 587256 143448 587308
rect 143500 587296 143506 587308
rect 166994 587296 167000 587308
rect 143500 587268 167000 587296
rect 143500 587256 143506 587268
rect 166994 587256 167000 587268
rect 167052 587256 167058 587308
rect 142706 587188 142712 587240
rect 142764 587228 142770 587240
rect 168098 587228 168104 587240
rect 142764 587200 168104 587228
rect 142764 587188 142770 587200
rect 168098 587188 168104 587200
rect 168156 587188 168162 587240
rect 140130 587120 140136 587172
rect 140188 587160 140194 587172
rect 168006 587160 168012 587172
rect 140188 587132 168012 587160
rect 140188 587120 140194 587132
rect 168006 587120 168012 587132
rect 168064 587120 168070 587172
rect 137922 587052 137928 587104
rect 137980 587092 137986 587104
rect 167822 587092 167828 587104
rect 137980 587064 167828 587092
rect 137980 587052 137986 587064
rect 167822 587052 167828 587064
rect 167880 587052 167886 587104
rect 139026 586984 139032 587036
rect 139084 587024 139090 587036
rect 171410 587024 171416 587036
rect 139084 586996 171416 587024
rect 139084 586984 139090 586996
rect 171410 586984 171416 586996
rect 171468 586984 171474 587036
rect 136542 586916 136548 586968
rect 136600 586956 136606 586968
rect 169754 586956 169760 586968
rect 136600 586928 169760 586956
rect 136600 586916 136606 586928
rect 169754 586916 169760 586928
rect 169812 586916 169818 586968
rect 133138 586848 133144 586900
rect 133196 586888 133202 586900
rect 167914 586888 167920 586900
rect 133196 586860 167920 586888
rect 133196 586848 133202 586860
rect 167914 586848 167920 586860
rect 167972 586848 167978 586900
rect 129642 586780 129648 586832
rect 129700 586820 129706 586832
rect 172790 586820 172796 586832
rect 129700 586792 172796 586820
rect 129700 586780 129706 586792
rect 172790 586780 172796 586792
rect 172848 586780 172854 586832
rect 126882 586712 126888 586764
rect 126940 586752 126946 586764
rect 173526 586752 173532 586764
rect 126940 586724 173532 586752
rect 126940 586712 126946 586724
rect 173526 586712 173532 586724
rect 173584 586712 173590 586764
rect 100570 586644 100576 586696
rect 100628 586684 100634 586696
rect 170766 586684 170772 586696
rect 100628 586656 170772 586684
rect 100628 586644 100634 586656
rect 170766 586644 170772 586656
rect 170824 586644 170830 586696
rect 28534 586576 28540 586628
rect 28592 586616 28598 586628
rect 43070 586616 43076 586628
rect 28592 586588 43076 586616
rect 28592 586576 28598 586588
rect 43070 586576 43076 586588
rect 43128 586576 43134 586628
rect 103146 586576 103152 586628
rect 103204 586616 103210 586628
rect 174630 586616 174636 586628
rect 103204 586588 174636 586616
rect 103204 586576 103210 586588
rect 174630 586576 174636 586588
rect 174688 586576 174694 586628
rect 28442 586508 28448 586560
rect 28500 586548 28506 586560
rect 43530 586548 43536 586560
rect 28500 586520 43536 586548
rect 28500 586508 28506 586520
rect 43530 586508 43536 586520
rect 43588 586508 43594 586560
rect 150710 586508 150716 586560
rect 150768 586548 150774 586560
rect 167086 586548 167092 586560
rect 150768 586520 167092 586548
rect 150768 586508 150774 586520
rect 167086 586508 167092 586520
rect 167144 586508 167150 586560
rect 139302 585828 139308 585880
rect 139360 585868 139366 585880
rect 181530 585868 181536 585880
rect 139360 585840 181536 585868
rect 139360 585828 139366 585840
rect 181530 585828 181536 585840
rect 181588 585828 181594 585880
rect 105078 585760 105084 585812
rect 105136 585800 105142 585812
rect 174722 585800 174728 585812
rect 105136 585772 174728 585800
rect 105136 585760 105142 585772
rect 174722 585760 174728 585772
rect 174780 585760 174786 585812
rect 339218 585760 339224 585812
rect 339276 585800 339282 585812
rect 407114 585800 407120 585812
rect 339276 585772 407120 585800
rect 339276 585760 339282 585772
rect 407114 585760 407120 585772
rect 407172 585760 407178 585812
rect 130562 585080 130568 585132
rect 130620 585120 130626 585132
rect 172882 585120 172888 585132
rect 130620 585092 172888 585120
rect 130620 585080 130626 585092
rect 172882 585080 172888 585092
rect 172940 585080 172946 585132
rect 120534 585012 120540 585064
rect 120592 585052 120598 585064
rect 167178 585052 167184 585064
rect 120592 585024 167184 585052
rect 120592 585012 120598 585024
rect 167178 585012 167184 585024
rect 167236 585012 167242 585064
rect 125042 584944 125048 584996
rect 125100 584984 125106 584996
rect 175366 584984 175372 584996
rect 125100 584956 175372 584984
rect 125100 584944 125106 584956
rect 175366 584944 175372 584956
rect 175424 584944 175430 584996
rect 129366 584876 129372 584928
rect 129424 584916 129430 584928
rect 180794 584916 180800 584928
rect 129424 584888 180800 584916
rect 129424 584876 129430 584888
rect 180794 584876 180800 584888
rect 180852 584876 180858 584928
rect 122650 584808 122656 584860
rect 122708 584848 122714 584860
rect 178034 584848 178040 584860
rect 122708 584820 178040 584848
rect 122708 584808 122714 584820
rect 178034 584808 178040 584820
rect 178092 584808 178098 584860
rect 117130 584740 117136 584792
rect 117188 584780 117194 584792
rect 172514 584780 172520 584792
rect 117188 584752 172520 584780
rect 117188 584740 117194 584752
rect 172514 584740 172520 584752
rect 172572 584740 172578 584792
rect 114830 584672 114836 584724
rect 114888 584712 114894 584724
rect 171226 584712 171232 584724
rect 114888 584684 171232 584712
rect 114888 584672 114894 584684
rect 171226 584672 171232 584684
rect 171284 584672 171290 584724
rect 113818 584604 113824 584656
rect 113876 584644 113882 584656
rect 172606 584644 172612 584656
rect 113876 584616 172612 584644
rect 113876 584604 113882 584616
rect 172606 584604 172612 584616
rect 172664 584604 172670 584656
rect 109494 584536 109500 584588
rect 109552 584576 109558 584588
rect 171318 584576 171324 584588
rect 109552 584548 171324 584576
rect 109552 584536 109558 584548
rect 171318 584536 171324 584548
rect 171376 584536 171382 584588
rect 110506 584468 110512 584520
rect 110564 584508 110570 584520
rect 187142 584508 187148 584520
rect 110564 584480 187148 584508
rect 110564 584468 110570 584480
rect 187142 584468 187148 584480
rect 187200 584468 187206 584520
rect 62942 584400 62948 584452
rect 63000 584440 63006 584452
rect 196894 584440 196900 584452
rect 63000 584412 196900 584440
rect 63000 584400 63006 584412
rect 196894 584400 196900 584412
rect 196952 584400 196958 584452
rect 131114 584332 131120 584384
rect 131172 584372 131178 584384
rect 173250 584372 173256 584384
rect 131172 584344 173256 584372
rect 131172 584332 131178 584344
rect 173250 584332 173256 584344
rect 173308 584332 173314 584384
rect 136450 584264 136456 584316
rect 136508 584304 136514 584316
rect 167638 584304 167644 584316
rect 136508 584276 167644 584304
rect 136508 584264 136514 584276
rect 167638 584264 167644 584276
rect 167696 584264 167702 584316
rect 147674 584196 147680 584248
rect 147732 584236 147738 584248
rect 171502 584236 171508 584248
rect 147732 584208 171508 584236
rect 147732 584196 147738 584208
rect 171502 584196 171508 584208
rect 171560 584196 171566 584248
rect 132586 582972 132592 583024
rect 132644 583012 132650 583024
rect 178954 583012 178960 583024
rect 132644 582984 178960 583012
rect 132644 582972 132650 582984
rect 178954 582972 178960 582984
rect 179012 582972 179018 583024
rect 339402 582972 339408 583024
rect 339460 583012 339466 583024
rect 407114 583012 407120 583024
rect 339460 582984 407120 583012
rect 339460 582972 339466 582984
rect 407114 582972 407120 582984
rect 407172 582972 407178 583024
rect 122834 581680 122840 581732
rect 122892 581720 122898 581732
rect 180058 581720 180064 581732
rect 122892 581692 180064 581720
rect 122892 581680 122898 581692
rect 180058 581680 180064 581692
rect 180116 581680 180122 581732
rect 95234 581612 95240 581664
rect 95292 581652 95298 581664
rect 185670 581652 185676 581664
rect 95292 581624 185676 581652
rect 95292 581612 95298 581624
rect 185670 581612 185676 581624
rect 185728 581612 185734 581664
rect 64874 580252 64880 580304
rect 64932 580292 64938 580304
rect 189810 580292 189816 580304
rect 64932 580264 189816 580292
rect 64932 580252 64938 580264
rect 189810 580252 189816 580264
rect 189868 580252 189874 580304
rect 3142 579640 3148 579692
rect 3200 579680 3206 579692
rect 181438 579680 181444 579692
rect 3200 579652 181444 579680
rect 3200 579640 3206 579652
rect 181438 579640 181444 579652
rect 181496 579640 181502 579692
rect 120166 578960 120172 579012
rect 120224 579000 120230 579012
rect 191190 579000 191196 579012
rect 120224 578972 191196 579000
rect 120224 578960 120230 578972
rect 191190 578960 191196 578972
rect 191248 578960 191254 579012
rect 83826 578892 83832 578944
rect 83884 578932 83890 578944
rect 194042 578932 194048 578944
rect 83884 578904 194048 578932
rect 83884 578892 83890 578904
rect 194042 578892 194048 578904
rect 194100 578892 194106 578944
rect 114554 577532 114560 577584
rect 114612 577572 114618 577584
rect 184290 577572 184296 577584
rect 114612 577544 184296 577572
rect 114612 577532 114618 577544
rect 184290 577532 184296 577544
rect 184348 577532 184354 577584
rect 86402 577464 86408 577516
rect 86460 577504 86466 577516
rect 195422 577504 195428 577516
rect 86460 577476 195428 577504
rect 86460 577464 86466 577476
rect 195422 577464 195428 577476
rect 195480 577464 195486 577516
rect 565078 576852 565084 576904
rect 565136 576892 565142 576904
rect 580166 576892 580172 576904
rect 565136 576864 580172 576892
rect 565136 576852 565142 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 113082 576172 113088 576224
rect 113140 576212 113146 576224
rect 177482 576212 177488 576224
rect 113140 576184 177488 576212
rect 113140 576172 113146 576184
rect 177482 576172 177488 576184
rect 177540 576172 177546 576224
rect 93762 576104 93768 576156
rect 93820 576144 93826 576156
rect 196802 576144 196808 576156
rect 93820 576116 196808 576144
rect 93820 576104 93826 576116
rect 196802 576104 196808 576116
rect 196860 576104 196866 576156
rect 338022 575492 338028 575544
rect 338080 575532 338086 575544
rect 425054 575532 425060 575544
rect 338080 575504 425060 575532
rect 338080 575492 338086 575504
rect 425054 575492 425060 575504
rect 425112 575492 425118 575544
rect 330202 575424 330208 575476
rect 330260 575464 330266 575476
rect 337102 575464 337108 575476
rect 330260 575436 337108 575464
rect 330260 575424 330266 575436
rect 337102 575424 337108 575436
rect 337160 575464 337166 575476
rect 408218 575464 408224 575476
rect 337160 575436 408224 575464
rect 337160 575424 337166 575436
rect 408218 575424 408224 575436
rect 408276 575464 408282 575476
rect 415394 575464 415400 575476
rect 408276 575436 415400 575464
rect 408276 575424 408282 575436
rect 415394 575424 415400 575436
rect 415452 575424 415458 575476
rect 199378 575152 199384 575204
rect 199436 575192 199442 575204
rect 293954 575192 293960 575204
rect 199436 575164 293960 575192
rect 199436 575152 199442 575164
rect 293954 575152 293960 575164
rect 294012 575152 294018 575204
rect 195698 575084 195704 575136
rect 195756 575124 195762 575136
rect 289814 575124 289820 575136
rect 195756 575096 289820 575124
rect 195756 575084 195762 575096
rect 289814 575084 289820 575096
rect 289872 575084 289878 575136
rect 198642 575016 198648 575068
rect 198700 575056 198706 575068
rect 293954 575056 293960 575068
rect 198700 575028 293960 575056
rect 198700 575016 198706 575028
rect 293954 575016 293960 575028
rect 294012 575016 294018 575068
rect 301866 575016 301872 575068
rect 301924 575056 301930 575068
rect 342346 575056 342352 575068
rect 301924 575028 342352 575056
rect 301924 575016 301930 575028
rect 342346 575016 342352 575028
rect 342404 575016 342410 575068
rect 199838 574948 199844 575000
rect 199896 574988 199902 575000
rect 280154 574988 280160 575000
rect 199896 574960 280160 574988
rect 199896 574948 199902 574960
rect 280154 574948 280160 574960
rect 280212 574948 280218 575000
rect 320450 574948 320456 575000
rect 320508 574988 320514 575000
rect 330478 574988 330484 575000
rect 320508 574960 330484 574988
rect 320508 574948 320514 574960
rect 330478 574948 330484 574960
rect 330536 574948 330542 575000
rect 340138 574948 340144 575000
rect 340196 574988 340202 575000
rect 466454 574988 466460 575000
rect 340196 574960 466460 574988
rect 340196 574948 340202 574960
rect 466454 574948 466460 574960
rect 466512 574948 466518 575000
rect 195882 574880 195888 574932
rect 195940 574920 195946 574932
rect 280246 574920 280252 574932
rect 195940 574892 280252 574920
rect 195940 574880 195946 574892
rect 280246 574880 280252 574892
rect 280304 574880 280310 574932
rect 307570 574880 307576 574932
rect 307628 574920 307634 574932
rect 339586 574920 339592 574932
rect 307628 574892 339592 574920
rect 307628 574880 307634 574892
rect 339586 574880 339592 574892
rect 339644 574880 339650 574932
rect 409414 574880 409420 574932
rect 409472 574920 409478 574932
rect 426434 574920 426440 574932
rect 409472 574892 426440 574920
rect 409472 574880 409478 574892
rect 426434 574880 426440 574892
rect 426492 574880 426498 574932
rect 118602 574812 118608 574864
rect 118660 574852 118666 574864
rect 188430 574852 188436 574864
rect 118660 574824 188436 574852
rect 118660 574812 118666 574824
rect 188430 574812 188436 574824
rect 188488 574812 188494 574864
rect 197078 574812 197084 574864
rect 197136 574852 197142 574864
rect 281534 574852 281540 574864
rect 197136 574824 281540 574852
rect 197136 574812 197142 574824
rect 281534 574812 281540 574824
rect 281592 574812 281598 574864
rect 304626 574812 304632 574864
rect 304684 574852 304690 574864
rect 336826 574852 336832 574864
rect 304684 574824 336832 574852
rect 304684 574812 304690 574824
rect 336826 574812 336832 574824
rect 336884 574812 336890 574864
rect 409506 574812 409512 574864
rect 409564 574852 409570 574864
rect 437474 574852 437480 574864
rect 409564 574824 437480 574852
rect 409564 574812 409570 574824
rect 437474 574812 437480 574824
rect 437532 574812 437538 574864
rect 81342 574744 81348 574796
rect 81400 574784 81406 574796
rect 191282 574784 191288 574796
rect 81400 574756 191288 574784
rect 81400 574744 81406 574756
rect 191282 574744 191288 574756
rect 191340 574744 191346 574796
rect 197170 574744 197176 574796
rect 197228 574784 197234 574796
rect 284294 574784 284300 574796
rect 197228 574756 284300 574784
rect 197228 574744 197234 574756
rect 284294 574744 284300 574756
rect 284352 574744 284358 574796
rect 305546 574744 305552 574796
rect 305604 574784 305610 574796
rect 339678 574784 339684 574796
rect 305604 574756 339684 574784
rect 305604 574744 305610 574756
rect 339678 574744 339684 574756
rect 339736 574744 339742 574796
rect 406562 574744 406568 574796
rect 406620 574784 406626 574796
rect 438854 574784 438860 574796
rect 406620 574756 438860 574784
rect 406620 574744 406626 574756
rect 438854 574744 438860 574756
rect 438912 574744 438918 574796
rect 195606 574676 195612 574728
rect 195664 574716 195670 574728
rect 284386 574716 284392 574728
rect 195664 574688 284392 574716
rect 195664 574676 195670 574688
rect 284386 574676 284392 574688
rect 284444 574676 284450 574728
rect 306282 574676 306288 574728
rect 306340 574716 306346 574728
rect 339770 574716 339776 574728
rect 306340 574688 339776 574716
rect 306340 574676 306346 574688
rect 339770 574676 339776 574688
rect 339828 574676 339834 574728
rect 406470 574676 406476 574728
rect 406528 574716 406534 574728
rect 444374 574716 444380 574728
rect 406528 574688 444380 574716
rect 406528 574676 406534 574688
rect 444374 574676 444380 574688
rect 444432 574676 444438 574728
rect 285306 574608 285312 574660
rect 285364 574648 285370 574660
rect 339954 574648 339960 574660
rect 285364 574620 339960 574648
rect 285364 574608 285370 574620
rect 339954 574608 339960 574620
rect 340012 574608 340018 574660
rect 409230 574608 409236 574660
rect 409288 574648 409294 574660
rect 451274 574648 451280 574660
rect 409288 574620 451280 574648
rect 409288 574608 409294 574620
rect 451274 574608 451280 574620
rect 451332 574608 451338 574660
rect 195790 574540 195796 574592
rect 195848 574580 195854 574592
rect 287514 574580 287520 574592
rect 195848 574552 287520 574580
rect 195848 574540 195854 574552
rect 287514 574540 287520 574552
rect 287572 574540 287578 574592
rect 302878 574540 302884 574592
rect 302936 574580 302942 574592
rect 337470 574580 337476 574592
rect 302936 574552 337476 574580
rect 302936 574540 302942 574552
rect 337470 574540 337476 574552
rect 337528 574540 337534 574592
rect 405274 574540 405280 574592
rect 405332 574580 405338 574592
rect 448514 574580 448520 574592
rect 405332 574552 448520 574580
rect 405332 574540 405338 574552
rect 448514 574540 448520 574552
rect 448572 574540 448578 574592
rect 287882 574472 287888 574524
rect 287940 574512 287946 574524
rect 341426 574512 341432 574524
rect 287940 574484 341432 574512
rect 287940 574472 287946 574484
rect 341426 574472 341432 574484
rect 341484 574472 341490 574524
rect 405090 574472 405096 574524
rect 405148 574512 405154 574524
rect 451274 574512 451280 574524
rect 405148 574484 451280 574512
rect 405148 574472 405154 574484
rect 451274 574472 451280 574484
rect 451332 574472 451338 574524
rect 490558 574472 490564 574524
rect 490616 574512 490622 574524
rect 492674 574512 492680 574524
rect 490616 574484 492680 574512
rect 490616 574472 490622 574484
rect 492674 574472 492680 574484
rect 492732 574472 492738 574524
rect 198550 574404 198556 574456
rect 198608 574444 198614 574456
rect 291194 574444 291200 574456
rect 198608 574416 291200 574444
rect 198608 574404 198614 574416
rect 291194 574404 291200 574416
rect 291252 574404 291258 574456
rect 300670 574404 300676 574456
rect 300728 574444 300734 574456
rect 342438 574444 342444 574456
rect 300728 574416 342444 574444
rect 300728 574404 300734 574416
rect 342438 574404 342444 574416
rect 342496 574404 342502 574456
rect 406378 574404 406384 574456
rect 406436 574444 406442 574456
rect 455414 574444 455420 574456
rect 406436 574416 455420 574444
rect 406436 574404 406442 574416
rect 455414 574404 455420 574416
rect 455472 574404 455478 574456
rect 199746 574336 199752 574388
rect 199804 574376 199810 574388
rect 292574 574376 292580 574388
rect 199804 574348 292580 574376
rect 199804 574336 199810 574348
rect 292574 574336 292580 574348
rect 292632 574336 292638 574388
rect 297910 574336 297916 574388
rect 297968 574376 297974 574388
rect 340966 574376 340972 574388
rect 297968 574348 340972 574376
rect 297968 574336 297974 574348
rect 340966 574336 340972 574348
rect 341024 574336 341030 574388
rect 400858 574336 400864 574388
rect 400916 574376 400922 574388
rect 458174 574376 458180 574388
rect 400916 574348 458180 574376
rect 400916 574336 400922 574348
rect 458174 574336 458180 574348
rect 458232 574336 458238 574388
rect 284202 574268 284208 574320
rect 284260 574308 284266 574320
rect 342254 574308 342260 574320
rect 284260 574280 342260 574308
rect 284260 574268 284266 574280
rect 342254 574268 342260 574280
rect 342312 574268 342318 574320
rect 398098 574268 398104 574320
rect 398156 574308 398162 574320
rect 462866 574308 462872 574320
rect 398156 574280 462872 574308
rect 398156 574268 398162 574280
rect 462866 574268 462872 574280
rect 462924 574268 462930 574320
rect 480898 574268 480904 574320
rect 480956 574308 480962 574320
rect 492674 574308 492680 574320
rect 480956 574280 492680 574308
rect 480956 574268 480962 574280
rect 492674 574268 492680 574280
rect 492732 574268 492738 574320
rect 196710 574200 196716 574252
rect 196768 574240 196774 574252
rect 288434 574240 288440 574252
rect 196768 574212 288440 574240
rect 196768 574200 196774 574212
rect 288434 574200 288440 574212
rect 288492 574200 288498 574252
rect 292482 574200 292488 574252
rect 292540 574240 292546 574252
rect 339494 574240 339500 574252
rect 292540 574212 339500 574240
rect 292540 574200 292546 574212
rect 339494 574200 339500 574212
rect 339552 574200 339558 574252
rect 396810 574200 396816 574252
rect 396868 574240 396874 574252
rect 465074 574240 465080 574252
rect 396868 574212 465080 574240
rect 396868 574200 396874 574212
rect 465074 574200 465080 574212
rect 465132 574200 465138 574252
rect 487798 574200 487804 574252
rect 487856 574240 487862 574252
rect 492766 574240 492772 574252
rect 487856 574212 492772 574240
rect 487856 574200 487862 574212
rect 492766 574200 492772 574212
rect 492824 574200 492830 574252
rect 196986 574132 196992 574184
rect 197044 574172 197050 574184
rect 285674 574172 285680 574184
rect 197044 574144 285680 574172
rect 197044 574132 197050 574144
rect 285674 574132 285680 574144
rect 285732 574132 285738 574184
rect 286594 574132 286600 574184
rect 286652 574172 286658 574184
rect 341518 574172 341524 574184
rect 286652 574144 341524 574172
rect 286652 574132 286658 574144
rect 341518 574132 341524 574144
rect 341576 574132 341582 574184
rect 391198 574132 391204 574184
rect 391256 574172 391262 574184
rect 459554 574172 459560 574184
rect 391256 574144 459560 574172
rect 391256 574132 391262 574144
rect 459554 574132 459560 574144
rect 459612 574132 459618 574184
rect 485038 574132 485044 574184
rect 485096 574172 485102 574184
rect 492950 574172 492956 574184
rect 485096 574144 492956 574172
rect 485096 574132 485102 574144
rect 492950 574132 492956 574144
rect 493008 574132 493014 574184
rect 195514 574064 195520 574116
rect 195572 574104 195578 574116
rect 306466 574104 306472 574116
rect 195572 574076 306472 574104
rect 195572 574064 195578 574076
rect 306466 574064 306472 574076
rect 306524 574064 306530 574116
rect 68922 573384 68928 573436
rect 68980 573424 68986 573436
rect 177574 573424 177580 573436
rect 68980 573396 177580 573424
rect 68980 573384 68986 573396
rect 177574 573384 177580 573396
rect 177632 573384 177638 573436
rect 191742 573384 191748 573436
rect 191800 573424 191806 573436
rect 269114 573424 269120 573436
rect 191800 573396 269120 573424
rect 191800 573384 191806 573396
rect 269114 573384 269120 573396
rect 269172 573384 269178 573436
rect 360194 573384 360200 573436
rect 360252 573424 360258 573436
rect 447134 573424 447140 573436
rect 360252 573396 447140 573424
rect 360252 573384 360258 573396
rect 447134 573384 447140 573396
rect 447192 573384 447198 573436
rect 3602 573316 3608 573368
rect 3660 573356 3666 573368
rect 407850 573356 407856 573368
rect 3660 573328 407856 573356
rect 3660 573316 3666 573328
rect 407850 573316 407856 573328
rect 407908 573316 407914 573368
rect 199562 572636 199568 572688
rect 199620 572676 199626 572688
rect 276014 572676 276020 572688
rect 199620 572648 276020 572676
rect 199620 572636 199626 572648
rect 276014 572636 276020 572648
rect 276072 572636 276078 572688
rect 291010 572636 291016 572688
rect 291068 572676 291074 572688
rect 337102 572676 337108 572688
rect 291068 572648 337108 572676
rect 291068 572636 291074 572648
rect 337102 572636 337108 572648
rect 337160 572636 337166 572688
rect 402238 572636 402244 572688
rect 402296 572676 402302 572688
rect 443086 572676 443092 572688
rect 402296 572648 443092 572676
rect 402296 572636 402302 572648
rect 443086 572636 443092 572648
rect 443144 572636 443150 572688
rect 198458 572568 198464 572620
rect 198516 572608 198522 572620
rect 277670 572608 277676 572620
rect 198516 572580 277676 572608
rect 198516 572568 198522 572580
rect 277670 572568 277676 572580
rect 277728 572568 277734 572620
rect 291102 572568 291108 572620
rect 291160 572608 291166 572620
rect 337194 572608 337200 572620
rect 291160 572580 337200 572608
rect 291160 572568 291166 572580
rect 337194 572568 337200 572580
rect 337252 572568 337258 572620
rect 402422 572568 402428 572620
rect 402480 572608 402486 572620
rect 445846 572608 445852 572620
rect 402480 572580 445852 572608
rect 402480 572568 402486 572580
rect 445846 572568 445852 572580
rect 445904 572568 445910 572620
rect 196618 572500 196624 572552
rect 196676 572540 196682 572552
rect 278774 572540 278780 572552
rect 196676 572512 278780 572540
rect 196676 572500 196682 572512
rect 278774 572500 278780 572512
rect 278832 572500 278838 572552
rect 289722 572500 289728 572552
rect 289780 572540 289786 572552
rect 337286 572540 337292 572552
rect 289780 572512 337292 572540
rect 289780 572500 289786 572512
rect 337286 572500 337292 572512
rect 337344 572500 337350 572552
rect 402698 572500 402704 572552
rect 402756 572540 402762 572552
rect 447226 572540 447232 572552
rect 402756 572512 447232 572540
rect 402756 572500 402762 572512
rect 447226 572500 447232 572512
rect 447284 572500 447290 572552
rect 193030 572432 193036 572484
rect 193088 572472 193094 572484
rect 295334 572472 295340 572484
rect 193088 572444 295340 572472
rect 193088 572432 193094 572444
rect 295334 572432 295340 572444
rect 295392 572432 295398 572484
rect 296530 572432 296536 572484
rect 296588 572472 296594 572484
rect 340874 572472 340880 572484
rect 296588 572444 340880 572472
rect 296588 572432 296594 572444
rect 340874 572432 340880 572444
rect 340932 572432 340938 572484
rect 402330 572432 402336 572484
rect 402388 572472 402394 572484
rect 449986 572472 449992 572484
rect 402388 572444 449992 572472
rect 402388 572432 402394 572444
rect 449986 572432 449992 572444
rect 450044 572432 450050 572484
rect 194410 572364 194416 572416
rect 194468 572404 194474 572416
rect 298094 572404 298100 572416
rect 194468 572376 298100 572404
rect 194468 572364 194474 572376
rect 298094 572364 298100 572376
rect 298152 572364 298158 572416
rect 299198 572364 299204 572416
rect 299256 572404 299262 572416
rect 341334 572404 341340 572416
rect 299256 572376 341340 572404
rect 299256 572364 299262 572376
rect 341334 572364 341340 572376
rect 341392 572364 341398 572416
rect 402606 572364 402612 572416
rect 402664 572404 402670 572416
rect 452654 572404 452660 572416
rect 402664 572376 452660 572404
rect 402664 572364 402670 572376
rect 452654 572364 452660 572376
rect 452712 572364 452718 572416
rect 194318 572296 194324 572348
rect 194376 572336 194382 572348
rect 299474 572336 299480 572348
rect 194376 572308 299480 572336
rect 194376 572296 194382 572308
rect 299474 572296 299480 572308
rect 299532 572296 299538 572348
rect 399754 572296 399760 572348
rect 399812 572336 399818 572348
rect 454126 572336 454132 572348
rect 399812 572308 454132 572336
rect 399812 572296 399818 572308
rect 454126 572296 454132 572308
rect 454184 572296 454190 572348
rect 192938 572228 192944 572280
rect 192996 572268 193002 572280
rect 298186 572268 298192 572280
rect 192996 572240 298192 572268
rect 192996 572228 193002 572240
rect 298186 572228 298192 572240
rect 298244 572228 298250 572280
rect 298922 572228 298928 572280
rect 298980 572268 298986 572280
rect 342530 572268 342536 572280
rect 298980 572240 342536 572268
rect 298980 572228 298986 572240
rect 342530 572228 342536 572240
rect 342588 572228 342594 572280
rect 399570 572228 399576 572280
rect 399628 572268 399634 572280
rect 456886 572268 456892 572280
rect 399628 572240 456892 572268
rect 399628 572228 399634 572240
rect 456886 572228 456892 572240
rect 456944 572228 456950 572280
rect 194502 572160 194508 572212
rect 194560 572200 194566 572212
rect 302234 572200 302240 572212
rect 194560 572172 302240 572200
rect 194560 572160 194566 572172
rect 302234 572160 302240 572172
rect 302292 572160 302298 572212
rect 399662 572160 399668 572212
rect 399720 572200 399726 572212
rect 459278 572200 459284 572212
rect 399720 572172 459284 572200
rect 399720 572160 399726 572172
rect 459278 572160 459284 572172
rect 459336 572160 459342 572212
rect 193122 572092 193128 572144
rect 193180 572132 193186 572144
rect 300854 572132 300860 572144
rect 193180 572104 300860 572132
rect 193180 572092 193186 572104
rect 300854 572092 300860 572104
rect 300912 572092 300918 572144
rect 399938 572092 399944 572144
rect 399996 572132 400002 572144
rect 461302 572132 461308 572144
rect 399996 572104 461308 572132
rect 399996 572092 400002 572104
rect 461302 572092 461308 572104
rect 461360 572092 461366 572144
rect 192754 572024 192760 572076
rect 192812 572064 192818 572076
rect 303614 572064 303620 572076
rect 192812 572036 303620 572064
rect 192812 572024 192818 572036
rect 303614 572024 303620 572036
rect 303672 572024 303678 572076
rect 399478 572024 399484 572076
rect 399536 572064 399542 572076
rect 463786 572064 463792 572076
rect 399536 572036 463792 572064
rect 399536 572024 399542 572036
rect 463786 572024 463792 572036
rect 463844 572024 463850 572076
rect 71682 571956 71688 572008
rect 71740 571996 71746 572008
rect 182910 571996 182916 572008
rect 71740 571968 182916 571996
rect 71740 571956 71746 571968
rect 182910 571956 182916 571968
rect 182968 571956 182974 572008
rect 194134 571956 194140 572008
rect 194192 571996 194198 572008
rect 304994 571996 305000 572008
rect 194192 571968 305000 571996
rect 194192 571956 194198 571968
rect 304994 571956 305000 571968
rect 305052 571956 305058 572008
rect 399846 571956 399852 572008
rect 399904 571996 399910 572008
rect 466454 571996 466460 572008
rect 399904 571968 466460 571996
rect 399904 571956 399910 571968
rect 466454 571956 466460 571968
rect 466512 571956 466518 572008
rect 199470 571888 199476 571940
rect 199528 571928 199534 571940
rect 274634 571928 274640 571940
rect 199528 571900 274640 571928
rect 199528 571888 199534 571900
rect 274634 571888 274640 571900
rect 274692 571888 274698 571940
rect 293770 571888 293776 571940
rect 293828 571928 293834 571940
rect 338574 571928 338580 571940
rect 293828 571900 338580 571928
rect 293828 571888 293834 571900
rect 338574 571888 338580 571900
rect 338632 571888 338638 571940
rect 402514 571888 402520 571940
rect 402572 571928 402578 571940
rect 441798 571928 441804 571940
rect 402572 571900 441804 571928
rect 402572 571888 402578 571900
rect 441798 571888 441804 571900
rect 441856 571888 441862 571940
rect 199654 571820 199660 571872
rect 199712 571860 199718 571872
rect 273254 571860 273260 571872
rect 199712 571832 273260 571860
rect 199712 571820 199718 571832
rect 273254 571820 273260 571832
rect 273312 571820 273318 571872
rect 294690 571820 294696 571872
rect 294748 571860 294754 571872
rect 339862 571860 339868 571872
rect 294748 571832 339868 571860
rect 294748 571820 294754 571832
rect 339862 571820 339868 571832
rect 339920 571820 339926 571872
rect 405458 571820 405464 571872
rect 405516 571860 405522 571872
rect 440326 571860 440332 571872
rect 405516 571832 440332 571860
rect 405516 571820 405522 571832
rect 440326 571820 440332 571832
rect 440384 571820 440390 571872
rect 405642 571752 405648 571804
rect 405700 571792 405706 571804
rect 436186 571792 436192 571804
rect 405700 571764 436192 571792
rect 405700 571752 405706 571764
rect 436186 571752 436192 571764
rect 436244 571752 436250 571804
rect 125502 570664 125508 570716
rect 125560 570704 125566 570716
rect 193950 570704 193956 570716
rect 125560 570676 193956 570704
rect 125560 570664 125566 570676
rect 193950 570664 193956 570676
rect 194008 570664 194014 570716
rect 88242 570596 88248 570648
rect 88300 570636 88306 570648
rect 181622 570636 181628 570648
rect 88300 570608 181628 570636
rect 88300 570596 88306 570608
rect 181622 570596 181628 570608
rect 181680 570596 181686 570648
rect 237190 570596 237196 570648
rect 237248 570636 237254 570648
rect 344370 570636 344376 570648
rect 237248 570608 344376 570636
rect 237248 570596 237254 570608
rect 344370 570596 344376 570608
rect 344428 570596 344434 570648
rect 365254 570596 365260 570648
rect 365312 570636 365318 570648
rect 452746 570636 452752 570648
rect 365312 570608 452752 570636
rect 365312 570596 365318 570608
rect 452746 570596 452752 570608
rect 452804 570596 452810 570648
rect 128262 569440 128268 569492
rect 128320 569480 128326 569492
rect 195330 569480 195336 569492
rect 128320 569452 195336 569480
rect 128320 569440 128326 569452
rect 195330 569440 195336 569452
rect 195388 569440 195394 569492
rect 194226 569372 194232 569424
rect 194284 569412 194290 569424
rect 270494 569412 270500 569424
rect 194284 569384 270500 569412
rect 194284 569372 194290 569384
rect 270494 569372 270500 569384
rect 270552 569372 270558 569424
rect 191650 569304 191656 569356
rect 191708 569344 191714 569356
rect 269206 569344 269212 569356
rect 191708 569316 269212 569344
rect 191708 569304 191714 569316
rect 269206 569304 269212 569316
rect 269264 569304 269270 569356
rect 192846 569236 192852 569288
rect 192904 569276 192910 569288
rect 271874 569276 271880 569288
rect 192904 569248 271880 569276
rect 192904 569236 192910 569248
rect 271874 569236 271880 569248
rect 271932 569236 271938 569288
rect 91002 569168 91008 569220
rect 91060 569208 91066 569220
rect 192478 569208 192484 569220
rect 91060 569180 192484 569208
rect 91060 569168 91066 569180
rect 192478 569168 192484 569180
rect 192536 569168 192542 569220
rect 253750 569168 253756 569220
rect 253808 569208 253814 569220
rect 347038 569208 347044 569220
rect 253808 569180 347044 569208
rect 253808 569168 253814 569180
rect 347038 569168 347044 569180
rect 347096 569168 347102 569220
rect 367738 569168 367744 569220
rect 367796 569208 367802 569220
rect 455506 569208 455512 569220
rect 367796 569180 455512 569208
rect 367796 569168 367802 569180
rect 455506 569168 455512 569180
rect 455564 569168 455570 569220
rect 131022 567876 131028 567928
rect 131080 567916 131086 567928
rect 167730 567916 167736 567928
rect 131080 567888 167736 567916
rect 131080 567876 131086 567888
rect 167730 567876 167736 567888
rect 167788 567876 167794 567928
rect 108942 567808 108948 567860
rect 109000 567848 109006 567860
rect 176194 567848 176200 567860
rect 109000 567820 176200 567848
rect 109000 567808 109006 567820
rect 176194 567808 176200 567820
rect 176252 567808 176258 567860
rect 253106 567808 253112 567860
rect 253164 567848 253170 567860
rect 347130 567848 347136 567860
rect 253164 567820 347136 567848
rect 253164 567808 253170 567820
rect 347130 567808 347136 567820
rect 347188 567808 347194 567860
rect 373994 567808 374000 567860
rect 374052 567848 374058 567860
rect 461118 567848 461124 567860
rect 374052 567820 461124 567848
rect 374052 567808 374058 567820
rect 461118 567808 461124 567820
rect 461176 567808 461182 567860
rect 74442 566448 74448 566500
rect 74500 566488 74506 566500
rect 184474 566488 184480 566500
rect 74500 566460 184480 566488
rect 74500 566448 74506 566460
rect 184474 566448 184480 566460
rect 184532 566448 184538 566500
rect 356422 566448 356428 566500
rect 356480 566488 356486 566500
rect 444466 566488 444472 566500
rect 356480 566460 444472 566488
rect 356480 566448 356486 566460
rect 444466 566448 444472 566460
rect 444524 566448 444530 566500
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 400950 565876 400956 565888
rect 3476 565848 400956 565876
rect 3476 565836 3482 565848
rect 400950 565836 400956 565848
rect 401008 565836 401014 565888
rect 75822 565156 75828 565208
rect 75880 565196 75886 565208
rect 188522 565196 188528 565208
rect 75880 565168 188528 565196
rect 75880 565156 75886 565168
rect 188522 565156 188528 565168
rect 188580 565156 188586 565208
rect 3510 565088 3516 565140
rect 3568 565128 3574 565140
rect 408034 565128 408040 565140
rect 3568 565100 408040 565128
rect 3568 565088 3574 565100
rect 408034 565088 408040 565100
rect 408092 565088 408098 565140
rect 142062 563796 142068 563848
rect 142120 563836 142126 563848
rect 168190 563836 168196 563848
rect 142120 563808 168196 563836
rect 142120 563796 142126 563808
rect 168190 563796 168196 563808
rect 168248 563796 168254 563848
rect 78582 563728 78588 563780
rect 78640 563768 78646 563780
rect 170950 563768 170956 563780
rect 78640 563740 170956 563768
rect 78640 563728 78646 563740
rect 170950 563728 170956 563740
rect 171008 563728 171014 563780
rect 357710 563728 357716 563780
rect 357768 563768 357774 563780
rect 444558 563768 444564 563780
rect 357768 563740 444564 563768
rect 357768 563728 357774 563740
rect 444558 563728 444564 563740
rect 444616 563728 444622 563780
rect 3786 563660 3792 563712
rect 3844 563700 3850 563712
rect 408126 563700 408132 563712
rect 3844 563672 408132 563700
rect 3844 563660 3850 563672
rect 408126 563660 408132 563672
rect 408184 563660 408190 563712
rect 29730 563116 29736 563168
rect 29788 563156 29794 563168
rect 29788 563128 35894 563156
rect 29788 563116 29794 563128
rect 29638 563048 29644 563100
rect 29696 563088 29702 563100
rect 35710 563088 35716 563100
rect 29696 563060 35716 563088
rect 29696 563048 29702 563060
rect 35710 563048 35716 563060
rect 35768 563048 35774 563100
rect 35866 563088 35894 563128
rect 46750 563088 46756 563100
rect 35866 563060 46756 563088
rect 46750 563048 46756 563060
rect 46808 563048 46814 563100
rect 566458 563048 566464 563100
rect 566516 563088 566522 563100
rect 580166 563088 580172 563100
rect 566516 563060 580172 563088
rect 566516 563048 566522 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 28718 562572 28724 562624
rect 28776 562612 28782 562624
rect 29730 562612 29736 562624
rect 28776 562584 29736 562612
rect 28776 562572 28782 562584
rect 29730 562572 29736 562584
rect 29788 562572 29794 562624
rect 28810 562300 28816 562352
rect 28868 562340 28874 562352
rect 29822 562340 29828 562352
rect 28868 562312 29828 562340
rect 28868 562300 28874 562312
rect 29822 562300 29828 562312
rect 29880 562340 29886 562352
rect 48038 562340 48044 562352
rect 29880 562312 48044 562340
rect 29880 562300 29886 562312
rect 48038 562300 48044 562312
rect 48096 562300 48102 562352
rect 60642 562300 60648 562352
rect 60700 562340 60706 562352
rect 179046 562340 179052 562352
rect 60700 562312 179052 562340
rect 60700 562300 60706 562312
rect 179046 562300 179052 562312
rect 179104 562300 179110 562352
rect 253842 562300 253848 562352
rect 253900 562340 253906 562352
rect 348510 562340 348516 562352
rect 253900 562312 348516 562340
rect 253900 562300 253906 562312
rect 348510 562300 348516 562312
rect 348568 562300 348574 562352
rect 351362 562300 351368 562352
rect 351420 562340 351426 562352
rect 438946 562340 438952 562352
rect 351420 562312 438952 562340
rect 351420 562300 351426 562312
rect 438946 562300 438952 562312
rect 439004 562300 439010 562352
rect 28626 561960 28632 562012
rect 28684 562000 28690 562012
rect 29638 562000 29644 562012
rect 28684 561972 29644 562000
rect 28684 561960 28690 561972
rect 29638 561960 29644 561972
rect 29696 561960 29702 562012
rect 375282 560940 375288 560992
rect 375340 560980 375346 560992
rect 462406 560980 462412 560992
rect 375340 560952 462412 560980
rect 375340 560940 375346 560952
rect 462406 560940 462412 560952
rect 462464 560940 462470 560992
rect 377766 559512 377772 559564
rect 377824 559552 377830 559564
rect 464338 559552 464344 559564
rect 377824 559524 464344 559552
rect 377824 559512 377830 559524
rect 464338 559512 464344 559524
rect 464396 559512 464402 559564
rect 379054 558152 379060 558204
rect 379112 558192 379118 558204
rect 466638 558192 466644 558204
rect 379112 558164 466644 558192
rect 379112 558152 379118 558164
rect 466638 558152 466644 558164
rect 466696 558152 466702 558204
rect 355134 556792 355140 556844
rect 355192 556832 355198 556844
rect 442994 556832 443000 556844
rect 355192 556804 443000 556832
rect 355192 556792 355198 556804
rect 442994 556792 443000 556804
rect 443052 556792 443058 556844
rect 381538 555432 381544 555484
rect 381596 555472 381602 555484
rect 468478 555472 468484 555484
rect 381596 555444 468484 555472
rect 381596 555432 381602 555444
rect 468478 555432 468484 555444
rect 468536 555432 468542 555484
rect 380342 554004 380348 554056
rect 380400 554044 380406 554056
rect 467834 554044 467840 554056
rect 380400 554016 467840 554044
rect 380400 554004 380406 554016
rect 467834 554004 467840 554016
rect 467892 554004 467898 554056
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 28258 553432 28264 553444
rect 3476 553404 28264 553432
rect 3476 553392 3482 553404
rect 28258 553392 28264 553404
rect 28316 553392 28322 553444
rect 376570 552644 376576 552696
rect 376628 552684 376634 552696
rect 463694 552684 463700 552696
rect 376628 552656 463700 552684
rect 376628 552644 376634 552656
rect 463694 552644 463700 552656
rect 463752 552644 463758 552696
rect 369026 551284 369032 551336
rect 369084 551324 369090 551336
rect 455598 551324 455604 551336
rect 369084 551296 455604 551324
rect 369084 551284 369090 551296
rect 455598 551284 455604 551296
rect 455656 551284 455662 551336
rect 348510 550536 348516 550588
rect 348568 550576 348574 550588
rect 485038 550576 485044 550588
rect 348568 550548 485044 550576
rect 348568 550536 348574 550548
rect 485038 550536 485044 550548
rect 485096 550536 485102 550588
rect 347130 549176 347136 549228
rect 347188 549216 347194 549228
rect 347590 549216 347596 549228
rect 347188 549188 347596 549216
rect 347188 549176 347194 549188
rect 347590 549176 347596 549188
rect 347648 549216 347654 549228
rect 487798 549216 487804 549228
rect 347648 549188 487804 549216
rect 347648 549176 347654 549188
rect 487798 549176 487804 549188
rect 487856 549176 487862 549228
rect 347038 547816 347044 547868
rect 347096 547856 347102 547868
rect 490558 547856 490564 547868
rect 347096 547828 490564 547856
rect 347096 547816 347102 547828
rect 490558 547816 490564 547828
rect 490616 547816 490622 547868
rect 346394 546456 346400 546508
rect 346452 546496 346458 546508
rect 347038 546496 347044 546508
rect 346452 546468 347044 546496
rect 346452 546456 346458 546468
rect 347038 546456 347044 546468
rect 347096 546456 347102 546508
rect 254578 545708 254584 545760
rect 254636 545748 254642 545760
rect 345106 545748 345112 545760
rect 254636 545720 345112 545748
rect 254636 545708 254642 545720
rect 345106 545708 345112 545720
rect 345164 545748 345170 545760
rect 480898 545748 480904 545760
rect 345164 545720 480904 545748
rect 345164 545708 345170 545720
rect 480898 545708 480904 545720
rect 480956 545708 480962 545760
rect 343818 545028 343824 545080
rect 343876 545068 343882 545080
rect 344370 545068 344376 545080
rect 343876 545040 344376 545068
rect 343876 545028 343882 545040
rect 344370 545028 344376 545040
rect 344428 545068 344434 545080
rect 507946 545068 507952 545080
rect 344428 545040 507952 545068
rect 344428 545028 344434 545040
rect 507946 545028 507952 545040
rect 508004 545028 508010 545080
rect 238570 544348 238576 544400
rect 238628 544388 238634 544400
rect 342622 544388 342628 544400
rect 238628 544360 342628 544388
rect 238628 544348 238634 544360
rect 342622 544348 342628 544360
rect 342680 544348 342686 544400
rect 342622 543668 342628 543720
rect 342680 543708 342686 543720
rect 506474 543708 506480 543720
rect 342680 543680 506480 543708
rect 342680 543668 342686 543680
rect 506474 543668 506480 543680
rect 506532 543668 506538 543720
rect 238662 542988 238668 543040
rect 238720 543028 238726 543040
rect 341610 543028 341616 543040
rect 238720 543000 341616 543028
rect 238720 542988 238726 543000
rect 341610 542988 341616 543000
rect 341668 542988 341674 543040
rect 358906 541696 358912 541748
rect 358964 541736 358970 541748
rect 445754 541736 445760 541748
rect 358964 541708 445760 541736
rect 358964 541696 358970 541708
rect 445754 541696 445760 541708
rect 445812 541696 445818 541748
rect 361482 541628 361488 541680
rect 361540 541668 361546 541680
rect 448606 541668 448612 541680
rect 361540 541640 448612 541668
rect 361540 541628 361546 541640
rect 448606 541628 448612 541640
rect 448664 541628 448670 541680
rect 384114 540812 384120 540864
rect 384172 540852 384178 540864
rect 470686 540852 470692 540864
rect 384172 540824 470692 540852
rect 384172 540812 384178 540824
rect 470686 540812 470692 540824
rect 470744 540812 470750 540864
rect 385310 540744 385316 540796
rect 385368 540784 385374 540796
rect 471974 540784 471980 540796
rect 385368 540756 471980 540784
rect 385368 540744 385374 540756
rect 471974 540744 471980 540756
rect 472032 540744 472038 540796
rect 386598 540676 386604 540728
rect 386656 540716 386662 540728
rect 473354 540716 473360 540728
rect 386656 540688 473360 540716
rect 386656 540676 386662 540688
rect 473354 540676 473360 540688
rect 473412 540676 473418 540728
rect 387886 540608 387892 540660
rect 387944 540648 387950 540660
rect 474734 540648 474740 540660
rect 387944 540620 474740 540648
rect 387944 540608 387950 540620
rect 474734 540608 474740 540620
rect 474792 540608 474798 540660
rect 389082 540540 389088 540592
rect 389140 540580 389146 540592
rect 476114 540580 476120 540592
rect 389140 540552 476120 540580
rect 389140 540540 389146 540552
rect 476114 540540 476120 540552
rect 476172 540540 476178 540592
rect 352650 540472 352656 540524
rect 352708 540512 352714 540524
rect 440234 540512 440240 540524
rect 352708 540484 440240 540512
rect 352708 540472 352714 540484
rect 440234 540472 440240 540484
rect 440292 540472 440298 540524
rect 280062 540404 280068 540456
rect 280120 540444 280126 540456
rect 338758 540444 338764 540456
rect 280120 540416 338764 540444
rect 280120 540404 280126 540416
rect 338758 540404 338764 540416
rect 338816 540404 338822 540456
rect 382826 540404 382832 540456
rect 382884 540444 382890 540456
rect 470594 540444 470600 540456
rect 382884 540416 470600 540444
rect 382884 540404 382890 540416
rect 470594 540404 470600 540416
rect 470652 540404 470658 540456
rect 278682 540336 278688 540388
rect 278740 540376 278746 540388
rect 338666 540376 338672 540388
rect 278740 540348 338672 540376
rect 278740 540336 278746 540348
rect 338666 540336 338672 540348
rect 338724 540336 338730 540388
rect 353294 540336 353300 540388
rect 353352 540376 353358 540388
rect 441614 540376 441620 540388
rect 353352 540348 441620 540376
rect 353352 540336 353358 540348
rect 441614 540336 441620 540348
rect 441672 540336 441678 540388
rect 218054 540268 218060 540320
rect 218112 540308 218118 540320
rect 527174 540308 527180 540320
rect 218112 540280 527180 540308
rect 218112 540268 218118 540280
rect 527174 540268 527180 540280
rect 527232 540268 527238 540320
rect 217594 540200 217600 540252
rect 217652 540240 217658 540252
rect 528830 540240 528836 540252
rect 217652 540212 528836 540240
rect 217652 540200 217658 540212
rect 528830 540200 528836 540212
rect 528888 540200 528894 540252
rect 187050 539928 187056 539980
rect 187108 539968 187114 539980
rect 205726 539968 205732 539980
rect 187108 539940 205732 539968
rect 187108 539928 187114 539940
rect 205726 539928 205732 539940
rect 205784 539928 205790 539980
rect 190362 539860 190368 539912
rect 190420 539900 190426 539912
rect 218054 539900 218060 539912
rect 190420 539872 218060 539900
rect 190420 539860 190426 539872
rect 218054 539860 218060 539872
rect 218112 539860 218118 539912
rect 169294 539792 169300 539844
rect 169352 539832 169358 539844
rect 338850 539832 338856 539844
rect 169352 539804 338856 539832
rect 169352 539792 169358 539804
rect 338850 539792 338856 539804
rect 338908 539792 338914 539844
rect 169202 539724 169208 539776
rect 169260 539764 169266 539776
rect 340046 539764 340052 539776
rect 169260 539736 340052 539764
rect 169260 539724 169266 539736
rect 340046 539724 340052 539736
rect 340104 539724 340110 539776
rect 169110 539656 169116 539708
rect 169168 539696 169174 539708
rect 340322 539696 340328 539708
rect 169168 539668 340328 539696
rect 169168 539656 169174 539668
rect 340322 539656 340328 539668
rect 340380 539656 340386 539708
rect 169018 539588 169024 539640
rect 169076 539628 169082 539640
rect 340230 539628 340236 539640
rect 169076 539600 340236 539628
rect 169076 539588 169082 539600
rect 340230 539588 340236 539600
rect 340288 539588 340294 539640
rect 370222 539316 370228 539368
rect 370280 539356 370286 539368
rect 456794 539356 456800 539368
rect 370280 539328 456800 539356
rect 370280 539316 370286 539328
rect 456794 539316 456800 539328
rect 456852 539316 456858 539368
rect 371510 539248 371516 539300
rect 371568 539288 371574 539300
rect 458358 539288 458364 539300
rect 371568 539260 458364 539288
rect 371568 539248 371574 539260
rect 458358 539248 458364 539260
rect 458416 539248 458422 539300
rect 372798 539180 372804 539232
rect 372856 539220 372862 539232
rect 459646 539220 459652 539232
rect 372856 539192 459652 539220
rect 372856 539180 372862 539192
rect 459646 539180 459652 539192
rect 459704 539180 459710 539232
rect 362678 539112 362684 539164
rect 362736 539152 362742 539164
rect 449894 539152 449900 539164
rect 362736 539124 449900 539152
rect 362736 539112 362742 539124
rect 449894 539112 449900 539124
rect 449952 539112 449958 539164
rect 318702 539044 318708 539096
rect 318760 539084 318766 539096
rect 342714 539084 342720 539096
rect 318760 539056 342720 539084
rect 318760 539044 318766 539056
rect 342714 539044 342720 539056
rect 342772 539044 342778 539096
rect 363966 539044 363972 539096
rect 364024 539084 364030 539096
rect 451274 539084 451280 539096
rect 364024 539056 451280 539084
rect 364024 539044 364030 539056
rect 451274 539044 451280 539056
rect 451332 539044 451338 539096
rect 284202 538976 284208 539028
rect 284260 539016 284266 539028
rect 342806 539016 342812 539028
rect 284260 538988 342812 539016
rect 284260 538976 284266 538988
rect 342806 538976 342812 538988
rect 342864 538976 342870 539028
rect 350166 538976 350172 539028
rect 350224 539016 350230 539028
rect 437566 539016 437572 539028
rect 350224 538988 437572 539016
rect 350224 538976 350230 538988
rect 437566 538976 437572 538988
rect 437624 538976 437630 539028
rect 282822 538908 282828 538960
rect 282880 538948 282886 538960
rect 342898 538948 342904 538960
rect 282880 538920 342904 538948
rect 282880 538908 282886 538920
rect 342898 538908 342904 538920
rect 342956 538908 342962 538960
rect 366450 538908 366456 538960
rect 366508 538948 366514 538960
rect 454034 538948 454040 538960
rect 366508 538920 454040 538948
rect 366508 538908 366514 538920
rect 454034 538908 454040 538920
rect 454092 538908 454098 538960
rect 281442 538840 281448 538892
rect 281500 538880 281506 538892
rect 341702 538880 341708 538892
rect 281500 538852 341708 538880
rect 281500 538840 281506 538852
rect 341702 538840 341708 538852
rect 341760 538840 341766 538892
rect 407666 538840 407672 538892
rect 407724 538880 407730 538892
rect 540790 538880 540796 538892
rect 407724 538852 540796 538880
rect 407724 538840 407730 538852
rect 540790 538840 540796 538852
rect 540848 538840 540854 538892
rect 570690 524424 570696 524476
rect 570748 524464 570754 524476
rect 580166 524464 580172 524476
rect 570748 524436 580172 524464
rect 570748 524424 570754 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 18598 514808 18604 514820
rect 3568 514780 18604 514808
rect 3568 514768 3574 514780
rect 18598 514768 18604 514780
rect 18656 514768 18662 514820
rect 565170 510620 565176 510672
rect 565228 510660 565234 510672
rect 580166 510660 580172 510672
rect 565228 510632 580172 510660
rect 565228 510620 565234 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 28718 501004 28724 501016
rect 3108 500976 28724 501004
rect 3108 500964 3114 500976
rect 28718 500964 28724 500976
rect 28776 500964 28782 501016
rect 339310 491240 339316 491292
rect 339368 491280 339374 491292
rect 340322 491280 340328 491292
rect 339368 491252 340328 491280
rect 339368 491240 339374 491252
rect 340322 491240 340328 491252
rect 340380 491280 340386 491292
rect 407206 491280 407212 491292
rect 340380 491252 407212 491280
rect 340380 491240 340386 491252
rect 407206 491240 407212 491252
rect 407264 491240 407270 491292
rect 339402 491172 339408 491224
rect 339460 491212 339466 491224
rect 340230 491212 340236 491224
rect 339460 491184 340236 491212
rect 339460 491172 339466 491184
rect 340230 491172 340236 491184
rect 340288 491212 340294 491224
rect 407114 491212 407120 491224
rect 340288 491184 407120 491212
rect 340288 491172 340294 491184
rect 407114 491172 407120 491184
rect 407172 491172 407178 491224
rect 340046 488452 340052 488504
rect 340104 488492 340110 488504
rect 407114 488492 407120 488504
rect 340104 488464 407120 488492
rect 340104 488452 340110 488464
rect 407114 488452 407120 488464
rect 407172 488452 407178 488504
rect 169662 487092 169668 487144
rect 169720 487132 169726 487144
rect 187050 487132 187056 487144
rect 169720 487104 187056 487132
rect 169720 487092 169726 487104
rect 187050 487092 187056 487104
rect 187108 487092 187114 487144
rect 338850 487092 338856 487144
rect 338908 487132 338914 487144
rect 407114 487132 407120 487144
rect 338908 487104 407120 487132
rect 338908 487092 338914 487104
rect 407114 487092 407120 487104
rect 407172 487092 407178 487144
rect 168834 486412 168840 486464
rect 168892 486452 168898 486464
rect 178678 486452 178684 486464
rect 168892 486424 178684 486452
rect 168892 486412 168898 486424
rect 178678 486412 178684 486424
rect 178736 486412 178742 486464
rect 339402 484372 339408 484424
rect 339460 484412 339466 484424
rect 340230 484412 340236 484424
rect 339460 484384 340236 484412
rect 339460 484372 339466 484384
rect 340230 484372 340236 484384
rect 340288 484412 340294 484424
rect 407114 484412 407120 484424
rect 340288 484384 407120 484412
rect 340288 484372 340294 484384
rect 407114 484372 407120 484384
rect 407172 484372 407178 484424
rect 577590 484372 577596 484424
rect 577648 484412 577654 484424
rect 580626 484412 580632 484424
rect 577648 484384 580632 484412
rect 577648 484372 577654 484384
rect 580626 484372 580632 484384
rect 580684 484372 580690 484424
rect 340046 483012 340052 483064
rect 340104 483052 340110 483064
rect 407114 483052 407120 483064
rect 340104 483024 407120 483052
rect 340104 483012 340110 483024
rect 407114 483012 407120 483024
rect 407172 483012 407178 483064
rect 338850 481652 338856 481704
rect 338908 481692 338914 481704
rect 407114 481692 407120 481704
rect 338908 481664 407120 481692
rect 338908 481652 338914 481664
rect 407114 481652 407120 481664
rect 407172 481652 407178 481704
rect 165522 476076 165528 476128
rect 165580 476116 165586 476128
rect 167178 476116 167184 476128
rect 165580 476088 167184 476116
rect 165580 476076 165586 476088
rect 167178 476076 167184 476088
rect 167236 476076 167242 476128
rect 3510 475532 3516 475584
rect 3568 475572 3574 475584
rect 166718 475572 166724 475584
rect 3568 475544 166724 475572
rect 3568 475532 3574 475544
rect 166718 475532 166724 475544
rect 166776 475532 166782 475584
rect 28534 475464 28540 475516
rect 28592 475504 28598 475516
rect 42794 475504 42800 475516
rect 28592 475476 42800 475504
rect 28592 475464 28598 475476
rect 42794 475464 42800 475476
rect 42852 475464 42858 475516
rect 151354 475396 151360 475448
rect 151412 475436 151418 475448
rect 151722 475436 151728 475448
rect 151412 475408 151728 475436
rect 151412 475396 151418 475408
rect 151722 475396 151728 475408
rect 151780 475436 151786 475448
rect 167086 475436 167092 475448
rect 151780 475408 167092 475436
rect 151780 475396 151786 475408
rect 167086 475396 167092 475408
rect 167144 475396 167150 475448
rect 29638 475328 29644 475380
rect 29696 475368 29702 475380
rect 34514 475368 34520 475380
rect 29696 475340 34520 475368
rect 29696 475328 29702 475340
rect 34514 475328 34520 475340
rect 34572 475328 34578 475380
rect 42794 475368 42800 475380
rect 35866 475340 42800 475368
rect 28442 475260 28448 475312
rect 28500 475300 28506 475312
rect 35866 475300 35894 475340
rect 42794 475328 42800 475340
rect 42852 475328 42858 475380
rect 141786 475328 141792 475380
rect 141844 475368 141850 475380
rect 175918 475368 175924 475380
rect 141844 475340 175924 475368
rect 141844 475328 141850 475340
rect 175918 475328 175924 475340
rect 175976 475328 175982 475380
rect 28500 475272 35894 475300
rect 28500 475260 28506 475272
rect 129642 475260 129648 475312
rect 129700 475300 129706 475312
rect 173894 475300 173900 475312
rect 129700 475272 173900 475300
rect 129700 475260 129706 475272
rect 173894 475260 173900 475272
rect 173952 475300 173958 475312
rect 174906 475300 174912 475312
rect 173952 475272 174912 475300
rect 173952 475260 173958 475272
rect 174906 475260 174912 475272
rect 174964 475260 174970 475312
rect 126882 475192 126888 475244
rect 126940 475232 126946 475244
rect 176654 475232 176660 475244
rect 126940 475204 176660 475232
rect 126940 475192 126946 475204
rect 176654 475192 176660 475204
rect 176712 475192 176718 475244
rect 131022 475124 131028 475176
rect 131080 475164 131086 475176
rect 181898 475164 181904 475176
rect 131080 475136 181904 475164
rect 131080 475124 131086 475136
rect 181898 475124 181904 475136
rect 181956 475124 181962 475176
rect 128262 475056 128268 475108
rect 128320 475096 128326 475108
rect 187694 475096 187700 475108
rect 128320 475068 187700 475096
rect 128320 475056 128326 475068
rect 187694 475056 187700 475068
rect 187752 475056 187758 475108
rect 115474 474988 115480 475040
rect 115532 475028 115538 475040
rect 175274 475028 175280 475040
rect 115532 475000 175280 475028
rect 115532 474988 115538 475000
rect 175274 474988 175280 475000
rect 175332 474988 175338 475040
rect 110322 474920 110328 474972
rect 110380 474960 110386 474972
rect 171778 474960 171784 474972
rect 110380 474932 171784 474960
rect 110380 474920 110386 474932
rect 171778 474920 171784 474932
rect 171836 474960 171842 474972
rect 172422 474960 172428 474972
rect 171836 474932 172428 474960
rect 171836 474920 171842 474932
rect 172422 474920 172428 474932
rect 172480 474920 172486 474972
rect 121178 474852 121184 474904
rect 121236 474892 121242 474904
rect 128998 474892 129004 474904
rect 121236 474864 129004 474892
rect 121236 474852 121242 474864
rect 128998 474852 129004 474864
rect 129056 474852 129062 474904
rect 129550 474852 129556 474904
rect 129608 474892 129614 474904
rect 193858 474892 193864 474904
rect 129608 474864 193864 474892
rect 129608 474852 129614 474864
rect 193858 474852 193864 474864
rect 193916 474852 193922 474904
rect 60642 474784 60648 474836
rect 60700 474824 60706 474836
rect 167546 474824 167552 474836
rect 60700 474796 167552 474824
rect 60700 474784 60706 474796
rect 167546 474784 167552 474796
rect 167604 474784 167610 474836
rect 175918 474784 175924 474836
rect 175976 474824 175982 474836
rect 199194 474824 199200 474836
rect 175976 474796 199200 474824
rect 175976 474784 175982 474796
rect 199194 474784 199200 474796
rect 199252 474784 199258 474836
rect 121362 474716 121368 474768
rect 121420 474756 121426 474768
rect 126238 474756 126244 474768
rect 121420 474728 126244 474756
rect 121420 474716 121426 474728
rect 126238 474716 126244 474728
rect 126296 474716 126302 474768
rect 174906 474716 174912 474768
rect 174964 474756 174970 474768
rect 199286 474756 199292 474768
rect 174964 474728 199292 474756
rect 174964 474716 174970 474728
rect 199286 474716 199292 474728
rect 199344 474716 199350 474768
rect 28442 474648 28448 474700
rect 28500 474688 28506 474700
rect 29638 474688 29644 474700
rect 28500 474660 29644 474688
rect 28500 474648 28506 474660
rect 29638 474648 29644 474660
rect 29696 474648 29702 474700
rect 136542 474172 136548 474224
rect 136600 474212 136606 474224
rect 137278 474212 137284 474224
rect 136600 474184 137284 474212
rect 136600 474172 136606 474184
rect 137278 474172 137284 474184
rect 137336 474172 137342 474224
rect 139302 474104 139308 474156
rect 139360 474144 139366 474156
rect 181714 474144 181720 474156
rect 139360 474116 181720 474144
rect 139360 474104 139366 474116
rect 181714 474104 181720 474116
rect 181772 474104 181778 474156
rect 136358 474036 136364 474088
rect 136416 474076 136422 474088
rect 192570 474076 192576 474088
rect 136416 474048 192576 474076
rect 136416 474036 136422 474048
rect 192570 474036 192576 474048
rect 192628 474036 192634 474088
rect 96522 473968 96528 474020
rect 96580 474008 96586 474020
rect 179138 474008 179144 474020
rect 96580 473980 179144 474008
rect 96580 473968 96586 473980
rect 179138 473968 179144 473980
rect 179196 473968 179202 474020
rect 143350 472744 143356 472796
rect 143408 472784 143414 472796
rect 177390 472784 177396 472796
rect 143408 472756 177396 472784
rect 143408 472744 143414 472756
rect 177390 472744 177396 472756
rect 177448 472744 177454 472796
rect 133690 472676 133696 472728
rect 133748 472716 133754 472728
rect 191374 472716 191380 472728
rect 133748 472688 191380 472716
rect 133748 472676 133754 472688
rect 191374 472676 191380 472688
rect 191432 472676 191438 472728
rect 93762 472608 93768 472660
rect 93820 472648 93826 472660
rect 180150 472648 180156 472660
rect 93820 472620 180156 472648
rect 93820 472608 93826 472620
rect 180150 472608 180156 472620
rect 180208 472608 180214 472660
rect 177390 471996 177396 472048
rect 177448 472036 177454 472048
rect 195238 472036 195244 472048
rect 177448 472008 195244 472036
rect 177448 471996 177454 472008
rect 195238 471996 195244 472008
rect 195296 471996 195302 472048
rect 131022 471384 131028 471436
rect 131080 471424 131086 471436
rect 189902 471424 189908 471436
rect 131080 471396 189908 471424
rect 131080 471384 131086 471396
rect 189902 471384 189908 471396
rect 189960 471384 189966 471436
rect 112990 471316 112996 471368
rect 113048 471356 113054 471368
rect 180242 471356 180248 471368
rect 113048 471328 180248 471356
rect 113048 471316 113054 471328
rect 180242 471316 180248 471328
rect 180300 471316 180306 471368
rect 86862 471248 86868 471300
rect 86920 471288 86926 471300
rect 183094 471288 183100 471300
rect 86920 471260 183100 471288
rect 86920 471248 86926 471260
rect 183094 471248 183100 471260
rect 183152 471248 183158 471300
rect 566550 470568 566556 470620
rect 566608 470608 566614 470620
rect 580166 470608 580172 470620
rect 566608 470580 580172 470608
rect 566608 470568 566614 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 124030 469956 124036 470008
rect 124088 469996 124094 470008
rect 174814 469996 174820 470008
rect 124088 469968 174820 469996
rect 124088 469956 124094 469968
rect 174814 469956 174820 469968
rect 174872 469956 174878 470008
rect 111610 469888 111616 469940
rect 111668 469928 111674 469940
rect 191466 469928 191472 469940
rect 111668 469900 191472 469928
rect 111668 469888 111674 469900
rect 191466 469888 191472 469900
rect 191524 469888 191530 469940
rect 84102 469820 84108 469872
rect 84160 469860 84166 469872
rect 185854 469860 185860 469872
rect 84160 469832 185860 469860
rect 84160 469820 84166 469832
rect 185854 469820 185860 469832
rect 185912 469820 185918 469872
rect 121270 468596 121276 468648
rect 121328 468636 121334 468648
rect 192662 468636 192668 468648
rect 121328 468608 192668 468636
rect 121328 468596 121334 468608
rect 192662 468596 192668 468608
rect 192720 468596 192726 468648
rect 108850 468528 108856 468580
rect 108908 468568 108914 468580
rect 187234 468568 187240 468580
rect 108908 468540 187240 468568
rect 108908 468528 108914 468540
rect 187234 468528 187240 468540
rect 187292 468528 187298 468580
rect 75822 468460 75828 468512
rect 75880 468500 75886 468512
rect 193766 468500 193772 468512
rect 75880 468472 193772 468500
rect 75880 468460 75886 468472
rect 193766 468460 193772 468472
rect 193824 468460 193830 468512
rect 115750 467236 115756 467288
rect 115808 467276 115814 467288
rect 176286 467276 176292 467288
rect 115808 467248 176292 467276
rect 115808 467236 115814 467248
rect 176286 467236 176292 467248
rect 176344 467236 176350 467288
rect 106182 467168 106188 467220
rect 106240 467208 106246 467220
rect 184658 467208 184664 467220
rect 106240 467180 184664 467208
rect 106240 467168 106246 467180
rect 184658 467168 184664 467180
rect 184716 467168 184722 467220
rect 78582 467100 78588 467152
rect 78640 467140 78646 467152
rect 195146 467140 195152 467152
rect 78640 467112 195152 467140
rect 78640 467100 78646 467112
rect 195146 467100 195152 467112
rect 195204 467100 195210 467152
rect 74442 465672 74448 465724
rect 74500 465712 74506 465724
rect 177758 465712 177764 465724
rect 74500 465684 177764 465712
rect 74500 465672 74506 465684
rect 177758 465672 177764 465684
rect 177816 465672 177822 465724
rect 136542 464448 136548 464500
rect 136600 464488 136606 464500
rect 169846 464488 169852 464500
rect 136600 464460 169852 464488
rect 136600 464448 136606 464460
rect 169846 464448 169852 464460
rect 169904 464448 169910 464500
rect 100662 464380 100668 464432
rect 100720 464420 100726 464432
rect 177666 464420 177672 464432
rect 100720 464392 177672 464420
rect 100720 464380 100726 464392
rect 177666 464380 177672 464392
rect 177724 464380 177730 464432
rect 68922 464312 68928 464364
rect 68980 464352 68986 464364
rect 187418 464352 187424 464364
rect 68980 464324 187424 464352
rect 68980 464312 68986 464324
rect 187418 464312 187424 464324
rect 187476 464312 187482 464364
rect 169846 463700 169852 463752
rect 169904 463740 169910 463752
rect 170398 463740 170404 463752
rect 169904 463712 170404 463740
rect 169904 463700 169910 463712
rect 170398 463700 170404 463712
rect 170456 463740 170462 463752
rect 176470 463740 176476 463752
rect 170456 463712 176476 463740
rect 170456 463700 170462 463712
rect 176470 463700 176476 463712
rect 176528 463700 176534 463752
rect 339402 463700 339408 463752
rect 339460 463740 339466 463752
rect 340322 463740 340328 463752
rect 339460 463712 340328 463740
rect 339460 463700 339466 463712
rect 340322 463700 340328 463712
rect 340380 463740 340386 463752
rect 407114 463740 407120 463752
rect 340380 463712 407120 463740
rect 340380 463700 340386 463712
rect 407114 463700 407120 463712
rect 407172 463700 407178 463752
rect 339126 462952 339132 463004
rect 339184 462992 339190 463004
rect 407114 462992 407120 463004
rect 339184 462964 407120 462992
rect 339184 462952 339190 462964
rect 407114 462952 407120 462964
rect 407172 462992 407178 463004
rect 407666 462992 407672 463004
rect 407172 462964 407672 462992
rect 407172 462952 407178 462964
rect 407666 462952 407672 462964
rect 407724 462952 407730 463004
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 191558 462380 191564 462392
rect 3568 462352 191564 462380
rect 3568 462340 3574 462352
rect 191558 462340 191564 462352
rect 191616 462340 191622 462392
rect 103422 461660 103428 461712
rect 103480 461700 103486 461712
rect 188614 461700 188620 461712
rect 103480 461672 188620 461700
rect 103480 461660 103486 461672
rect 188614 461660 188620 461672
rect 188672 461660 188678 461712
rect 81342 461592 81348 461644
rect 81400 461632 81406 461644
rect 189994 461632 190000 461644
rect 81400 461604 190000 461632
rect 81400 461592 81406 461604
rect 189994 461592 190000 461604
rect 190052 461592 190058 461644
rect 339034 461592 339040 461644
rect 339092 461632 339098 461644
rect 407114 461632 407120 461644
rect 339092 461604 407120 461632
rect 339092 461592 339098 461604
rect 407114 461592 407120 461604
rect 407172 461592 407178 461644
rect 128262 460232 128268 460284
rect 128320 460272 128326 460284
rect 183002 460272 183008 460284
rect 128320 460244 183008 460272
rect 128320 460232 128326 460244
rect 183002 460232 183008 460244
rect 183060 460232 183066 460284
rect 88242 460164 88248 460216
rect 88300 460204 88306 460216
rect 174906 460204 174912 460216
rect 88300 460176 174912 460204
rect 88300 460164 88306 460176
rect 174906 460164 174912 460176
rect 174964 460164 174970 460216
rect 118510 458872 118516 458924
rect 118568 458912 118574 458924
rect 185762 458912 185768 458924
rect 118568 458884 185768 458912
rect 118568 458872 118574 458884
rect 185762 458872 185768 458884
rect 185820 458872 185826 458924
rect 91002 458804 91008 458856
rect 91060 458844 91066 458856
rect 176378 458844 176384 458856
rect 91060 458816 176384 458844
rect 91060 458804 91066 458816
rect 176378 458804 176384 458816
rect 176436 458804 176442 458856
rect 195054 457716 195060 457768
rect 195112 457756 195118 457768
rect 195514 457756 195520 457768
rect 195112 457728 195520 457756
rect 195112 457716 195118 457728
rect 195514 457716 195520 457728
rect 195572 457716 195578 457768
rect 195238 457580 195244 457632
rect 195296 457620 195302 457632
rect 195514 457620 195520 457632
rect 195296 457592 195520 457620
rect 195296 457580 195302 457592
rect 195514 457580 195520 457592
rect 195572 457580 195578 457632
rect 125502 457512 125508 457564
rect 125560 457552 125566 457564
rect 168282 457552 168288 457564
rect 125560 457524 168288 457552
rect 125560 457512 125566 457524
rect 168282 457512 168288 457524
rect 168340 457512 168346 457564
rect 99282 457444 99288 457496
rect 99340 457484 99346 457496
rect 181806 457484 181812 457496
rect 99340 457456 181812 457484
rect 99340 457444 99346 457456
rect 181806 457444 181812 457456
rect 181864 457444 181870 457496
rect 561030 456764 561036 456816
rect 561088 456804 561094 456816
rect 580166 456804 580172 456816
rect 561088 456776 580172 456804
rect 561088 456764 561094 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 135162 456696 135168 456748
rect 135220 456736 135226 456748
rect 168742 456736 168748 456748
rect 135220 456708 168748 456736
rect 135220 456696 135226 456708
rect 168742 456696 168748 456708
rect 168800 456696 168806 456748
rect 197078 456152 197084 456204
rect 197136 456152 197142 456204
rect 137922 456084 137928 456136
rect 137980 456124 137986 456136
rect 172422 456124 172428 456136
rect 137980 456096 172428 456124
rect 137980 456084 137986 456096
rect 172422 456084 172428 456096
rect 172480 456084 172486 456136
rect 63402 456016 63408 456068
rect 63460 456056 63466 456068
rect 188706 456056 188712 456068
rect 63460 456028 188712 456056
rect 63460 456016 63466 456028
rect 188706 456016 188712 456028
rect 188764 456016 188770 456068
rect 197096 455988 197124 456152
rect 197170 455988 197176 456000
rect 197096 455960 197176 455988
rect 197170 455948 197176 455960
rect 197228 455948 197234 456000
rect 171870 455472 171876 455524
rect 171928 455512 171934 455524
rect 172422 455512 172428 455524
rect 171928 455484 172428 455512
rect 171928 455472 171934 455484
rect 172422 455472 172428 455484
rect 172480 455512 172486 455524
rect 195238 455512 195244 455524
rect 172480 455484 195244 455512
rect 172480 455472 172486 455484
rect 195238 455472 195244 455484
rect 195296 455472 195302 455524
rect 168742 455404 168748 455456
rect 168800 455444 168806 455456
rect 196066 455444 196072 455456
rect 168800 455416 196072 455444
rect 168800 455404 168806 455416
rect 196066 455404 196072 455416
rect 196124 455404 196130 455456
rect 169846 455336 169852 455388
rect 169904 455376 169910 455388
rect 171042 455376 171048 455388
rect 169904 455348 171048 455376
rect 169904 455336 169910 455348
rect 171042 455336 171048 455348
rect 171100 455376 171106 455388
rect 171594 455376 171600 455388
rect 171100 455348 171600 455376
rect 171100 455336 171106 455348
rect 171594 455336 171600 455348
rect 171652 455336 171658 455388
rect 150342 454928 150348 454980
rect 150400 454968 150406 454980
rect 169846 454968 169852 454980
rect 150400 454940 169852 454968
rect 150400 454928 150406 454940
rect 169846 454928 169852 454940
rect 169904 454928 169910 454980
rect 148318 454860 148324 454912
rect 148376 454900 148382 454912
rect 183462 454900 183468 454912
rect 148376 454872 183468 454900
rect 148376 454860 148382 454872
rect 183462 454860 183468 454872
rect 183520 454860 183526 454912
rect 113082 454792 113088 454844
rect 113140 454832 113146 454844
rect 172422 454832 172428 454844
rect 113140 454804 172428 454832
rect 113140 454792 113146 454804
rect 172422 454792 172428 454804
rect 172480 454792 172486 454844
rect 114370 454724 114376 454776
rect 114428 454764 114434 454776
rect 176102 454764 176108 454776
rect 114428 454736 176108 454764
rect 114428 454724 114434 454736
rect 176102 454724 176108 454736
rect 176160 454724 176166 454776
rect 71682 454656 71688 454708
rect 71740 454696 71746 454708
rect 184750 454696 184756 454708
rect 71740 454668 184756 454696
rect 71740 454656 71746 454668
rect 184750 454656 184756 454668
rect 184808 454656 184814 454708
rect 183186 454180 183192 454232
rect 183244 454220 183250 454232
rect 183462 454220 183468 454232
rect 183244 454192 183468 454220
rect 183244 454180 183250 454192
rect 183462 454180 183468 454192
rect 183520 454220 183526 454232
rect 197354 454220 197360 454232
rect 183520 454192 197360 454220
rect 183520 454180 183526 454192
rect 197354 454180 197360 454192
rect 197412 454180 197418 454232
rect 176102 454112 176108 454164
rect 176160 454152 176166 454164
rect 198734 454152 198740 454164
rect 176160 454124 198740 454152
rect 176160 454112 176166 454124
rect 198734 454112 198740 454124
rect 198792 454112 198798 454164
rect 172054 454044 172060 454096
rect 172112 454084 172118 454096
rect 172422 454084 172428 454096
rect 172112 454056 172428 454084
rect 172112 454044 172118 454056
rect 172422 454044 172428 454056
rect 172480 454084 172486 454096
rect 195974 454084 195980 454096
rect 172480 454056 195980 454084
rect 172480 454044 172486 454056
rect 195974 454044 195980 454056
rect 196032 454044 196038 454096
rect 193582 453976 193588 454028
rect 193640 454016 193646 454028
rect 193858 454016 193864 454028
rect 193640 453988 193864 454016
rect 193640 453976 193646 453988
rect 193858 453976 193864 453988
rect 193916 453976 193922 454028
rect 143442 453908 143448 453960
rect 143500 453948 143506 453960
rect 176010 453948 176016 453960
rect 143500 453920 176016 453948
rect 143500 453908 143506 453920
rect 176010 453908 176016 453920
rect 176068 453908 176074 453960
rect 128998 453840 129004 453892
rect 129056 453880 129062 453892
rect 172698 453880 172704 453892
rect 129056 453852 172704 453880
rect 129056 453840 129062 453852
rect 172698 453840 172704 453852
rect 172756 453840 172762 453892
rect 336274 453840 336280 453892
rect 336332 453880 336338 453892
rect 336918 453880 336924 453892
rect 336332 453852 336924 453880
rect 336332 453840 336338 453852
rect 336918 453840 336924 453852
rect 336976 453840 336982 453892
rect 126238 453772 126244 453824
rect 126296 453812 126302 453824
rect 173434 453812 173440 453824
rect 126296 453784 173440 453812
rect 126296 453772 126302 453784
rect 173434 453772 173440 453784
rect 173492 453772 173498 453824
rect 122742 453704 122748 453756
rect 122800 453744 122806 453756
rect 169846 453744 169852 453756
rect 122800 453716 169852 453744
rect 122800 453704 122806 453716
rect 169846 453704 169852 453716
rect 169904 453704 169910 453756
rect 291010 453704 291016 453756
rect 291068 453744 291074 453756
rect 338666 453744 338672 453756
rect 291068 453716 338672 453744
rect 291068 453704 291074 453716
rect 338666 453704 338672 453716
rect 338724 453704 338730 453756
rect 124122 453636 124128 453688
rect 124180 453676 124186 453688
rect 179414 453676 179420 453688
rect 124180 453648 179420 453676
rect 124180 453636 124186 453648
rect 179414 453636 179420 453648
rect 179472 453636 179478 453688
rect 289814 453636 289820 453688
rect 289872 453676 289878 453688
rect 338758 453676 338764 453688
rect 289872 453648 338764 453676
rect 289872 453636 289878 453648
rect 338758 453636 338764 453648
rect 338816 453636 338822 453688
rect 117222 453568 117228 453620
rect 117280 453608 117286 453620
rect 174078 453608 174084 453620
rect 117280 453580 174084 453608
rect 117280 453568 117286 453580
rect 174078 453568 174084 453580
rect 174136 453568 174142 453620
rect 324958 453568 324964 453620
rect 325016 453608 325022 453620
rect 399938 453608 399944 453620
rect 325016 453580 399944 453608
rect 325016 453568 325022 453580
rect 399938 453568 399944 453580
rect 399996 453568 400002 453620
rect 132402 453500 132408 453552
rect 132460 453540 132466 453552
rect 191098 453540 191104 453552
rect 132460 453512 191104 453540
rect 132460 453500 132466 453512
rect 191098 453500 191104 453512
rect 191156 453540 191162 453552
rect 278038 453540 278044 453552
rect 191156 453512 278044 453540
rect 191156 453500 191162 453512
rect 278038 453500 278044 453512
rect 278096 453500 278102 453552
rect 311158 453500 311164 453552
rect 311216 453540 311222 453552
rect 405274 453540 405280 453552
rect 311216 453512 405280 453540
rect 311216 453500 311222 453512
rect 405274 453500 405280 453512
rect 405332 453500 405338 453552
rect 114462 453432 114468 453484
rect 114520 453472 114526 453484
rect 174538 453472 174544 453484
rect 114520 453444 174544 453472
rect 114520 453432 114526 453444
rect 174538 453432 174544 453444
rect 174596 453432 174602 453484
rect 281442 453472 281448 453484
rect 190426 453444 281448 453472
rect 118602 453364 118608 453416
rect 118660 453404 118666 453416
rect 185946 453404 185952 453416
rect 118660 453376 185952 453404
rect 118660 453364 118666 453376
rect 185946 453364 185952 453376
rect 186004 453404 186010 453416
rect 190426 453404 190454 453444
rect 281442 453432 281448 453444
rect 281500 453432 281506 453484
rect 301222 453432 301228 453484
rect 301280 453472 301286 453484
rect 406562 453472 406568 453484
rect 301280 453444 406568 453472
rect 301280 453432 301286 453444
rect 406562 453432 406568 453444
rect 406620 453432 406626 453484
rect 186004 453376 190454 453404
rect 186004 453364 186010 453376
rect 196158 453364 196164 453416
rect 196216 453404 196222 453416
rect 294782 453404 294788 453416
rect 196216 453376 294788 453404
rect 196216 453364 196222 453376
rect 294782 453364 294788 453376
rect 294840 453364 294846 453416
rect 298554 453364 298560 453416
rect 298612 453404 298618 453416
rect 405642 453404 405648 453416
rect 298612 453376 405648 453404
rect 298612 453364 298618 453376
rect 405642 453364 405648 453376
rect 405700 453364 405706 453416
rect 119982 453296 119988 453348
rect 120040 453336 120046 453348
rect 189718 453336 189724 453348
rect 120040 453308 189724 453336
rect 120040 453296 120046 453308
rect 189718 453296 189724 453308
rect 189776 453336 189782 453348
rect 288894 453336 288900 453348
rect 189776 453308 288900 453336
rect 189776 453296 189782 453308
rect 288894 453296 288900 453308
rect 288952 453296 288958 453348
rect 299842 453296 299848 453348
rect 299900 453336 299906 453348
rect 409506 453336 409512 453348
rect 299900 453308 409512 453336
rect 299900 453296 299906 453308
rect 409506 453296 409512 453308
rect 409564 453296 409570 453348
rect 409690 453296 409696 453348
rect 409748 453336 409754 453348
rect 468294 453336 468300 453348
rect 409748 453308 468300 453336
rect 409748 453296 409754 453308
rect 468294 453296 468300 453308
rect 468352 453296 468358 453348
rect 199286 453228 199292 453280
rect 199344 453268 199350 453280
rect 298462 453268 298468 453280
rect 199344 453240 298468 453268
rect 199344 453228 199350 453240
rect 298462 453228 298468 453240
rect 298520 453228 298526 453280
rect 193582 453160 193588 453212
rect 193640 453200 193646 453212
rect 299566 453200 299572 453212
rect 193640 453172 299572 453200
rect 193640 453160 193646 453172
rect 299566 453160 299572 453172
rect 299624 453160 299630 453212
rect 174538 453092 174544 453144
rect 174596 453132 174602 453144
rect 284294 453132 284300 453144
rect 174596 453104 284300 453132
rect 174596 453092 174602 453104
rect 284294 453092 284300 453104
rect 284352 453092 284358 453144
rect 199194 453024 199200 453076
rect 199252 453064 199258 453076
rect 311066 453064 311072 453076
rect 199252 453036 311072 453064
rect 199252 453024 199258 453036
rect 311066 453024 311072 453036
rect 311124 453024 311130 453076
rect 174078 452956 174084 453008
rect 174136 452996 174142 453008
rect 286778 452996 286784 453008
rect 174136 452968 286784 452996
rect 174136 452956 174142 452968
rect 286778 452956 286784 452968
rect 286836 452956 286842 453008
rect 179414 452888 179420 452940
rect 179472 452928 179478 452940
rect 293678 452928 293684 452940
rect 179472 452900 293684 452928
rect 179472 452888 179478 452900
rect 293678 452888 293684 452900
rect 293736 452888 293742 452940
rect 172698 452820 172704 452872
rect 172756 452860 172762 452872
rect 290182 452860 290188 452872
rect 172756 452832 290188 452860
rect 172756 452820 172762 452832
rect 290182 452820 290188 452832
rect 290240 452820 290246 452872
rect 173434 452752 173440 452804
rect 173492 452792 173498 452804
rect 291194 452792 291200 452804
rect 173492 452764 291200 452792
rect 173492 452752 173498 452764
rect 291194 452752 291200 452764
rect 291252 452752 291258 452804
rect 169846 452684 169852 452736
rect 169904 452724 169910 452736
rect 170674 452724 170680 452736
rect 169904 452696 170680 452724
rect 169904 452684 169910 452696
rect 170674 452684 170680 452696
rect 170732 452724 170738 452736
rect 292574 452724 292580 452736
rect 170732 452696 292580 452724
rect 170732 452684 170738 452696
rect 292574 452684 292580 452696
rect 292632 452684 292638 452736
rect 335078 452684 335084 452736
rect 335136 452724 335142 452736
rect 337378 452724 337384 452736
rect 335136 452696 337384 452724
rect 335136 452684 335142 452696
rect 337378 452684 337384 452696
rect 337436 452684 337442 452736
rect 176010 452616 176016 452668
rect 176068 452656 176074 452668
rect 312354 452656 312360 452668
rect 176068 452628 312360 452656
rect 176068 452616 176074 452628
rect 312354 452616 312360 452628
rect 312412 452616 312418 452668
rect 29546 452548 29552 452600
rect 29604 452588 29610 452600
rect 29730 452588 29736 452600
rect 29604 452560 29736 452588
rect 29604 452548 29610 452560
rect 29730 452548 29736 452560
rect 29788 452548 29794 452600
rect 140682 452548 140688 452600
rect 140740 452588 140746 452600
rect 167270 452588 167276 452600
rect 140740 452560 167276 452588
rect 140740 452548 140746 452560
rect 167270 452548 167276 452560
rect 167328 452548 167334 452600
rect 176470 452548 176476 452600
rect 176528 452588 176534 452600
rect 305270 452588 305276 452600
rect 176528 452560 305276 452588
rect 176528 452548 176534 452560
rect 305270 452548 305276 452560
rect 305328 452548 305334 452600
rect 195514 452480 195520 452532
rect 195572 452520 195578 452532
rect 313366 452520 313372 452532
rect 195572 452492 313372 452520
rect 195572 452480 195578 452492
rect 313366 452480 313372 452492
rect 313424 452480 313430 452532
rect 330018 452480 330024 452532
rect 330076 452520 330082 452532
rect 399846 452520 399852 452532
rect 330076 452492 399852 452520
rect 330076 452480 330082 452492
rect 399846 452480 399852 452492
rect 399904 452480 399910 452532
rect 466178 452480 466184 452532
rect 466236 452520 466242 452532
rect 467098 452520 467104 452532
rect 466236 452492 467104 452520
rect 466236 452480 466242 452492
rect 467098 452480 467104 452492
rect 467156 452480 467162 452532
rect 473538 452480 473544 452532
rect 473596 452520 473602 452532
rect 476758 452520 476764 452532
rect 473596 452492 476764 452520
rect 473596 452480 473602 452492
rect 476758 452480 476764 452492
rect 476816 452480 476822 452532
rect 481082 452480 481088 452532
rect 481140 452520 481146 452532
rect 485130 452520 485136 452532
rect 481140 452492 485136 452520
rect 481140 452480 481146 452492
rect 485130 452480 485136 452492
rect 485188 452480 485194 452532
rect 493594 452480 493600 452532
rect 493652 452520 493658 452532
rect 497458 452520 497464 452532
rect 493652 452492 497464 452520
rect 493652 452480 493658 452492
rect 497458 452480 497464 452492
rect 497516 452480 497522 452532
rect 503530 452480 503536 452532
rect 503588 452520 503594 452532
rect 504358 452520 504364 452532
rect 503588 452492 504364 452520
rect 503588 452480 503594 452492
rect 504358 452480 504364 452492
rect 504416 452480 504422 452532
rect 505922 452480 505928 452532
rect 505980 452520 505986 452532
rect 507118 452520 507124 452532
rect 505980 452492 507124 452520
rect 505980 452480 505986 452492
rect 507118 452480 507124 452492
rect 507176 452480 507182 452532
rect 197354 452412 197360 452464
rect 197412 452452 197418 452464
rect 314654 452452 314660 452464
rect 197412 452424 314660 452452
rect 197412 452412 197418 452424
rect 314654 452412 314660 452424
rect 314712 452412 314718 452464
rect 317414 452412 317420 452464
rect 317472 452452 317478 452464
rect 399754 452452 399760 452464
rect 317472 452424 399760 452452
rect 317472 452412 317478 452424
rect 399754 452412 399760 452424
rect 399812 452412 399818 452464
rect 483474 452412 483480 452464
rect 483532 452452 483538 452464
rect 487798 452452 487804 452464
rect 483532 452424 487804 452452
rect 483532 452412 483538 452424
rect 487798 452412 487804 452424
rect 487856 452412 487862 452464
rect 195238 452344 195244 452396
rect 195296 452384 195302 452396
rect 307846 452384 307852 452396
rect 195296 452356 307852 452384
rect 195296 452344 195302 452356
rect 307846 452344 307852 452356
rect 307904 452344 307910 452396
rect 316218 452344 316224 452396
rect 316276 452384 316282 452396
rect 402606 452384 402612 452396
rect 316276 452356 402612 452384
rect 316276 452344 316282 452356
rect 402606 452344 402612 452356
rect 402664 452344 402670 452396
rect 196066 452276 196072 452328
rect 196124 452316 196130 452328
rect 304166 452316 304172 452328
rect 196124 452288 304172 452316
rect 196124 452276 196130 452288
rect 304166 452276 304172 452288
rect 304224 452276 304230 452328
rect 312446 452276 312452 452328
rect 312504 452316 312510 452328
rect 402330 452316 402336 452328
rect 312504 452288 402336 452316
rect 312504 452276 312510 452288
rect 402330 452276 402336 452288
rect 402388 452276 402394 452328
rect 151722 452208 151728 452260
rect 151780 452248 151786 452260
rect 169938 452248 169944 452260
rect 151780 452220 169944 452248
rect 151780 452208 151786 452220
rect 169938 452208 169944 452220
rect 169996 452208 170002 452260
rect 195974 452208 195980 452260
rect 196032 452248 196038 452260
rect 282086 452248 282092 452260
rect 196032 452220 282092 452248
rect 196032 452208 196038 452220
rect 282086 452208 282092 452220
rect 282144 452208 282150 452260
rect 309962 452208 309968 452260
rect 310020 452248 310026 452260
rect 402698 452248 402704 452260
rect 310020 452220 402704 452248
rect 310020 452208 310026 452220
rect 402698 452208 402704 452220
rect 402756 452208 402762 452260
rect 139210 452140 139216 452192
rect 139268 452180 139274 452192
rect 171962 452180 171968 452192
rect 139268 452152 171968 452180
rect 139268 452140 139274 452152
rect 171962 452140 171968 452152
rect 172020 452140 172026 452192
rect 198734 452140 198740 452192
rect 198792 452180 198798 452192
rect 283190 452180 283196 452192
rect 198792 452152 283196 452180
rect 198792 452140 198798 452152
rect 283190 452140 283196 452152
rect 283248 452140 283254 452192
rect 308674 452140 308680 452192
rect 308732 452180 308738 452192
rect 402422 452180 402428 452192
rect 308732 452152 402428 452180
rect 308732 452140 308738 452152
rect 402422 452140 402428 452152
rect 402480 452140 402486 452192
rect 137278 452072 137284 452124
rect 137336 452112 137342 452124
rect 170490 452112 170496 452124
rect 137336 452084 170496 452112
rect 137336 452072 137342 452084
rect 170490 452072 170496 452084
rect 170548 452072 170554 452124
rect 278038 452072 278044 452124
rect 278096 452112 278102 452124
rect 301958 452112 301964 452124
rect 278096 452084 301964 452112
rect 278096 452072 278102 452084
rect 301958 452072 301964 452084
rect 302016 452072 302022 452124
rect 306098 452072 306104 452124
rect 306156 452112 306162 452124
rect 402238 452112 402244 452124
rect 306156 452084 402244 452112
rect 306156 452072 306162 452084
rect 402238 452072 402244 452084
rect 402296 452072 402302 452124
rect 133782 452004 133788 452056
rect 133840 452044 133846 452056
rect 187050 452044 187056 452056
rect 133840 452016 187056 452044
rect 133840 452004 133846 452016
rect 187050 452004 187056 452016
rect 187108 452004 187114 452056
rect 303614 452004 303620 452056
rect 303672 452044 303678 452056
rect 402514 452044 402520 452056
rect 303672 452016 402520 452044
rect 303672 452004 303678 452016
rect 402514 452004 402520 452016
rect 402572 452004 402578 452056
rect 28534 451936 28540 451988
rect 28592 451976 28598 451988
rect 34514 451976 34520 451988
rect 28592 451948 34520 451976
rect 28592 451936 28598 451948
rect 34514 451936 34520 451948
rect 34572 451936 34578 451988
rect 66162 451936 66168 451988
rect 66220 451976 66226 451988
rect 174998 451976 175004 451988
rect 66220 451948 175004 451976
rect 66220 451936 66226 451948
rect 174998 451936 175004 451948
rect 175056 451936 175062 451988
rect 302326 451936 302332 451988
rect 302384 451976 302390 451988
rect 405458 451976 405464 451988
rect 302384 451948 405464 451976
rect 302384 451936 302390 451948
rect 405458 451936 405464 451948
rect 405516 451936 405522 451988
rect 29546 451868 29552 451920
rect 29604 451908 29610 451920
rect 45646 451908 45652 451920
rect 29604 451880 45652 451908
rect 29604 451868 29610 451880
rect 45646 451868 45652 451880
rect 45704 451868 45710 451920
rect 167270 451868 167276 451920
rect 167328 451908 167334 451920
rect 309870 451908 309876 451920
rect 167328 451880 309876 451908
rect 167328 451868 167334 451880
rect 309870 451868 309876 451880
rect 309928 451868 309934 451920
rect 320174 451868 320180 451920
rect 320232 451908 320238 451920
rect 425422 451908 425428 451920
rect 320232 451880 425428 451908
rect 320232 451868 320238 451880
rect 425422 451868 425428 451880
rect 425480 451868 425486 451920
rect 280982 451800 280988 451852
rect 281040 451840 281046 451852
rect 341426 451840 341432 451852
rect 281040 451812 341432 451840
rect 281040 451800 281046 451812
rect 341426 451800 341432 451812
rect 341484 451800 341490 451852
rect 282270 451732 282276 451784
rect 282328 451772 282334 451784
rect 341518 451772 341524 451784
rect 282328 451744 341524 451772
rect 282328 451732 282334 451744
rect 341518 451732 341524 451744
rect 341576 451732 341582 451784
rect 283466 451664 283472 451716
rect 283524 451704 283530 451716
rect 339954 451704 339960 451716
rect 283524 451676 339960 451704
rect 283524 451664 283530 451676
rect 339954 451664 339960 451676
rect 340012 451664 340018 451716
rect 195054 451596 195060 451648
rect 195112 451636 195118 451648
rect 201770 451636 201776 451648
rect 195112 451608 201776 451636
rect 195112 451596 195118 451608
rect 201770 451596 201776 451608
rect 201828 451596 201834 451648
rect 198366 451528 198372 451580
rect 198424 451568 198430 451580
rect 200206 451568 200212 451580
rect 198424 451540 200212 451568
rect 198424 451528 198430 451540
rect 200206 451528 200212 451540
rect 200264 451528 200270 451580
rect 187050 451460 187056 451512
rect 187108 451500 187114 451512
rect 303062 451500 303068 451512
rect 187108 451472 303068 451500
rect 187108 451460 187114 451472
rect 303062 451460 303068 451472
rect 303120 451460 303126 451512
rect 171962 451392 171968 451444
rect 172020 451432 172026 451444
rect 308950 451432 308956 451444
rect 172020 451404 308956 451432
rect 172020 451392 172026 451404
rect 308950 451392 308956 451404
rect 309008 451392 309014 451444
rect 170490 451324 170496 451376
rect 170548 451364 170554 451376
rect 306374 451364 306380 451376
rect 170548 451336 306380 451364
rect 170548 451324 170554 451336
rect 306374 451324 306380 451336
rect 306432 451324 306438 451376
rect 318794 451324 318800 451376
rect 318852 451364 318858 451376
rect 319438 451364 319444 451376
rect 318852 451336 319444 451364
rect 318852 451324 318858 451336
rect 319438 451324 319444 451336
rect 319496 451364 319502 451376
rect 426894 451364 426900 451376
rect 319496 451336 426900 451364
rect 319496 451324 319502 451336
rect 426894 451324 426900 451336
rect 426952 451324 426958 451376
rect 495986 451324 495992 451376
rect 496044 451364 496050 451376
rect 530578 451364 530584 451376
rect 496044 451336 530584 451364
rect 496044 451324 496050 451336
rect 530578 451324 530584 451336
rect 530636 451324 530642 451376
rect 169938 451256 169944 451308
rect 169996 451296 170002 451308
rect 320174 451296 320180 451308
rect 169996 451268 320180 451296
rect 169996 451256 170002 451268
rect 320174 451256 320180 451268
rect 320232 451256 320238 451308
rect 468662 451256 468668 451308
rect 468720 451296 468726 451308
rect 473998 451296 474004 451308
rect 468720 451268 474004 451296
rect 468720 451256 468726 451268
rect 473998 451256 474004 451268
rect 474056 451256 474062 451308
rect 476022 451256 476028 451308
rect 476080 451296 476086 451308
rect 480898 451296 480904 451308
rect 476080 451268 480904 451296
rect 476080 451256 476086 451268
rect 480898 451256 480904 451268
rect 480956 451256 480962 451308
rect 29822 451188 29828 451240
rect 29880 451228 29886 451240
rect 48038 451228 48044 451240
rect 29880 451200 48044 451228
rect 29880 451188 29886 451200
rect 48038 451188 48044 451200
rect 48096 451188 48102 451240
rect 170306 451188 170312 451240
rect 170364 451228 170370 451240
rect 452838 451228 452844 451240
rect 170364 451200 452844 451228
rect 170364 451188 170370 451200
rect 452838 451188 452844 451200
rect 452896 451188 452902 451240
rect 173802 451120 173808 451172
rect 173860 451160 173866 451172
rect 450262 451160 450268 451172
rect 173860 451132 450268 451160
rect 173860 451120 173866 451132
rect 450262 451120 450268 451132
rect 450320 451120 450326 451172
rect 169294 451052 169300 451104
rect 169352 451092 169358 451104
rect 340230 451092 340236 451104
rect 169352 451064 340236 451092
rect 169352 451052 169358 451064
rect 340230 451052 340236 451064
rect 340288 451052 340294 451104
rect 194134 450916 194140 450968
rect 194192 450956 194198 450968
rect 203058 450956 203064 450968
rect 194192 450928 203064 450956
rect 194192 450916 194198 450928
rect 203058 450916 203064 450928
rect 203116 450916 203122 450968
rect 168006 450848 168012 450900
rect 168064 450888 168070 450900
rect 193674 450888 193680 450900
rect 168064 450860 193680 450888
rect 168064 450848 168070 450860
rect 193674 450848 193680 450860
rect 193732 450888 193738 450900
rect 436278 450888 436284 450900
rect 193732 450860 436284 450888
rect 193732 450848 193738 450860
rect 436278 450848 436284 450860
rect 436336 450848 436342 450900
rect 168190 450780 168196 450832
rect 168248 450820 168254 450832
rect 187326 450820 187332 450832
rect 168248 450792 187332 450820
rect 168248 450780 168254 450792
rect 187326 450780 187332 450792
rect 187384 450820 187390 450832
rect 434714 450820 434720 450832
rect 187384 450792 434720 450820
rect 187384 450780 187390 450792
rect 434714 450780 434720 450792
rect 434772 450780 434778 450832
rect 168098 450712 168104 450764
rect 168156 450752 168162 450764
rect 179230 450752 179236 450764
rect 168156 450724 179236 450752
rect 168156 450712 168162 450724
rect 179230 450712 179236 450724
rect 179288 450752 179294 450764
rect 433702 450752 433708 450764
rect 179288 450724 433708 450752
rect 179288 450712 179294 450724
rect 433702 450712 433708 450724
rect 433760 450712 433766 450764
rect 165522 450644 165528 450696
rect 165580 450684 165586 450696
rect 184566 450684 184572 450696
rect 165580 450656 184572 450684
rect 165580 450644 165586 450656
rect 184566 450644 184572 450656
rect 184624 450684 184630 450696
rect 454126 450684 454132 450696
rect 184624 450656 454132 450684
rect 184624 450644 184630 450656
rect 454126 450644 454132 450656
rect 454184 450644 454190 450696
rect 516042 450644 516048 450696
rect 516100 450684 516106 450696
rect 556338 450684 556344 450696
rect 516100 450656 556344 450684
rect 516100 450644 516106 450656
rect 556338 450644 556344 450656
rect 556396 450644 556402 450696
rect 28718 450576 28724 450628
rect 28776 450616 28782 450628
rect 429378 450616 429384 450628
rect 28776 450588 429384 450616
rect 28776 450576 28782 450588
rect 429378 450576 429384 450588
rect 429436 450576 429442 450628
rect 443638 450576 443644 450628
rect 443696 450616 443702 450628
rect 519906 450616 519912 450628
rect 443696 450588 519912 450616
rect 443696 450576 443702 450588
rect 519906 450576 519912 450588
rect 519964 450576 519970 450628
rect 18598 450508 18604 450560
rect 18656 450548 18662 450560
rect 430574 450548 430580 450560
rect 18656 450520 430580 450548
rect 18656 450508 18662 450520
rect 430574 450508 430580 450520
rect 430632 450508 430638 450560
rect 438670 450508 438676 450560
rect 438728 450548 438734 450560
rect 517330 450548 517336 450560
rect 438728 450520 517336 450548
rect 438728 450508 438734 450520
rect 517330 450508 517336 450520
rect 517388 450508 517394 450560
rect 169294 450168 169300 450220
rect 169352 450208 169358 450220
rect 169478 450208 169484 450220
rect 169352 450180 169484 450208
rect 169352 450168 169358 450180
rect 169478 450168 169484 450180
rect 169536 450168 169542 450220
rect 28350 450100 28356 450152
rect 28408 450140 28414 450152
rect 421834 450140 421840 450152
rect 28408 450112 421840 450140
rect 28408 450100 28414 450112
rect 421834 450100 421840 450112
rect 421892 450100 421898 450152
rect 28442 450032 28448 450084
rect 28500 450072 28506 450084
rect 423030 450072 423036 450084
rect 28500 450044 423036 450072
rect 28500 450032 28506 450044
rect 423030 450032 423036 450044
rect 423088 450032 423094 450084
rect 3326 449964 3332 450016
rect 3384 450004 3390 450016
rect 410518 450004 410524 450016
rect 3384 449976 410524 450004
rect 3384 449964 3390 449976
rect 410518 449964 410524 449976
rect 410576 449964 410582 450016
rect 3510 449896 3516 449948
rect 3568 449936 3574 449948
rect 413278 449936 413284 449948
rect 3568 449908 413284 449936
rect 3568 449896 3574 449908
rect 413278 449896 413284 449908
rect 413336 449896 413342 449948
rect 169018 449828 169024 449880
rect 169076 449868 169082 449880
rect 340046 449868 340052 449880
rect 169076 449840 340052 449868
rect 169076 449828 169082 449840
rect 340046 449828 340052 449840
rect 340104 449828 340110 449880
rect 171042 449760 171048 449812
rect 171100 449800 171106 449812
rect 318794 449800 318800 449812
rect 171100 449772 318800 449800
rect 171100 449760 171106 449772
rect 318794 449760 318800 449772
rect 318852 449760 318858 449812
rect 182082 449692 182088 449744
rect 182140 449732 182146 449744
rect 300118 449732 300124 449744
rect 182140 449704 300124 449732
rect 182140 449692 182146 449704
rect 300118 449692 300124 449704
rect 300176 449692 300182 449744
rect 247034 449420 247040 449472
rect 247092 449460 247098 449472
rect 338298 449460 338304 449472
rect 247092 449432 338304 449460
rect 247092 449420 247098 449432
rect 338298 449420 338304 449432
rect 338356 449420 338362 449472
rect 175182 449352 175188 449404
rect 175240 449392 175246 449404
rect 338850 449392 338856 449404
rect 175240 449364 338856 449392
rect 175240 449352 175246 449364
rect 338850 449352 338856 449364
rect 338908 449352 338914 449404
rect 396718 449352 396724 449404
rect 396776 449392 396782 449404
rect 464522 449392 464528 449404
rect 396776 449364 464528 449392
rect 396776 449352 396782 449364
rect 464522 449352 464528 449364
rect 464580 449352 464586 449404
rect 280154 449284 280160 449336
rect 280212 449324 280218 449336
rect 490926 449324 490932 449336
rect 280212 449296 490932 449324
rect 280212 449284 280218 449296
rect 490926 449284 490932 449296
rect 490984 449284 490990 449336
rect 166718 449216 166724 449268
rect 166776 449256 166782 449268
rect 424318 449256 424324 449268
rect 166776 449228 424324 449256
rect 166776 449216 166782 449228
rect 424318 449216 424324 449228
rect 424376 449216 424382 449268
rect 478414 449216 478420 449268
rect 478472 449256 478478 449268
rect 537478 449256 537484 449268
rect 478472 449228 537484 449256
rect 478472 449216 478478 449228
rect 537478 449216 537484 449228
rect 537536 449216 537542 449268
rect 169110 449148 169116 449200
rect 169168 449188 169174 449200
rect 174170 449188 174176 449200
rect 169168 449160 174176 449188
rect 169168 449148 169174 449160
rect 174170 449148 174176 449160
rect 174228 449188 174234 449200
rect 175182 449188 175188 449200
rect 174228 449160 175188 449188
rect 174228 449148 174234 449160
rect 175182 449148 175188 449160
rect 175240 449148 175246 449200
rect 243170 449148 243176 449200
rect 243228 449188 243234 449200
rect 509786 449188 509792 449200
rect 243228 449160 509792 449188
rect 243228 449148 243234 449160
rect 509786 449148 509792 449160
rect 509844 449148 509850 449200
rect 197906 448468 197912 448520
rect 197964 448508 197970 448520
rect 549714 448508 549720 448520
rect 197964 448480 549720 448508
rect 197964 448468 197970 448480
rect 549714 448468 549720 448480
rect 549772 448468 549778 448520
rect 169386 448400 169392 448452
rect 169444 448440 169450 448452
rect 340322 448440 340328 448452
rect 169444 448412 340328 448440
rect 169444 448400 169450 448412
rect 340322 448400 340328 448412
rect 340380 448400 340386 448452
rect 169294 448332 169300 448384
rect 169352 448372 169358 448384
rect 169662 448372 169668 448384
rect 169352 448344 169668 448372
rect 169352 448332 169358 448344
rect 169662 448332 169668 448344
rect 169720 448372 169726 448384
rect 339034 448372 339040 448384
rect 169720 448344 339040 448372
rect 169720 448332 169726 448344
rect 339034 448332 339040 448344
rect 339092 448332 339098 448384
rect 199378 448264 199384 448316
rect 199436 448304 199442 448316
rect 214374 448304 214380 448316
rect 199436 448276 214380 448304
rect 199436 448264 199442 448276
rect 214374 448264 214380 448276
rect 214432 448264 214438 448316
rect 199746 448196 199752 448248
rect 199804 448236 199810 448248
rect 215570 448236 215576 448248
rect 199804 448208 215576 448236
rect 199804 448196 199810 448208
rect 215570 448196 215576 448208
rect 215628 448196 215634 448248
rect 198550 448128 198556 448180
rect 198608 448168 198614 448180
rect 216858 448168 216864 448180
rect 198608 448140 216864 448168
rect 198608 448128 198614 448140
rect 216858 448128 216864 448140
rect 216916 448128 216922 448180
rect 264606 448128 264612 448180
rect 264664 448168 264670 448180
rect 337470 448168 337476 448180
rect 264664 448140 337476 448168
rect 264664 448128 264670 448140
rect 337470 448128 337476 448140
rect 337528 448128 337534 448180
rect 196710 448060 196716 448112
rect 196768 448100 196774 448112
rect 219342 448100 219348 448112
rect 196768 448072 219348 448100
rect 196768 448060 196774 448072
rect 219342 448060 219348 448072
rect 219400 448060 219406 448112
rect 322474 448060 322480 448112
rect 322532 448100 322538 448112
rect 399662 448100 399668 448112
rect 322532 448072 399668 448100
rect 322532 448060 322538 448072
rect 399662 448060 399668 448072
rect 399720 448060 399726 448112
rect 195698 447992 195704 448044
rect 195756 448032 195762 448044
rect 218146 448032 218152 448044
rect 195756 448004 218152 448032
rect 195756 447992 195762 448004
rect 218146 447992 218152 448004
rect 218204 447992 218210 448044
rect 319990 447992 319996 448044
rect 320048 448032 320054 448044
rect 399570 448032 399576 448044
rect 320048 448004 399576 448032
rect 320048 447992 320054 448004
rect 399570 447992 399576 448004
rect 399628 447992 399634 448044
rect 195790 447924 195796 447976
rect 195848 447964 195854 447976
rect 220630 447964 220636 447976
rect 195848 447936 220636 447964
rect 195848 447924 195854 447936
rect 220630 447924 220636 447936
rect 220688 447924 220694 447976
rect 252094 447924 252100 447976
rect 252152 447964 252158 447976
rect 337562 447964 337568 447976
rect 252152 447936 337568 447964
rect 252152 447924 252158 447936
rect 337562 447924 337568 447936
rect 337620 447924 337626 447976
rect 351178 447924 351184 447976
rect 351236 447964 351242 447976
rect 459554 447964 459560 447976
rect 351236 447936 459560 447964
rect 351236 447924 351242 447936
rect 459554 447924 459560 447936
rect 459612 447924 459618 447976
rect 501230 447924 501236 447976
rect 501288 447964 501294 447976
rect 548794 447964 548800 447976
rect 501288 447936 548800 447964
rect 501288 447924 501294 447936
rect 548794 447924 548800 447936
rect 548852 447924 548858 447976
rect 196986 447856 196992 447908
rect 197044 447896 197050 447908
rect 221918 447896 221924 447908
rect 197044 447868 221924 447896
rect 197044 447856 197050 447868
rect 221918 447856 221924 447868
rect 221976 447856 221982 447908
rect 296070 447856 296076 447908
rect 296128 447896 296134 447908
rect 405182 447896 405188 447908
rect 296128 447868 405188 447896
rect 296128 447856 296134 447868
rect 405182 447856 405188 447868
rect 405240 447856 405246 447908
rect 448514 447856 448520 447908
rect 448572 447896 448578 447908
rect 522390 447896 522396 447908
rect 448572 447868 522396 447896
rect 448572 447856 448578 447868
rect 522390 447856 522396 447868
rect 522448 447856 522454 447908
rect 195606 447788 195612 447840
rect 195664 447828 195670 447840
rect 223114 447828 223120 447840
rect 195664 447800 223120 447828
rect 195664 447788 195670 447800
rect 223114 447788 223120 447800
rect 223172 447788 223178 447840
rect 255682 447788 255688 447840
rect 255740 447828 255746 447840
rect 503530 447828 503536 447840
rect 255740 447800 503536 447828
rect 255740 447788 255746 447800
rect 503530 447788 503536 447800
rect 503588 447788 503594 447840
rect 198642 447720 198648 447772
rect 198700 447760 198706 447772
rect 213086 447760 213092 447772
rect 198700 447732 213092 447760
rect 198700 447720 198706 447732
rect 213086 447720 213092 447732
rect 213144 447720 213150 447772
rect 192754 447652 192760 447704
rect 192812 447692 192818 447704
rect 204254 447692 204260 447704
rect 192812 447664 204260 447692
rect 192812 447652 192818 447664
rect 204254 447652 204260 447664
rect 204312 447652 204318 447704
rect 194502 447584 194508 447636
rect 194560 447624 194566 447636
rect 205542 447624 205548 447636
rect 194560 447596 205548 447624
rect 194560 447584 194566 447596
rect 205542 447584 205548 447596
rect 205600 447584 205606 447636
rect 204530 447108 204536 447160
rect 204588 447148 204594 447160
rect 449434 447148 449440 447160
rect 204588 447120 449440 447148
rect 204588 447108 204594 447120
rect 449434 447108 449440 447120
rect 449492 447108 449498 447160
rect 244550 446564 244556 446616
rect 244608 446604 244614 446616
rect 338390 446604 338396 446616
rect 244608 446576 338396 446604
rect 244608 446564 244614 446576
rect 338390 446564 338396 446576
rect 338448 446564 338454 446616
rect 397454 446564 397460 446616
rect 397512 446604 397518 446616
rect 466454 446604 466460 446616
rect 397512 446576 466460 446604
rect 397512 446564 397518 446576
rect 466454 446564 466460 446576
rect 466512 446564 466518 446616
rect 293034 446496 293040 446548
rect 293092 446536 293098 446548
rect 436738 446536 436744 446548
rect 293092 446508 436744 446536
rect 293092 446496 293098 446508
rect 436738 446496 436744 446508
rect 436796 446496 436802 446548
rect 491018 446496 491024 446548
rect 491076 446536 491082 446548
rect 543734 446536 543740 446548
rect 491076 446508 543740 446536
rect 491076 446496 491082 446508
rect 543734 446496 543740 446508
rect 543792 446496 543798 446548
rect 273162 446428 273168 446480
rect 273220 446468 273226 446480
rect 494698 446468 494704 446480
rect 273220 446440 494704 446468
rect 273220 446428 273226 446440
rect 494698 446428 494704 446440
rect 494756 446428 494762 446480
rect 184198 446360 184204 446412
rect 184256 446400 184262 446412
rect 452010 446400 452016 446412
rect 184256 446372 452016 446400
rect 184256 446360 184262 446372
rect 452010 446360 452016 446372
rect 452068 446360 452074 446412
rect 453666 446360 453672 446412
rect 453724 446400 453730 446412
rect 524874 446400 524880 446412
rect 453724 446372 524880 446400
rect 453724 446360 453730 446372
rect 524874 446360 524880 446372
rect 524932 446360 524938 446412
rect 199838 445680 199844 445732
rect 199896 445720 199902 445732
rect 226886 445720 226892 445732
rect 199896 445692 226892 445720
rect 199896 445680 199902 445692
rect 226886 445680 226892 445692
rect 226944 445680 226950 445732
rect 268378 445680 268384 445732
rect 268436 445720 268442 445732
rect 341334 445720 341340 445732
rect 268436 445692 341340 445720
rect 268436 445680 268442 445692
rect 341334 445680 341340 445692
rect 341392 445680 341398 445732
rect 197170 445612 197176 445664
rect 197228 445652 197234 445664
rect 225690 445652 225696 445664
rect 197228 445624 225696 445652
rect 197228 445612 197234 445624
rect 225690 445612 225696 445624
rect 225748 445612 225754 445664
rect 262122 445612 262128 445664
rect 262180 445652 262186 445664
rect 339678 445652 339684 445664
rect 262180 445624 339684 445652
rect 262180 445612 262186 445624
rect 339678 445612 339684 445624
rect 339736 445612 339742 445664
rect 195882 445544 195888 445596
rect 195940 445584 195946 445596
rect 228174 445584 228180 445596
rect 195940 445556 228180 445584
rect 195940 445544 195946 445556
rect 228174 445544 228180 445556
rect 228232 445544 228238 445596
rect 260834 445544 260840 445596
rect 260892 445584 260898 445596
rect 339770 445584 339776 445596
rect 260892 445556 339776 445584
rect 260892 445544 260898 445556
rect 339770 445544 339776 445556
rect 339828 445544 339834 445596
rect 198458 445476 198464 445528
rect 198516 445516 198522 445528
rect 230658 445516 230664 445528
rect 198516 445488 230664 445516
rect 198516 445476 198522 445488
rect 230658 445476 230664 445488
rect 230716 445476 230722 445528
rect 259638 445476 259644 445528
rect 259696 445516 259702 445528
rect 339586 445516 339592 445528
rect 259696 445488 339592 445516
rect 259696 445476 259702 445488
rect 339586 445476 339592 445488
rect 339644 445476 339650 445528
rect 199562 445408 199568 445460
rect 199620 445448 199626 445460
rect 231946 445448 231952 445460
rect 199620 445420 231952 445448
rect 199620 445408 199626 445420
rect 231946 445408 231952 445420
rect 232004 445408 232010 445460
rect 258350 445408 258356 445460
rect 258408 445448 258414 445460
rect 341150 445448 341156 445460
rect 258408 445420 341156 445448
rect 258408 445408 258414 445420
rect 341150 445408 341156 445420
rect 341208 445408 341214 445460
rect 196618 445340 196624 445392
rect 196676 445380 196682 445392
rect 229462 445380 229468 445392
rect 196676 445352 229468 445380
rect 196676 445340 196682 445352
rect 229462 445340 229468 445352
rect 229520 445340 229526 445392
rect 253290 445340 253296 445392
rect 253348 445380 253354 445392
rect 337010 445380 337016 445392
rect 253348 445352 337016 445380
rect 253348 445340 253354 445352
rect 337010 445340 337016 445352
rect 337068 445340 337074 445392
rect 199654 445272 199660 445324
rect 199712 445312 199718 445324
rect 234430 445312 234436 445324
rect 199712 445284 234436 445312
rect 199712 445272 199718 445284
rect 234430 445272 234436 445284
rect 234488 445272 234494 445324
rect 254578 445272 254584 445324
rect 254636 445312 254642 445324
rect 338482 445312 338488 445324
rect 254636 445284 338488 445312
rect 254636 445272 254642 445284
rect 338482 445272 338488 445284
rect 338540 445272 338546 445324
rect 199470 445204 199476 445256
rect 199528 445244 199534 445256
rect 233234 445244 233240 445256
rect 199528 445216 233240 445244
rect 199528 445204 199534 445216
rect 233234 445204 233240 445216
rect 233292 445204 233298 445256
rect 257062 445204 257068 445256
rect 257120 445244 257126 445256
rect 341058 445244 341064 445256
rect 257120 445216 341064 445244
rect 257120 445204 257126 445216
rect 341058 445204 341064 445216
rect 341116 445204 341122 445256
rect 192846 445136 192852 445188
rect 192904 445176 192910 445188
rect 235718 445176 235724 445188
rect 192904 445148 235724 445176
rect 192904 445136 192910 445148
rect 235718 445136 235724 445148
rect 235776 445136 235782 445188
rect 255866 445136 255872 445188
rect 255924 445176 255930 445188
rect 341242 445176 341248 445188
rect 255924 445148 341248 445176
rect 255924 445136 255930 445148
rect 341242 445136 341248 445148
rect 341300 445136 341306 445188
rect 194226 445068 194232 445120
rect 194284 445108 194290 445120
rect 237006 445108 237012 445120
rect 194284 445080 237012 445108
rect 194284 445068 194290 445080
rect 237006 445068 237012 445080
rect 237064 445068 237070 445120
rect 243262 445068 243268 445120
rect 243320 445108 243326 445120
rect 338206 445108 338212 445120
rect 243320 445080 338212 445108
rect 243320 445068 243326 445080
rect 338206 445068 338212 445080
rect 338264 445068 338270 445120
rect 344278 445068 344284 445120
rect 344336 445108 344342 445120
rect 460750 445108 460756 445120
rect 344336 445080 460756 445108
rect 344336 445068 344342 445080
rect 460750 445068 460756 445080
rect 460808 445068 460814 445120
rect 463602 445068 463608 445120
rect 463660 445108 463666 445120
rect 529934 445108 529940 445120
rect 463660 445080 529940 445108
rect 463660 445068 463666 445080
rect 529934 445068 529940 445080
rect 529992 445068 529998 445120
rect 191650 445000 191656 445052
rect 191708 445040 191714 445052
rect 238202 445040 238208 445052
rect 191708 445012 238208 445040
rect 191708 445000 191714 445012
rect 238202 445000 238208 445012
rect 238260 445000 238266 445052
rect 265618 445000 265624 445052
rect 265676 445040 265682 445052
rect 498470 445040 498476 445052
rect 265676 445012 498476 445040
rect 265676 445000 265682 445012
rect 498470 445000 498476 445012
rect 498528 445000 498534 445052
rect 197078 444932 197084 444984
rect 197136 444972 197142 444984
rect 224402 444972 224408 444984
rect 197136 444944 224408 444972
rect 197136 444932 197142 444944
rect 224402 444932 224408 444944
rect 224460 444932 224466 444984
rect 269666 444932 269672 444984
rect 269724 444972 269730 444984
rect 342530 444972 342536 444984
rect 269724 444944 342536 444972
rect 269724 444932 269730 444944
rect 342530 444932 342536 444944
rect 342588 444932 342594 444984
rect 193030 444864 193036 444916
rect 193088 444904 193094 444916
rect 211798 444904 211804 444916
rect 193088 444876 211804 444904
rect 193088 444864 193094 444876
rect 211798 444864 211804 444876
rect 211856 444864 211862 444916
rect 327534 444864 327540 444916
rect 327592 444904 327598 444916
rect 399478 444904 399484 444916
rect 327592 444876 399484 444904
rect 327592 444864 327598 444876
rect 399478 444864 399484 444876
rect 399536 444864 399542 444916
rect 194410 444796 194416 444848
rect 194468 444836 194474 444848
rect 210602 444836 210608 444848
rect 194468 444808 210608 444836
rect 194468 444796 194474 444808
rect 210602 444796 210608 444808
rect 210660 444796 210666 444848
rect 270954 444796 270960 444848
rect 271012 444836 271018 444848
rect 340966 444836 340972 444848
rect 271012 444808 340972 444836
rect 271012 444796 271018 444808
rect 340966 444796 340972 444808
rect 341024 444796 341030 444848
rect 348418 443776 348424 443828
rect 348476 443816 348482 443828
rect 456978 443816 456984 443828
rect 348476 443788 456984 443816
rect 348476 443776 348482 443788
rect 456978 443776 456984 443788
rect 457036 443776 457042 443828
rect 263502 443708 263508 443760
rect 263560 443748 263566 443760
rect 499758 443748 499764 443760
rect 263560 443720 499764 443748
rect 263560 443708 263566 443720
rect 499758 443708 499764 443720
rect 499816 443708 499822 443760
rect 507118 443708 507124 443760
rect 507176 443748 507182 443760
rect 551278 443748 551284 443760
rect 507176 443720 551284 443748
rect 507176 443708 507182 443720
rect 551278 443708 551284 443720
rect 551336 443708 551342 443760
rect 178770 443640 178776 443692
rect 178828 443680 178834 443692
rect 439406 443680 439412 443692
rect 178828 443652 439412 443680
rect 178828 443640 178834 443652
rect 439406 443640 439412 443652
rect 439464 443640 439470 443692
rect 456702 443640 456708 443692
rect 456760 443680 456766 443692
rect 526162 443680 526168 443692
rect 456760 443652 526168 443680
rect 456760 443640 456766 443652
rect 526162 443640 526168 443652
rect 526220 443640 526226 443692
rect 277210 442892 277216 442944
rect 277268 442932 277274 442944
rect 337102 442932 337108 442944
rect 277268 442904 337108 442932
rect 277268 442892 277274 442904
rect 337102 442892 337108 442904
rect 337160 442892 337166 442944
rect 275922 442824 275928 442876
rect 275980 442864 275986 442876
rect 339494 442864 339500 442876
rect 275980 442836 339500 442864
rect 275980 442824 275986 442836
rect 339494 442824 339500 442836
rect 339552 442824 339558 442876
rect 274726 442756 274732 442808
rect 274784 442796 274790 442808
rect 338574 442796 338580 442808
rect 274784 442768 338580 442796
rect 274784 442756 274790 442768
rect 338574 442756 338580 442768
rect 338632 442756 338638 442808
rect 273438 442688 273444 442740
rect 273496 442728 273502 442740
rect 339862 442728 339868 442740
rect 273496 442700 339868 442728
rect 273496 442688 273502 442700
rect 339862 442688 339868 442700
rect 339920 442688 339926 442740
rect 272150 442620 272156 442672
rect 272208 442660 272214 442672
rect 340874 442660 340880 442672
rect 272208 442632 340880 442660
rect 272208 442620 272214 442632
rect 340874 442620 340880 442632
rect 340932 442620 340938 442672
rect 263410 442552 263416 442604
rect 263468 442592 263474 442604
rect 336826 442592 336832 442604
rect 263468 442564 336832 442592
rect 263468 442552 263474 442564
rect 336826 442552 336832 442564
rect 336884 442552 336890 442604
rect 267182 442484 267188 442536
rect 267240 442524 267246 442536
rect 342438 442524 342444 442536
rect 267240 442496 342444 442524
rect 267240 442484 267246 442496
rect 342438 442484 342444 442496
rect 342496 442484 342502 442536
rect 265894 442416 265900 442468
rect 265952 442456 265958 442468
rect 342346 442456 342352 442468
rect 265952 442428 342352 442456
rect 265952 442416 265958 442428
rect 342346 442416 342352 442428
rect 342404 442416 342410 442468
rect 400950 442416 400956 442468
rect 401008 442456 401014 442468
rect 434346 442456 434352 442468
rect 401008 442428 434352 442456
rect 401008 442416 401014 442428
rect 434346 442416 434352 442428
rect 434404 442416 434410 442468
rect 191742 442348 191748 442400
rect 191800 442388 191806 442400
rect 239490 442388 239496 442400
rect 191800 442360 239496 442388
rect 191800 442348 191806 442360
rect 239490 442348 239496 442360
rect 239548 442348 239554 442400
rect 278682 442348 278688 442400
rect 278740 442388 278746 442400
rect 492214 442388 492220 442400
rect 278740 442360 492220 442388
rect 278740 442348 278746 442360
rect 492214 442348 492220 442360
rect 492272 442348 492278 442400
rect 177298 442280 177304 442332
rect 177356 442320 177362 442332
rect 450722 442320 450728 442332
rect 177356 442292 450728 442320
rect 177356 442280 177362 442292
rect 450722 442280 450728 442292
rect 450780 442280 450786 442332
rect 487062 442280 487068 442332
rect 487120 442320 487126 442332
rect 541250 442320 541256 442332
rect 487120 442292 541256 442320
rect 487120 442280 487126 442292
rect 541250 442280 541256 442292
rect 541308 442280 541314 442332
rect 234522 442212 234528 442264
rect 234580 442252 234586 442264
rect 514846 442252 514852 442264
rect 234580 442224 514852 442252
rect 234580 442212 234586 442224
rect 514846 442212 514852 442224
rect 514904 442212 514910 442264
rect 278498 442144 278504 442196
rect 278556 442184 278562 442196
rect 337194 442184 337200 442196
rect 278556 442156 337200 442184
rect 278556 442144 278562 442156
rect 337194 442144 337200 442156
rect 337252 442144 337258 442196
rect 279694 442076 279700 442128
rect 279752 442116 279758 442128
rect 337286 442116 337292 442128
rect 279752 442088 337292 442116
rect 279752 442076 279758 442088
rect 337286 442076 337292 442088
rect 337344 442076 337350 442128
rect 167914 441532 167920 441584
rect 167972 441572 167978 441584
rect 442994 441572 443000 441584
rect 167972 441544 443000 441572
rect 167972 441532 167978 441544
rect 442994 441532 443000 441544
rect 443052 441532 443058 441584
rect 358078 441056 358084 441108
rect 358136 441096 358142 441108
rect 454494 441096 454500 441108
rect 358136 441068 454500 441096
rect 358136 441056 358142 441068
rect 454494 441056 454500 441068
rect 454552 441056 454558 441108
rect 285582 440988 285588 441040
rect 285640 441028 285646 441040
rect 471238 441028 471244 441040
rect 285640 441000 471244 441028
rect 285640 440988 285646 441000
rect 471238 440988 471244 441000
rect 471296 440988 471302 441040
rect 260742 440920 260748 440972
rect 260800 440960 260806 440972
rect 501046 440960 501052 440972
rect 260800 440932 501052 440960
rect 260800 440920 260806 440932
rect 501046 440920 501052 440932
rect 501104 440920 501110 440972
rect 186958 440852 186964 440904
rect 187016 440892 187022 440904
rect 448238 440892 448244 440904
rect 187016 440864 448244 440892
rect 187016 440852 187022 440864
rect 448238 440852 448244 440864
rect 448296 440852 448302 440904
rect 471882 440852 471888 440904
rect 471940 440892 471946 440904
rect 533706 440892 533712 440904
rect 471940 440864 533712 440892
rect 471940 440852 471946 440864
rect 533706 440852 533712 440864
rect 533764 440852 533770 440904
rect 167822 440172 167828 440224
rect 167880 440212 167886 440224
rect 437658 440212 437664 440224
rect 167880 440184 437664 440212
rect 167880 440172 167886 440184
rect 437658 440172 437664 440184
rect 437716 440172 437722 440224
rect 169754 440104 169760 440156
rect 169812 440144 169818 440156
rect 438946 440144 438952 440156
rect 169812 440116 438952 440144
rect 169812 440104 169818 440116
rect 438946 440104 438952 440116
rect 439004 440104 439010 440156
rect 333790 439764 333796 439816
rect 333848 439804 333854 439816
rect 409414 439804 409420 439816
rect 333848 439776 409420 439804
rect 333848 439764 333854 439776
rect 409414 439764 409420 439776
rect 409472 439764 409478 439816
rect 356698 439696 356704 439748
rect 356756 439736 356762 439748
rect 458174 439736 458180 439748
rect 356756 439708 458180 439736
rect 356756 439696 356762 439708
rect 458174 439696 458180 439708
rect 458232 439696 458238 439748
rect 187786 439628 187792 439680
rect 187844 439668 187850 439680
rect 444466 439668 444472 439680
rect 187844 439640 444472 439668
rect 187844 439628 187850 439640
rect 444466 439628 444472 439640
rect 444524 439628 444530 439680
rect 476758 439628 476764 439680
rect 476816 439668 476822 439680
rect 534994 439668 535000 439680
rect 476816 439640 535000 439668
rect 476816 439628 476822 439640
rect 534994 439628 535000 439640
rect 535052 439628 535058 439680
rect 306282 439560 306288 439612
rect 306340 439600 306346 439612
rect 478414 439600 478420 439612
rect 306340 439572 478420 439600
rect 306340 439560 306346 439572
rect 478414 439560 478420 439572
rect 478472 439560 478478 439612
rect 188338 439492 188344 439544
rect 188396 439532 188402 439544
rect 444466 439532 444472 439544
rect 188396 439504 444472 439532
rect 188396 439492 188402 439504
rect 444466 439492 444472 439504
rect 444524 439492 444530 439544
rect 447042 439492 447048 439544
rect 447100 439532 447106 439544
rect 521102 439532 521108 439544
rect 447100 439504 521108 439532
rect 447100 439492 447106 439504
rect 521102 439492 521108 439504
rect 521160 439492 521166 439544
rect 168006 438880 168012 438932
rect 168064 438920 168070 438932
rect 169754 438920 169760 438932
rect 168064 438892 169760 438920
rect 168064 438880 168070 438892
rect 169754 438880 169760 438892
rect 169812 438880 169818 438932
rect 173250 438812 173256 438864
rect 173308 438852 173314 438864
rect 187786 438852 187792 438864
rect 173308 438824 187792 438852
rect 173308 438812 173314 438824
rect 187786 438812 187792 438824
rect 187844 438812 187850 438864
rect 393958 438336 393964 438388
rect 394016 438376 394022 438388
rect 462038 438376 462044 438388
rect 394016 438348 462044 438376
rect 394016 438336 394022 438348
rect 462038 438336 462044 438348
rect 462096 438336 462102 438388
rect 288342 438268 288348 438320
rect 288400 438308 288406 438320
rect 485038 438308 485044 438320
rect 288400 438280 485044 438308
rect 288400 438268 288406 438280
rect 485038 438268 485044 438280
rect 485096 438268 485102 438320
rect 275830 438200 275836 438252
rect 275888 438240 275894 438252
rect 493502 438240 493508 438252
rect 275888 438212 493508 438240
rect 275888 438200 275894 438212
rect 493502 438200 493508 438212
rect 493560 438200 493566 438252
rect 497458 438200 497464 438252
rect 497516 438240 497522 438252
rect 545022 438240 545028 438252
rect 497516 438212 545028 438240
rect 497516 438200 497522 438212
rect 545022 438200 545028 438212
rect 545080 438200 545086 438252
rect 186958 438132 186964 438184
rect 187016 438172 187022 438184
rect 432046 438172 432052 438184
rect 187016 438144 432052 438172
rect 187016 438132 187022 438144
rect 432046 438132 432052 438144
rect 432104 438132 432110 438184
rect 459462 438132 459468 438184
rect 459520 438172 459526 438184
rect 527450 438172 527456 438184
rect 459520 438144 527456 438172
rect 459520 438132 459526 438144
rect 527450 438132 527456 438144
rect 527508 438132 527514 438184
rect 314930 436840 314936 436892
rect 314988 436880 314994 436892
rect 409230 436880 409236 436892
rect 314988 436852 409236 436880
rect 314988 436840 314994 436852
rect 409230 436840 409236 436852
rect 409288 436840 409294 436892
rect 485130 436840 485136 436892
rect 485188 436880 485194 436892
rect 538766 436880 538772 436892
rect 485188 436852 538772 436880
rect 485188 436840 485194 436852
rect 538766 436840 538772 436852
rect 538824 436840 538830 436892
rect 284202 436772 284208 436824
rect 284260 436812 284266 436824
rect 489730 436812 489736 436824
rect 284260 436784 489736 436812
rect 284260 436772 284266 436784
rect 489730 436772 489736 436784
rect 489788 436772 489794 436824
rect 248230 436704 248236 436756
rect 248288 436744 248294 436756
rect 507302 436744 507308 436756
rect 248288 436716 507308 436744
rect 248288 436704 248294 436716
rect 507302 436704 507308 436716
rect 507360 436704 507366 436756
rect 473354 435480 473360 435532
rect 473412 435520 473418 435532
rect 548518 435520 548524 435532
rect 473412 435492 548524 435520
rect 473412 435480 473418 435492
rect 548518 435480 548524 435492
rect 548576 435480 548582 435532
rect 309042 435412 309048 435464
rect 309100 435452 309106 435464
rect 477126 435452 477132 435464
rect 309100 435424 477132 435452
rect 309100 435412 309106 435424
rect 477126 435412 477132 435424
rect 477184 435412 477190 435464
rect 251082 435344 251088 435396
rect 251140 435384 251146 435396
rect 506014 435384 506020 435396
rect 251140 435356 506020 435384
rect 251140 435344 251146 435356
rect 506014 435344 506020 435356
rect 506072 435344 506078 435396
rect 191558 434052 191564 434104
rect 191616 434092 191622 434104
rect 426802 434092 426808 434104
rect 191616 434064 426808 434092
rect 191616 434052 191622 434064
rect 426802 434052 426808 434064
rect 426860 434052 426866 434104
rect 451182 434052 451188 434104
rect 451240 434092 451246 434104
rect 523678 434092 523684 434104
rect 451240 434064 523684 434092
rect 451240 434052 451246 434064
rect 523678 434052 523684 434064
rect 523736 434052 523742 434104
rect 253842 433984 253848 434036
rect 253900 434024 253906 434036
rect 504818 434024 504824 434036
rect 253900 433996 504824 434024
rect 253900 433984 253906 433996
rect 504818 433984 504824 433996
rect 504876 433984 504882 434036
rect 511902 433984 511908 434036
rect 511960 434024 511966 434036
rect 553854 434024 553860 434036
rect 511960 433996 553860 434024
rect 511960 433984 511966 433996
rect 553854 433984 553860 433996
rect 553912 433984 553918 434036
rect 326246 432692 326252 432744
rect 326304 432732 326310 432744
rect 398098 432732 398104 432744
rect 326304 432704 398104 432732
rect 326304 432692 326310 432704
rect 398098 432692 398104 432704
rect 398156 432692 398162 432744
rect 292298 432624 292304 432676
rect 292356 432664 292362 432676
rect 409322 432664 409328 432676
rect 292356 432636 409328 432664
rect 292356 432624 292362 432636
rect 409322 432624 409328 432636
rect 409380 432624 409386 432676
rect 467098 432624 467104 432676
rect 467156 432664 467162 432676
rect 531222 432664 531228 432676
rect 467156 432636 531228 432664
rect 467156 432624 467162 432636
rect 531222 432624 531228 432636
rect 531280 432624 531286 432676
rect 245562 432556 245568 432608
rect 245620 432596 245626 432608
rect 508590 432596 508596 432608
rect 245620 432568 508596 432596
rect 245620 432556 245626 432568
rect 508590 432556 508596 432568
rect 508648 432556 508654 432608
rect 331306 431536 331312 431588
rect 331364 431576 331370 431588
rect 340138 431576 340144 431588
rect 331364 431548 340144 431576
rect 331364 431536 331370 431548
rect 340138 431536 340144 431548
rect 340196 431536 340202 431588
rect 241974 431468 241980 431520
rect 242032 431508 242038 431520
rect 336734 431508 336740 431520
rect 242032 431480 336740 431508
rect 242032 431468 242038 431480
rect 336734 431468 336740 431480
rect 336792 431468 336798 431520
rect 353938 431468 353944 431520
rect 353996 431508 354002 431520
rect 455782 431508 455788 431520
rect 353996 431480 455788 431508
rect 353996 431468 354002 431480
rect 455782 431468 455788 431480
rect 455840 431468 455846 431520
rect 462222 431468 462228 431520
rect 462280 431508 462286 431520
rect 528646 431508 528652 431520
rect 462280 431480 528652 431508
rect 462280 431468 462286 431480
rect 528646 431468 528652 431480
rect 528704 431468 528710 431520
rect 259362 431400 259368 431452
rect 259420 431440 259426 431452
rect 502242 431440 502248 431452
rect 259420 431412 502248 431440
rect 259420 431400 259426 431412
rect 502242 431400 502248 431412
rect 502300 431400 502306 431452
rect 198550 431332 198556 431384
rect 198608 431372 198614 431384
rect 465074 431372 465080 431384
rect 198608 431344 465080 431372
rect 198608 431332 198614 431344
rect 465074 431332 465080 431344
rect 465132 431332 465138 431384
rect 199194 431264 199200 431316
rect 199252 431304 199258 431316
rect 468018 431304 468024 431316
rect 199252 431276 468024 431304
rect 199252 431264 199258 431276
rect 468018 431264 468024 431276
rect 468076 431264 468082 431316
rect 198366 431196 198372 431248
rect 198424 431236 198430 431248
rect 467926 431236 467932 431248
rect 198424 431208 467932 431236
rect 198424 431196 198430 431208
rect 467926 431196 467932 431208
rect 467984 431196 467990 431248
rect 567930 430584 567936 430636
rect 567988 430624 567994 430636
rect 579890 430624 579896 430636
rect 567988 430596 579896 430624
rect 567988 430584 567994 430596
rect 579890 430584 579896 430596
rect 579948 430584 579954 430636
rect 323762 430244 323768 430296
rect 323820 430284 323826 430296
rect 391198 430284 391204 430296
rect 323820 430256 391204 430284
rect 323820 430244 323826 430256
rect 391198 430244 391204 430256
rect 391256 430244 391262 430296
rect 404998 430244 405004 430296
rect 405056 430284 405062 430296
rect 463326 430284 463332 430296
rect 405056 430256 463332 430284
rect 405056 430244 405062 430256
rect 463326 430244 463332 430256
rect 463384 430244 463390 430296
rect 291102 430176 291108 430228
rect 291160 430216 291166 430228
rect 447778 430216 447784 430228
rect 291160 430188 447784 430216
rect 291160 430176 291166 430188
rect 447778 430176 447784 430188
rect 447836 430176 447842 430228
rect 198734 430108 198740 430160
rect 198792 430148 198798 430160
rect 459738 430148 459744 430160
rect 198792 430120 459744 430148
rect 198792 430108 198798 430120
rect 459738 430108 459744 430120
rect 459796 430108 459802 430160
rect 198918 430040 198924 430092
rect 198976 430080 198982 430092
rect 461026 430080 461032 430092
rect 198976 430052 461032 430080
rect 198976 430040 198982 430052
rect 461026 430040 461032 430052
rect 461084 430040 461090 430092
rect 199010 429972 199016 430024
rect 199068 430012 199074 430024
rect 462406 430012 462412 430024
rect 199068 429984 462412 430012
rect 199068 429972 199074 429984
rect 462406 429972 462412 429984
rect 462464 429972 462470 430024
rect 198642 429904 198648 429956
rect 198700 429944 198706 429956
rect 462314 429944 462320 429956
rect 198700 429916 462320 429944
rect 198700 429904 198706 429916
rect 462314 429904 462320 429916
rect 462372 429904 462378 429956
rect 199102 429836 199108 429888
rect 199160 429876 199166 429888
rect 466546 429876 466552 429888
rect 199160 429848 466552 429876
rect 199160 429836 199166 429848
rect 466546 429836 466552 429848
rect 466604 429836 466610 429888
rect 175366 429088 175372 429140
rect 175424 429128 175430 429140
rect 451366 429128 451372 429140
rect 175424 429100 451372 429128
rect 175424 429088 175430 429100
rect 451366 429088 451372 429100
rect 451424 429088 451430 429140
rect 178034 429020 178040 429072
rect 178092 429060 178098 429072
rect 452746 429060 452752 429072
rect 178092 429032 452752 429060
rect 178092 429020 178098 429032
rect 452746 429020 452752 429032
rect 452804 429020 452810 429072
rect 170306 428952 170312 429004
rect 170364 428992 170370 429004
rect 171502 428992 171508 429004
rect 170364 428964 171508 428992
rect 170364 428952 170370 428964
rect 171502 428952 171508 428964
rect 171560 428992 171566 429004
rect 428458 428992 428464 429004
rect 171560 428964 428464 428992
rect 171560 428952 171566 428964
rect 428458 428952 428464 428964
rect 428516 428952 428522 429004
rect 303522 428680 303528 428732
rect 303580 428720 303586 428732
rect 479610 428720 479616 428732
rect 303580 428692 479616 428720
rect 303580 428680 303586 428692
rect 479610 428680 479616 428692
rect 479668 428680 479674 428732
rect 198826 428612 198832 428664
rect 198884 428652 198890 428664
rect 458266 428652 458272 428664
rect 198884 428624 458272 428652
rect 198884 428612 198890 428624
rect 458266 428612 458272 428624
rect 458324 428612 458330 428664
rect 198458 428544 198464 428596
rect 198516 428584 198522 428596
rect 463786 428584 463792 428596
rect 198516 428556 463792 428584
rect 198516 428544 198522 428556
rect 463786 428544 463792 428556
rect 463844 428544 463850 428596
rect 177850 428476 177856 428528
rect 177908 428516 177914 428528
rect 455506 428516 455512 428528
rect 177908 428488 455512 428516
rect 177908 428476 177914 428488
rect 455506 428476 455512 428488
rect 455564 428476 455570 428528
rect 178770 428408 178776 428460
rect 178828 428448 178834 428460
rect 456886 428448 456892 428460
rect 178828 428420 456892 428448
rect 178828 428408 178834 428420
rect 456886 428408 456892 428420
rect 456944 428408 456950 428460
rect 473998 428408 474004 428460
rect 474056 428448 474062 428460
rect 532418 428448 532424 428460
rect 474056 428420 532424 428448
rect 474056 428408 474062 428420
rect 532418 428408 532424 428420
rect 532476 428408 532482 428460
rect 173618 427796 173624 427848
rect 173676 427836 173682 427848
rect 175366 427836 175372 427848
rect 173676 427808 175372 427836
rect 173676 427796 173682 427808
rect 175366 427796 175372 427808
rect 175424 427796 175430 427848
rect 177298 427796 177304 427848
rect 177356 427836 177362 427848
rect 178034 427836 178040 427848
rect 177356 427808 178040 427836
rect 177356 427796 177362 427808
rect 178034 427796 178040 427808
rect 178092 427796 178098 427848
rect 173710 427728 173716 427780
rect 173768 427768 173774 427780
rect 445846 427768 445852 427780
rect 173768 427740 445852 427768
rect 173768 427728 173774 427740
rect 445846 427728 445852 427740
rect 445904 427728 445910 427780
rect 180334 427660 180340 427712
rect 180392 427700 180398 427712
rect 180794 427700 180800 427712
rect 180392 427672 180800 427700
rect 180392 427660 180398 427672
rect 180794 427660 180800 427672
rect 180852 427700 180858 427712
rect 447226 427700 447232 427712
rect 180852 427672 447232 427700
rect 180852 427660 180858 427672
rect 447226 427660 447232 427672
rect 447284 427660 447290 427712
rect 172146 427592 172152 427644
rect 172204 427632 172210 427644
rect 198826 427632 198832 427644
rect 172204 427604 198832 427632
rect 172204 427592 172210 427604
rect 198826 427592 198832 427604
rect 198884 427592 198890 427644
rect 304902 427116 304908 427168
rect 304960 427156 304966 427168
rect 409138 427156 409144 427168
rect 304960 427128 409144 427156
rect 304960 427116 304966 427128
rect 409138 427116 409144 427128
rect 409196 427116 409202 427168
rect 441522 427116 441528 427168
rect 441580 427156 441586 427168
rect 518618 427156 518624 427168
rect 441580 427128 518624 427156
rect 441580 427116 441586 427128
rect 518618 427116 518624 427128
rect 518676 427116 518682 427168
rect 191742 427048 191748 427100
rect 191800 427088 191806 427100
rect 448606 427088 448612 427100
rect 191800 427060 448612 427088
rect 191800 427048 191806 427060
rect 448606 427048 448612 427060
rect 448664 427048 448670 427100
rect 488442 427048 488448 427100
rect 488500 427088 488506 427100
rect 542538 427088 542544 427100
rect 488500 427060 542544 427088
rect 488500 427048 488506 427060
rect 542538 427048 542544 427060
rect 542596 427048 542602 427100
rect 184198 426436 184204 426488
rect 184256 426476 184262 426488
rect 392854 426476 392860 426488
rect 184256 426448 392860 426476
rect 184256 426436 184262 426448
rect 392854 426436 392860 426448
rect 392912 426436 392918 426488
rect 172330 426368 172336 426420
rect 172388 426408 172394 426420
rect 172882 426408 172888 426420
rect 172388 426380 172888 426408
rect 172388 426368 172394 426380
rect 172882 426368 172888 426380
rect 172940 426408 172946 426420
rect 445754 426408 445760 426420
rect 172940 426380 445760 426408
rect 172940 426368 172946 426380
rect 445754 426368 445760 426380
rect 445812 426368 445818 426420
rect 173158 426300 173164 426352
rect 173216 426340 173222 426352
rect 190454 426340 190460 426352
rect 173216 426312 190460 426340
rect 173216 426300 173222 426312
rect 190454 426300 190460 426312
rect 190512 426340 190518 426352
rect 191742 426340 191748 426352
rect 190512 426312 191748 426340
rect 190512 426300 190518 426312
rect 191742 426300 191748 426312
rect 191800 426300 191806 426352
rect 328730 425892 328736 425944
rect 328788 425932 328794 425944
rect 396810 425932 396816 425944
rect 328788 425904 396816 425932
rect 328788 425892 328794 425904
rect 396810 425892 396816 425904
rect 396868 425892 396874 425944
rect 321186 425824 321192 425876
rect 321244 425864 321250 425876
rect 400858 425864 400864 425876
rect 321244 425836 400864 425864
rect 321244 425824 321250 425836
rect 400858 425824 400864 425836
rect 400916 425824 400922 425876
rect 318702 425756 318708 425808
rect 318760 425796 318766 425808
rect 406378 425796 406384 425808
rect 318760 425768 406384 425796
rect 318760 425756 318766 425768
rect 406378 425756 406384 425768
rect 406436 425756 406442 425808
rect 504358 425756 504364 425808
rect 504416 425796 504422 425808
rect 550082 425796 550088 425808
rect 504416 425768 550088 425796
rect 504416 425756 504422 425768
rect 550082 425756 550088 425768
rect 550140 425756 550146 425808
rect 313642 425688 313648 425740
rect 313700 425728 313706 425740
rect 405090 425728 405096 425740
rect 313700 425700 405096 425728
rect 313700 425688 313706 425700
rect 405090 425688 405096 425700
rect 405148 425688 405154 425740
rect 480898 425688 480904 425740
rect 480956 425728 480962 425740
rect 536190 425728 536196 425740
rect 480956 425700 536196 425728
rect 480956 425688 480962 425700
rect 536190 425688 536196 425700
rect 536248 425688 536254 425740
rect 332502 425008 332508 425060
rect 332560 425048 332566 425060
rect 342714 425048 342720 425060
rect 332560 425020 342720 425048
rect 332560 425008 332566 425020
rect 342714 425008 342720 425020
rect 342772 425008 342778 425060
rect 288526 424940 288532 424992
rect 288584 424980 288590 424992
rect 341702 424980 341708 424992
rect 288584 424952 341708 424980
rect 288584 424940 288590 424952
rect 341702 424940 341708 424952
rect 341760 424940 341766 424992
rect 287238 424872 287244 424924
rect 287296 424912 287302 424924
rect 342898 424912 342904 424924
rect 287296 424884 342904 424912
rect 287296 424872 287302 424884
rect 342898 424872 342904 424884
rect 342956 424872 342962 424924
rect 286042 424804 286048 424856
rect 286100 424844 286106 424856
rect 342806 424844 342812 424856
rect 286100 424816 342812 424844
rect 286100 424804 286106 424816
rect 342806 424804 342812 424816
rect 342864 424804 342870 424856
rect 300762 424736 300768 424788
rect 300820 424776 300826 424788
rect 480622 424776 480628 424788
rect 300820 424748 480628 424776
rect 300820 424736 300826 424748
rect 480622 424736 480628 424748
rect 480680 424736 480686 424788
rect 299382 424668 299388 424720
rect 299440 424708 299446 424720
rect 481910 424708 481916 424720
rect 299440 424680 481916 424708
rect 299440 424668 299446 424680
rect 481910 424668 481916 424680
rect 481968 424668 481974 424720
rect 296622 424600 296628 424652
rect 296680 424640 296686 424652
rect 483198 424640 483204 424652
rect 296680 424612 483204 424640
rect 296680 424600 296686 424612
rect 483198 424600 483204 424612
rect 483256 424600 483262 424652
rect 241422 424532 241428 424584
rect 241480 424572 241486 424584
rect 510798 424572 510804 424584
rect 241480 424544 510804 424572
rect 241480 424532 241486 424544
rect 510798 424532 510804 424544
rect 510856 424532 510862 424584
rect 238662 424464 238668 424516
rect 238720 424504 238726 424516
rect 512178 424504 512184 424516
rect 238720 424476 512184 424504
rect 238720 424464 238726 424476
rect 512178 424464 512184 424476
rect 512236 424464 512242 424516
rect 235902 424396 235908 424448
rect 235960 424436 235966 424448
rect 513374 424436 513380 424448
rect 235960 424408 513380 424436
rect 235960 424396 235966 424408
rect 513374 424396 513380 424408
rect 513432 424396 513438 424448
rect 231762 424328 231768 424380
rect 231820 424368 231826 424380
rect 516134 424368 516140 424380
rect 231820 424340 516140 424368
rect 231820 424328 231826 424340
rect 516134 424328 516140 424340
rect 516192 424328 516198 424380
rect 170122 423580 170128 423632
rect 170180 423620 170186 423632
rect 440234 423620 440240 423632
rect 170180 423592 440240 423620
rect 170180 423580 170186 423592
rect 440234 423580 440240 423592
rect 440292 423580 440298 423632
rect 171410 423512 171416 423564
rect 171468 423552 171474 423564
rect 437566 423552 437572 423564
rect 171468 423524 437572 423552
rect 171468 423512 171474 423524
rect 437566 423512 437572 423524
rect 437624 423512 437630 423564
rect 245746 423036 245752 423088
rect 245804 423076 245810 423088
rect 338114 423076 338120 423088
rect 245804 423048 338120 423076
rect 245804 423036 245810 423048
rect 338114 423036 338120 423048
rect 338172 423036 338178 423088
rect 487798 423036 487804 423088
rect 487856 423076 487862 423088
rect 539686 423076 539692 423088
rect 487856 423048 539692 423076
rect 487856 423036 487862 423048
rect 539686 423036 539692 423048
rect 539744 423036 539750 423088
rect 271782 422968 271788 423020
rect 271840 423008 271846 423020
rect 495710 423008 495716 423020
rect 271840 422980 495716 423008
rect 271840 422968 271846 422980
rect 495710 422968 495716 422980
rect 495768 422968 495774 423020
rect 199378 422900 199384 422952
rect 199436 422940 199442 422952
rect 213362 422940 213368 422952
rect 199436 422912 213368 422940
rect 199436 422900 199442 422912
rect 213362 422900 213368 422912
rect 213420 422900 213426 422952
rect 269022 422900 269028 422952
rect 269080 422940 269086 422952
rect 496998 422940 497004 422952
rect 269080 422912 497004 422940
rect 269080 422900 269086 422912
rect 496998 422900 497004 422912
rect 497056 422900 497062 422952
rect 168098 422288 168104 422340
rect 168156 422328 168162 422340
rect 171410 422328 171416 422340
rect 168156 422300 171416 422328
rect 168156 422288 168162 422300
rect 171410 422288 171416 422300
rect 171468 422288 171474 422340
rect 410518 422152 410524 422204
rect 410576 422192 410582 422204
rect 425238 422192 425244 422204
rect 410576 422164 425244 422192
rect 410576 422152 410582 422164
rect 425238 422152 425244 422164
rect 425296 422152 425302 422204
rect 407850 422084 407856 422136
rect 407908 422124 407914 422136
rect 435358 422124 435364 422136
rect 407908 422096 435364 422124
rect 407908 422084 407914 422096
rect 435358 422084 435364 422096
rect 435416 422084 435422 422136
rect 408126 422016 408132 422068
rect 408184 422056 408190 422068
rect 436646 422056 436652 422068
rect 408184 422028 436652 422056
rect 408184 422016 408190 422028
rect 436646 422016 436652 422028
rect 436704 422016 436710 422068
rect 407942 421948 407948 422000
rect 408000 421988 408006 422000
rect 440326 421988 440332 422000
rect 408000 421960 440332 421988
rect 408000 421948 408006 421960
rect 440326 421948 440332 421960
rect 440384 421948 440390 422000
rect 530578 421948 530584 422000
rect 530636 421988 530642 422000
rect 545942 421988 545948 422000
rect 530636 421960 545948 421988
rect 530636 421948 530642 421960
rect 545942 421948 545948 421960
rect 546000 421948 546006 422000
rect 408034 421880 408040 421932
rect 408092 421920 408098 421932
rect 441706 421920 441712 421932
rect 408092 421892 441712 421920
rect 408092 421880 408098 421892
rect 441706 421880 441712 421892
rect 441764 421880 441770 421932
rect 471238 421880 471244 421932
rect 471296 421920 471302 421932
rect 488166 421920 488172 421932
rect 471296 421892 488172 421920
rect 471296 421880 471302 421892
rect 488166 421880 488172 421892
rect 488224 421880 488230 421932
rect 514662 421880 514668 421932
rect 514720 421920 514726 421932
rect 554774 421920 554780 421932
rect 514720 421892 554780 421920
rect 514720 421880 514726 421892
rect 554774 421880 554780 421892
rect 554832 421880 554838 421932
rect 284754 421812 284760 421864
rect 284812 421852 284818 421864
rect 342254 421852 342260 421864
rect 284812 421824 342260 421852
rect 284812 421812 284818 421824
rect 342254 421812 342260 421824
rect 342312 421812 342318 421864
rect 407758 421812 407764 421864
rect 407816 421852 407822 421864
rect 446582 421852 446588 421864
rect 407816 421824 446588 421852
rect 407816 421812 407822 421824
rect 446582 421812 446588 421824
rect 446640 421812 446646 421864
rect 447778 421812 447784 421864
rect 447836 421852 447842 421864
rect 485774 421852 485780 421864
rect 447836 421824 485780 421852
rect 447836 421812 447842 421824
rect 485774 421812 485780 421824
rect 485832 421812 485838 421864
rect 509142 421812 509148 421864
rect 509200 421852 509206 421864
rect 552198 421852 552204 421864
rect 509200 421824 552204 421852
rect 509200 421812 509206 421824
rect 552198 421812 552204 421824
rect 552256 421812 552262 421864
rect 341518 421744 341524 421796
rect 341576 421784 341582 421796
rect 427814 421784 427820 421796
rect 341576 421756 427820 421784
rect 341576 421744 341582 421756
rect 427814 421744 427820 421756
rect 427872 421744 427878 421796
rect 436738 421744 436744 421796
rect 436796 421784 436802 421796
rect 484394 421784 484400 421796
rect 436796 421756 484400 421784
rect 436796 421744 436802 421756
rect 484394 421744 484400 421756
rect 484452 421744 484458 421796
rect 499482 421744 499488 421796
rect 499540 421784 499546 421796
rect 547230 421784 547236 421796
rect 499540 421756 547236 421784
rect 499540 421744 499546 421756
rect 547230 421744 547236 421756
rect 547288 421744 547294 421796
rect 196618 421676 196624 421728
rect 196676 421716 196682 421728
rect 397638 421716 397644 421728
rect 196676 421688 397644 421716
rect 196676 421676 196682 421688
rect 397638 421676 397644 421688
rect 397696 421676 397702 421728
rect 409782 421676 409788 421728
rect 409840 421716 409846 421728
rect 470686 421716 470692 421728
rect 409840 421688 470692 421716
rect 409840 421676 409846 421688
rect 470686 421676 470692 421688
rect 470744 421676 470750 421728
rect 474642 421676 474648 421728
rect 474700 421716 474706 421728
rect 546678 421716 546684 421728
rect 474700 421688 546684 421716
rect 474700 421676 474706 421688
rect 546678 421676 546684 421688
rect 546736 421676 546742 421728
rect 193858 421608 193864 421660
rect 193916 421648 193922 421660
rect 400214 421648 400220 421660
rect 193916 421620 400220 421648
rect 193916 421608 193922 421620
rect 400214 421608 400220 421620
rect 400272 421608 400278 421660
rect 408310 421608 408316 421660
rect 408368 421648 408374 421660
rect 471974 421648 471980 421660
rect 408368 421620 471980 421648
rect 408368 421608 408374 421620
rect 471974 421608 471980 421620
rect 472032 421608 472038 421660
rect 475838 421608 475844 421660
rect 475896 421648 475902 421660
rect 547874 421648 547880 421660
rect 475896 421620 547880 421648
rect 475896 421608 475902 421620
rect 547874 421608 547880 421620
rect 547932 421608 547938 421660
rect 199562 421540 199568 421592
rect 199620 421580 199626 421592
rect 407574 421580 407580 421592
rect 199620 421552 407580 421580
rect 199620 421540 199626 421552
rect 407574 421540 407580 421552
rect 407632 421540 407638 421592
rect 408402 421540 408408 421592
rect 408460 421580 408466 421592
rect 465534 421580 465540 421592
rect 408460 421552 465540 421580
rect 408460 421540 408466 421552
rect 465534 421540 465540 421552
rect 465592 421540 465598 421592
rect 469582 421540 469588 421592
rect 469640 421580 469646 421592
rect 546770 421580 546776 421592
rect 469640 421552 546776 421580
rect 469640 421540 469646 421552
rect 546770 421540 546776 421552
rect 546828 421540 546834 421592
rect 195238 421472 195244 421524
rect 195296 421512 195302 421524
rect 403894 421512 403900 421524
rect 195296 421484 403900 421512
rect 195296 421472 195302 421484
rect 403894 421472 403900 421484
rect 403952 421472 403958 421524
rect 196986 421404 196992 421456
rect 197044 421444 197050 421456
rect 408862 421444 408868 421456
rect 197044 421416 408868 421444
rect 197044 421404 197050 421416
rect 408862 421404 408868 421416
rect 408920 421404 408926 421456
rect 197078 421336 197084 421388
rect 197136 421376 197142 421388
rect 415394 421376 415400 421388
rect 197136 421348 415400 421376
rect 197136 421336 197142 421348
rect 415394 421336 415400 421348
rect 415452 421336 415458 421388
rect 197170 421268 197176 421320
rect 197228 421308 197234 421320
rect 416774 421308 416780 421320
rect 197228 421280 416780 421308
rect 197228 421268 197234 421280
rect 416774 421268 416780 421280
rect 416832 421268 416838 421320
rect 173158 421200 173164 421252
rect 173216 421240 173222 421252
rect 393774 421240 393780 421252
rect 173216 421212 393780 421240
rect 173216 421200 173222 421212
rect 393774 421200 393780 421212
rect 393832 421200 393838 421252
rect 173250 421132 173256 421184
rect 173308 421172 173314 421184
rect 398926 421172 398932 421184
rect 173308 421144 398932 421172
rect 173308 421132 173314 421144
rect 398926 421132 398932 421144
rect 398984 421132 398990 421184
rect 172146 421064 172152 421116
rect 172204 421104 172210 421116
rect 406470 421104 406476 421116
rect 172204 421076 406476 421104
rect 172204 421064 172210 421076
rect 406470 421064 406476 421076
rect 406528 421064 406534 421116
rect 172238 420996 172244 421048
rect 172296 421036 172302 421048
rect 412818 421036 412824 421048
rect 172296 421008 412824 421036
rect 172296 420996 172302 421008
rect 412818 420996 412824 421008
rect 412876 420996 412882 421048
rect 413278 420996 413284 421048
rect 413336 421036 413342 421048
rect 420270 421036 420276 421048
rect 413336 421008 420276 421036
rect 413336 420996 413342 421008
rect 420270 420996 420276 421008
rect 420328 420996 420334 421048
rect 173526 420928 173532 420980
rect 173584 420968 173590 420980
rect 414014 420968 414020 420980
rect 173584 420940 414020 420968
rect 173584 420928 173590 420940
rect 414014 420928 414020 420940
rect 414072 420928 414078 420980
rect 485038 420928 485044 420980
rect 485096 420968 485102 420980
rect 487154 420968 487160 420980
rect 485096 420940 487160 420968
rect 485096 420928 485102 420940
rect 487154 420928 487160 420940
rect 487212 420928 487218 420980
rect 199470 420180 199476 420232
rect 199528 420220 199534 420232
rect 213178 420220 213184 420232
rect 199528 420192 213184 420220
rect 199528 420180 199534 420192
rect 213178 420180 213184 420192
rect 213236 420180 213242 420232
rect 181438 419704 181444 419756
rect 181496 419744 181502 419756
rect 402974 419744 402980 419756
rect 181496 419716 402980 419744
rect 181496 419704 181502 419716
rect 402974 419704 402980 419716
rect 403032 419704 403038 419756
rect 195514 419636 195520 419688
rect 195572 419676 195578 419688
rect 418982 419676 418988 419688
rect 195572 419648 418988 419676
rect 195572 419636 195578 419648
rect 418982 419636 418988 419648
rect 419040 419636 419046 419688
rect 184382 419568 184388 419620
rect 184440 419608 184446 419620
rect 410150 419608 410156 419620
rect 184440 419580 410156 419608
rect 184440 419568 184446 419580
rect 410150 419568 410156 419580
rect 410208 419568 410214 419620
rect 187510 419500 187516 419552
rect 187568 419540 187574 419552
rect 417694 419540 417700 419552
rect 187568 419512 417700 419540
rect 187568 419500 187574 419512
rect 417694 419500 417700 419512
rect 417752 419500 417758 419552
rect 179046 419432 179052 419484
rect 179104 419472 179110 419484
rect 197354 419472 197360 419484
rect 179104 419444 197360 419472
rect 179104 419432 179110 419444
rect 197354 419432 197360 419444
rect 197412 419432 197418 419484
rect 189810 416712 189816 416764
rect 189868 416752 189874 416764
rect 197354 416752 197360 416764
rect 189868 416724 197360 416752
rect 189868 416712 189874 416724
rect 197354 416712 197360 416724
rect 197412 416712 197418 416764
rect 177574 415352 177580 415404
rect 177632 415392 177638 415404
rect 197354 415392 197360 415404
rect 177632 415364 197360 415392
rect 177632 415352 177638 415364
rect 197354 415352 197360 415364
rect 197412 415352 197418 415404
rect 560202 415352 560208 415404
rect 560260 415392 560266 415404
rect 580258 415392 580264 415404
rect 560260 415364 580264 415392
rect 560260 415352 560266 415364
rect 580258 415352 580264 415364
rect 580316 415352 580322 415404
rect 182910 413924 182916 413976
rect 182968 413964 182974 413976
rect 197354 413964 197360 413976
rect 182968 413936 197360 413964
rect 182968 413924 182974 413936
rect 197354 413924 197360 413936
rect 197412 413924 197418 413976
rect 184474 412564 184480 412616
rect 184532 412604 184538 412616
rect 197354 412604 197360 412616
rect 184532 412576 197360 412604
rect 184532 412564 184538 412576
rect 197354 412564 197360 412576
rect 197412 412564 197418 412616
rect 3418 411204 3424 411256
rect 3476 411244 3482 411256
rect 28442 411244 28448 411256
rect 3476 411216 28448 411244
rect 3476 411204 3482 411216
rect 28442 411204 28448 411216
rect 28500 411204 28506 411256
rect 188522 411204 188528 411256
rect 188580 411244 188586 411256
rect 197354 411244 197360 411256
rect 188580 411216 197360 411244
rect 188580 411204 188586 411216
rect 197354 411204 197360 411216
rect 197412 411204 197418 411256
rect 170950 409776 170956 409828
rect 171008 409816 171014 409828
rect 197354 409816 197360 409828
rect 171008 409788 197360 409816
rect 171008 409776 171014 409788
rect 197354 409776 197360 409788
rect 197412 409776 197418 409828
rect 191282 409708 191288 409760
rect 191340 409748 191346 409760
rect 197446 409748 197452 409760
rect 191340 409720 197452 409748
rect 191340 409708 191346 409720
rect 197446 409708 197452 409720
rect 197504 409708 197510 409760
rect 170214 408416 170220 408468
rect 170272 408456 170278 408468
rect 171318 408456 171324 408468
rect 170272 408428 171324 408456
rect 170272 408416 170278 408428
rect 171318 408416 171324 408428
rect 171376 408416 171382 408468
rect 194042 408416 194048 408468
rect 194100 408456 194106 408468
rect 197354 408456 197360 408468
rect 194100 408428 197360 408456
rect 194100 408416 194106 408428
rect 197354 408416 197360 408428
rect 197412 408416 197418 408468
rect 560110 408416 560116 408468
rect 560168 408456 560174 408468
rect 577498 408456 577504 408468
rect 560168 408428 577504 408456
rect 560168 408416 560174 408428
rect 577498 408416 577504 408428
rect 577556 408416 577562 408468
rect 195422 407056 195428 407108
rect 195480 407096 195486 407108
rect 197722 407096 197728 407108
rect 195480 407068 197728 407096
rect 195480 407056 195486 407068
rect 197722 407056 197728 407068
rect 197780 407056 197786 407108
rect 181622 405628 181628 405680
rect 181680 405668 181686 405680
rect 197354 405668 197360 405680
rect 181680 405640 197360 405668
rect 181680 405628 181686 405640
rect 197354 405628 197360 405640
rect 197412 405628 197418 405680
rect 574830 404336 574836 404388
rect 574888 404376 574894 404388
rect 580166 404376 580172 404388
rect 574888 404348 580172 404376
rect 574888 404336 574894 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 192478 404268 192484 404320
rect 192536 404308 192542 404320
rect 197354 404308 197360 404320
rect 192536 404280 197360 404308
rect 192536 404268 192542 404280
rect 197354 404268 197360 404280
rect 197412 404268 197418 404320
rect 185670 401548 185676 401600
rect 185728 401588 185734 401600
rect 197354 401588 197360 401600
rect 185728 401560 197360 401588
rect 185728 401548 185734 401560
rect 197354 401548 197360 401560
rect 197412 401548 197418 401600
rect 170858 400120 170864 400172
rect 170916 400160 170922 400172
rect 197354 400160 197360 400172
rect 170916 400132 197360 400160
rect 170916 400120 170922 400132
rect 197354 400120 197360 400132
rect 197412 400120 197418 400172
rect 560018 400120 560024 400172
rect 560076 400160 560082 400172
rect 570598 400160 570604 400172
rect 560076 400132 570604 400160
rect 560076 400120 560082 400132
rect 570598 400120 570604 400132
rect 570656 400120 570662 400172
rect 3234 398760 3240 398812
rect 3292 398800 3298 398812
rect 28350 398800 28356 398812
rect 3292 398772 28356 398800
rect 3292 398760 3298 398772
rect 28350 398760 28356 398772
rect 28408 398760 28414 398812
rect 170766 398760 170772 398812
rect 170824 398800 170830 398812
rect 197354 398800 197360 398812
rect 170824 398772 197360 398800
rect 170824 398760 170830 398772
rect 197354 398760 197360 398772
rect 197412 398760 197418 398812
rect 174630 398692 174636 398744
rect 174688 398732 174694 398744
rect 197446 398732 197452 398744
rect 174688 398704 197452 398732
rect 174688 398692 174694 398704
rect 197446 398692 197452 398704
rect 197504 398692 197510 398744
rect 168834 398284 168840 398336
rect 168892 398324 168898 398336
rect 169938 398324 169944 398336
rect 168892 398296 169944 398324
rect 168892 398284 168898 398296
rect 169938 398284 169944 398296
rect 169996 398284 170002 398336
rect 174722 397400 174728 397452
rect 174780 397440 174786 397452
rect 197354 397440 197360 397452
rect 174780 397412 197360 397440
rect 174780 397400 174786 397412
rect 197354 397400 197360 397412
rect 197412 397400 197418 397452
rect 176194 395972 176200 396024
rect 176252 396012 176258 396024
rect 197354 396012 197360 396024
rect 176252 395984 197360 396012
rect 176252 395972 176258 395984
rect 197354 395972 197360 395984
rect 197412 395972 197418 396024
rect 187142 394612 187148 394664
rect 187200 394652 187206 394664
rect 197354 394652 197360 394664
rect 187200 394624 197360 394652
rect 187200 394612 187206 394624
rect 197354 394612 197360 394624
rect 197412 394612 197418 394664
rect 169478 393252 169484 393304
rect 169536 393292 169542 393304
rect 174170 393292 174176 393304
rect 169536 393264 174176 393292
rect 169536 393252 169542 393264
rect 174170 393252 174176 393264
rect 174228 393252 174234 393304
rect 177482 393252 177488 393304
rect 177540 393292 177546 393304
rect 197354 393292 197360 393304
rect 177540 393264 197360 393292
rect 177540 393252 177546 393264
rect 197354 393252 197360 393264
rect 197412 393252 197418 393304
rect 169110 391960 169116 392012
rect 169168 392000 169174 392012
rect 169478 392000 169484 392012
rect 169168 391972 169484 392000
rect 169168 391960 169174 391972
rect 169478 391960 169484 391972
rect 169536 391960 169542 392012
rect 184290 391892 184296 391944
rect 184348 391932 184354 391944
rect 197354 391932 197360 391944
rect 184348 391904 197360 391932
rect 184348 391892 184354 391904
rect 197354 391892 197360 391904
rect 197412 391892 197418 391944
rect 560202 391892 560208 391944
rect 560260 391932 560266 391944
rect 578878 391932 578884 391944
rect 560260 391904 578884 391932
rect 560260 391892 560266 391904
rect 578878 391892 578884 391904
rect 578936 391892 578942 391944
rect 188430 390464 188436 390516
rect 188488 390504 188494 390516
rect 197354 390504 197360 390516
rect 188488 390476 197360 390504
rect 188488 390464 188494 390476
rect 197354 390464 197360 390476
rect 197412 390464 197418 390516
rect 191190 389104 191196 389156
rect 191248 389144 191254 389156
rect 197354 389144 197360 389156
rect 191248 389116 197360 389144
rect 191248 389104 191254 389116
rect 197354 389104 197360 389116
rect 197412 389104 197418 389156
rect 180058 387744 180064 387796
rect 180116 387784 180122 387796
rect 197354 387784 197360 387796
rect 180116 387756 197360 387784
rect 180116 387744 180122 387756
rect 197354 387744 197360 387756
rect 197412 387744 197418 387796
rect 195330 386316 195336 386368
rect 195388 386356 195394 386368
rect 197722 386356 197728 386368
rect 195388 386328 197728 386356
rect 195388 386316 195394 386328
rect 197722 386316 197728 386328
rect 197780 386316 197786 386368
rect 193950 386248 193956 386300
rect 194008 386288 194014 386300
rect 197354 386288 197360 386300
rect 194008 386260 197360 386288
rect 194008 386248 194014 386260
rect 197354 386248 197360 386260
rect 197412 386248 197418 386300
rect 167730 384956 167736 385008
rect 167788 384996 167794 385008
rect 197354 384996 197360 385008
rect 167788 384968 197360 384996
rect 167788 384956 167794 384968
rect 197354 384956 197360 384968
rect 197412 384956 197418 385008
rect 178954 383596 178960 383648
rect 179012 383636 179018 383648
rect 197354 383636 197360 383648
rect 179012 383608 197360 383636
rect 179012 383596 179018 383608
rect 197354 383596 197360 383608
rect 197412 383596 197418 383648
rect 559190 383392 559196 383444
rect 559248 383432 559254 383444
rect 560938 383432 560944 383444
rect 559248 383404 560944 383432
rect 559248 383392 559254 383404
rect 560938 383392 560944 383404
rect 560996 383392 561002 383444
rect 167638 382168 167644 382220
rect 167696 382208 167702 382220
rect 197354 382208 197360 382220
rect 167696 382180 197360 382208
rect 167696 382168 167702 382180
rect 197354 382168 197360 382180
rect 197412 382168 197418 382220
rect 181530 380808 181536 380860
rect 181588 380848 181594 380860
rect 197354 380848 197360 380860
rect 181588 380820 197360 380848
rect 181588 380808 181594 380820
rect 197354 380808 197360 380820
rect 197412 380808 197418 380860
rect 167546 379448 167552 379500
rect 167604 379488 167610 379500
rect 197354 379488 197360 379500
rect 167604 379460 197360 379488
rect 167604 379448 167610 379460
rect 197354 379448 197360 379460
rect 197412 379448 197418 379500
rect 570598 378156 570604 378208
rect 570656 378196 570662 378208
rect 580166 378196 580172 378208
rect 570656 378168 580172 378196
rect 570656 378156 570662 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 188706 378088 188712 378140
rect 188764 378128 188770 378140
rect 197354 378128 197360 378140
rect 188764 378100 197360 378128
rect 188764 378088 188770 378100
rect 197354 378088 197360 378100
rect 197412 378088 197418 378140
rect 174998 376660 175004 376712
rect 175056 376700 175062 376712
rect 197354 376700 197360 376712
rect 175056 376672 197360 376700
rect 175056 376660 175062 376672
rect 197354 376660 197360 376672
rect 197412 376660 197418 376712
rect 187418 375300 187424 375352
rect 187476 375340 187482 375352
rect 197354 375340 197360 375352
rect 187476 375312 197360 375340
rect 187476 375300 187482 375312
rect 197354 375300 197360 375312
rect 197412 375300 197418 375352
rect 560202 375300 560208 375352
rect 560260 375340 560266 375352
rect 567838 375340 567844 375352
rect 560260 375312 567844 375340
rect 560260 375300 560266 375312
rect 567838 375300 567844 375312
rect 567896 375300 567902 375352
rect 184750 373940 184756 373992
rect 184808 373980 184814 373992
rect 197354 373980 197360 373992
rect 184808 373952 197360 373980
rect 184808 373940 184814 373952
rect 197354 373940 197360 373952
rect 197412 373940 197418 373992
rect 177758 372512 177764 372564
rect 177816 372552 177822 372564
rect 197354 372552 197360 372564
rect 177816 372524 197360 372552
rect 177816 372512 177822 372524
rect 197354 372512 197360 372524
rect 197412 372512 197418 372564
rect 193766 372444 193772 372496
rect 193824 372484 193830 372496
rect 197446 372484 197452 372496
rect 193824 372456 197452 372484
rect 193824 372444 193830 372456
rect 197446 372444 197452 372456
rect 197504 372444 197510 372496
rect 195146 371152 195152 371204
rect 195204 371192 195210 371204
rect 197354 371192 197360 371204
rect 195204 371164 197360 371192
rect 195204 371152 195210 371164
rect 197354 371152 197360 371164
rect 197412 371152 197418 371204
rect 189994 369792 190000 369844
rect 190052 369832 190058 369844
rect 197354 369832 197360 369844
rect 190052 369804 197360 369832
rect 190052 369792 190058 369804
rect 197354 369792 197360 369804
rect 197412 369792 197418 369844
rect 185854 368432 185860 368484
rect 185912 368472 185918 368484
rect 197354 368472 197360 368484
rect 185912 368444 197360 368472
rect 185912 368432 185918 368444
rect 197354 368432 197360 368444
rect 197412 368432 197418 368484
rect 559190 367412 559196 367464
rect 559248 367452 559254 367464
rect 565078 367452 565084 367464
rect 559248 367424 565084 367452
rect 559248 367412 559254 367424
rect 565078 367412 565084 367424
rect 565136 367412 565142 367464
rect 183094 367004 183100 367056
rect 183152 367044 183158 367056
rect 197354 367044 197360 367056
rect 183152 367016 197360 367044
rect 183152 367004 183158 367016
rect 197354 367004 197360 367016
rect 197412 367004 197418 367056
rect 3418 365644 3424 365696
rect 3476 365684 3482 365696
rect 197170 365684 197176 365696
rect 3476 365656 197176 365684
rect 3476 365644 3482 365656
rect 197170 365644 197176 365656
rect 197228 365644 197234 365696
rect 174906 365576 174912 365628
rect 174964 365616 174970 365628
rect 197354 365616 197360 365628
rect 174964 365588 197360 365616
rect 174964 365576 174970 365588
rect 197354 365576 197360 365588
rect 197412 365576 197418 365628
rect 3418 365100 3424 365152
rect 3476 365140 3482 365152
rect 197814 365140 197820 365152
rect 3476 365112 197820 365140
rect 3476 365100 3482 365112
rect 197814 365100 197820 365112
rect 197872 365100 197878 365152
rect 3602 365032 3608 365084
rect 3660 365072 3666 365084
rect 199562 365072 199568 365084
rect 3660 365044 199568 365072
rect 3660 365032 3666 365044
rect 199562 365032 199568 365044
rect 199620 365032 199626 365084
rect 3510 364964 3516 365016
rect 3568 365004 3574 365016
rect 200114 365004 200120 365016
rect 3568 364976 200120 365004
rect 3568 364964 3574 364976
rect 200114 364964 200120 364976
rect 200172 364964 200178 365016
rect 559558 364352 559564 364404
rect 559616 364392 559622 364404
rect 579614 364392 579620 364404
rect 559616 364364 579620 364392
rect 559616 364352 559622 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 139210 364284 139216 364336
rect 139268 364324 139274 364336
rect 168098 364324 168104 364336
rect 139268 364296 168104 364324
rect 139268 364284 139274 364296
rect 168098 364284 168104 364296
rect 168156 364284 168162 364336
rect 176378 364284 176384 364336
rect 176436 364324 176442 364336
rect 197354 364324 197360 364336
rect 176436 364296 197360 364324
rect 176436 364284 176442 364296
rect 197354 364284 197360 364296
rect 197412 364284 197418 364336
rect 167178 364148 167184 364200
rect 167236 364188 167242 364200
rect 178770 364188 178776 364200
rect 167236 364160 178776 364188
rect 167236 364148 167242 364160
rect 178770 364148 178776 364160
rect 178828 364148 178834 364200
rect 136542 364080 136548 364132
rect 136600 364120 136606 364132
rect 168190 364120 168196 364132
rect 136600 364092 168196 364120
rect 136600 364080 136606 364092
rect 168190 364080 168196 364092
rect 168248 364080 168254 364132
rect 130930 363944 130936 363996
rect 130988 363984 130994 363996
rect 172330 363984 172336 363996
rect 130988 363956 172336 363984
rect 130988 363944 130994 363956
rect 172330 363944 172336 363956
rect 172388 363944 172394 363996
rect 125502 363876 125508 363928
rect 125560 363916 125566 363928
rect 173618 363916 173624 363928
rect 125560 363888 173624 363916
rect 125560 363876 125566 363888
rect 173618 363876 173624 363888
rect 173676 363876 173682 363928
rect 29638 363808 29644 363860
rect 29696 363848 29702 363860
rect 42794 363848 42800 363860
rect 29696 363820 42800 363848
rect 29696 363808 29702 363820
rect 42794 363808 42800 363820
rect 42852 363808 42858 363860
rect 129642 363808 129648 363860
rect 129700 363848 129706 363860
rect 180334 363848 180340 363860
rect 129700 363820 180340 363848
rect 129700 363808 129706 363820
rect 180334 363808 180340 363820
rect 180392 363808 180398 363860
rect 122742 363740 122748 363792
rect 122800 363780 122806 363792
rect 177298 363780 177304 363792
rect 122800 363752 177304 363780
rect 122800 363740 122806 363752
rect 177298 363740 177304 363752
rect 177356 363740 177362 363792
rect 28626 363672 28632 363724
rect 28684 363712 28690 363724
rect 42886 363712 42892 363724
rect 28684 363684 42892 363712
rect 28684 363672 28690 363684
rect 42886 363672 42892 363684
rect 42944 363672 42950 363724
rect 29730 363604 29736 363656
rect 29788 363644 29794 363656
rect 46934 363644 46940 363656
rect 29788 363616 46940 363644
rect 29788 363604 29794 363616
rect 46934 363604 46940 363616
rect 46992 363604 46998 363656
rect 128262 363604 128268 363656
rect 128320 363644 128326 363656
rect 190454 363644 190460 363656
rect 128320 363616 190460 363644
rect 128320 363604 128326 363616
rect 190454 363604 190460 363616
rect 190512 363604 190518 363656
rect 167730 363536 167736 363588
rect 167788 363576 167794 363588
rect 170950 363576 170956 363588
rect 167788 363548 170956 363576
rect 167788 363536 167794 363548
rect 170950 363536 170956 363548
rect 171008 363576 171014 363588
rect 177850 363576 177856 363588
rect 171008 363548 177856 363576
rect 171008 363536 171014 363548
rect 177850 363536 177856 363548
rect 177908 363536 177914 363588
rect 148962 363468 148968 363520
rect 149020 363508 149026 363520
rect 170306 363508 170312 363520
rect 149020 363480 170312 363508
rect 149020 363468 149026 363480
rect 170306 363468 170312 363480
rect 170364 363468 170370 363520
rect 136542 363332 136548 363384
rect 136600 363372 136606 363384
rect 146938 363372 146944 363384
rect 136600 363344 146944 363372
rect 136600 363332 136606 363344
rect 146938 363332 146944 363344
rect 146996 363332 147002 363384
rect 137922 363264 137928 363316
rect 137980 363304 137986 363316
rect 167822 363304 167828 363316
rect 137980 363276 167828 363304
rect 137980 363264 137986 363276
rect 167822 363264 167828 363276
rect 167880 363264 167886 363316
rect 29454 362924 29460 362976
rect 29512 362964 29518 362976
rect 29638 362964 29644 362976
rect 29512 362936 29644 362964
rect 29512 362924 29518 362936
rect 29638 362924 29644 362936
rect 29696 362924 29702 362976
rect 151170 362924 151176 362976
rect 151228 362964 151234 362976
rect 167086 362964 167092 362976
rect 151228 362936 167092 362964
rect 151228 362924 151234 362936
rect 167086 362924 167092 362936
rect 167144 362964 167150 362976
rect 169846 362964 169852 362976
rect 167144 362936 169852 362964
rect 167144 362924 167150 362936
rect 169846 362924 169852 362936
rect 169904 362924 169910 362976
rect 184934 362924 184940 362976
rect 184992 362964 184998 362976
rect 187786 362964 187792 362976
rect 184992 362936 187792 362964
rect 184992 362924 184998 362936
rect 187786 362924 187792 362936
rect 187844 362924 187850 362976
rect 180150 362856 180156 362908
rect 180208 362896 180214 362908
rect 197354 362896 197360 362908
rect 180208 362868 197360 362896
rect 180208 362856 180214 362868
rect 197354 362856 197360 362868
rect 197412 362856 197418 362908
rect 138290 362380 138296 362432
rect 138348 362420 138354 362432
rect 180334 362420 180340 362432
rect 138348 362392 180340 362420
rect 138348 362380 138354 362392
rect 180334 362380 180340 362392
rect 180392 362380 180398 362432
rect 124122 362312 124128 362364
rect 124180 362352 124186 362364
rect 170766 362352 170772 362364
rect 124180 362324 170772 362352
rect 124180 362312 124186 362324
rect 170766 362312 170772 362324
rect 170824 362312 170830 362364
rect 146938 362244 146944 362296
rect 146996 362284 147002 362296
rect 168006 362284 168012 362296
rect 146996 362256 168012 362284
rect 146996 362244 147002 362256
rect 168006 362244 168012 362256
rect 168064 362284 168070 362296
rect 184290 362284 184296 362296
rect 168064 362256 184296 362284
rect 168064 362244 168070 362256
rect 184290 362244 184296 362256
rect 184348 362244 184354 362296
rect 108850 362176 108856 362228
rect 108908 362216 108914 362228
rect 177298 362216 177304 362228
rect 108908 362188 177304 362216
rect 108908 362176 108914 362188
rect 177298 362176 177304 362188
rect 177356 362176 177362 362228
rect 167914 361496 167920 361548
rect 167972 361536 167978 361548
rect 169754 361536 169760 361548
rect 167972 361508 169760 361536
rect 167972 361496 167978 361508
rect 169754 361496 169760 361508
rect 169812 361496 169818 361548
rect 179138 361496 179144 361548
rect 179196 361536 179202 361548
rect 197354 361536 197360 361548
rect 179196 361508 197360 361536
rect 179196 361496 179202 361508
rect 197354 361496 197360 361508
rect 197412 361496 197418 361548
rect 181806 361428 181812 361480
rect 181864 361468 181870 361480
rect 197446 361468 197452 361480
rect 181864 361440 197452 361468
rect 181864 361428 181870 361440
rect 197446 361428 197452 361440
rect 197504 361428 197510 361480
rect 150434 361088 150440 361140
rect 150492 361128 150498 361140
rect 167178 361128 167184 361140
rect 150492 361100 167184 361128
rect 150492 361088 150498 361100
rect 167178 361088 167184 361100
rect 167236 361128 167242 361140
rect 171042 361128 171048 361140
rect 167236 361100 171048 361128
rect 167236 361088 167242 361100
rect 171042 361088 171048 361100
rect 171100 361088 171106 361140
rect 133138 361020 133144 361072
rect 133196 361060 133202 361072
rect 167914 361060 167920 361072
rect 133196 361032 167920 361060
rect 133196 361020 133202 361032
rect 167914 361020 167920 361032
rect 167972 361020 167978 361072
rect 127618 360952 127624 361004
rect 127676 360992 127682 361004
rect 170950 360992 170956 361004
rect 127676 360964 170956 360992
rect 127676 360952 127682 360964
rect 170950 360952 170956 360964
rect 171008 360952 171014 361004
rect 143350 360884 143356 360936
rect 143408 360924 143414 360936
rect 166994 360924 167000 360936
rect 143408 360896 167000 360924
rect 143408 360884 143414 360896
rect 166994 360884 167000 360896
rect 167052 360924 167058 360936
rect 186958 360924 186964 360936
rect 167052 360896 186964 360924
rect 167052 360884 167058 360896
rect 186958 360884 186964 360896
rect 187016 360924 187022 360936
rect 193214 360924 193220 360936
rect 187016 360896 193220 360924
rect 187016 360884 187022 360896
rect 193214 360884 193220 360896
rect 193272 360884 193278 360936
rect 73154 360816 73160 360868
rect 73212 360856 73218 360868
rect 176378 360856 176384 360868
rect 73212 360828 176384 360856
rect 73212 360816 73218 360828
rect 176378 360816 176384 360828
rect 176436 360816 176442 360868
rect 140314 360136 140320 360188
rect 140372 360176 140378 360188
rect 193674 360176 193680 360188
rect 140372 360148 193680 360176
rect 140372 360136 140378 360148
rect 193674 360136 193680 360148
rect 193732 360176 193738 360188
rect 194594 360176 194600 360188
rect 193732 360148 194600 360176
rect 193732 360136 193738 360148
rect 194594 360136 194600 360148
rect 194652 360136 194658 360188
rect 560202 360136 560208 360188
rect 560260 360176 560266 360188
rect 574738 360176 574744 360188
rect 560260 360148 574744 360176
rect 560260 360136 560266 360148
rect 574738 360136 574744 360148
rect 574796 360136 574802 360188
rect 125962 360068 125968 360120
rect 126020 360108 126026 360120
rect 173802 360108 173808 360120
rect 126020 360080 173808 360108
rect 126020 360068 126026 360080
rect 173802 360068 173808 360080
rect 173860 360108 173866 360120
rect 176746 360108 176752 360120
rect 173860 360080 176752 360108
rect 173860 360068 173866 360080
rect 176746 360068 176752 360080
rect 176804 360068 176810 360120
rect 177666 360068 177672 360120
rect 177724 360108 177730 360120
rect 197354 360108 197360 360120
rect 177724 360080 197360 360108
rect 177724 360068 177730 360080
rect 197354 360068 197360 360080
rect 197412 360068 197418 360120
rect 135898 359524 135904 359576
rect 135956 359564 135962 359576
rect 174722 359564 174728 359576
rect 135956 359536 174728 359564
rect 135956 359524 135962 359536
rect 174722 359524 174728 359536
rect 174780 359524 174786 359576
rect 103146 359456 103152 359508
rect 103204 359496 103210 359508
rect 167638 359496 167644 359508
rect 103204 359468 167644 359496
rect 103204 359456 103210 359468
rect 167638 359456 167644 359468
rect 167696 359456 167702 359508
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 195514 358748 195520 358760
rect 3384 358720 195520 358748
rect 3384 358708 3390 358720
rect 195514 358708 195520 358720
rect 195572 358708 195578 358760
rect 114370 358640 114376 358692
rect 114428 358680 114434 358692
rect 172606 358680 172612 358692
rect 114428 358652 172612 358680
rect 114428 358640 114434 358652
rect 172606 358640 172612 358652
rect 172664 358680 172670 358692
rect 173802 358680 173808 358692
rect 172664 358652 173808 358680
rect 172664 358640 172670 358652
rect 173802 358640 173808 358652
rect 173860 358640 173866 358692
rect 188614 358640 188620 358692
rect 188672 358680 188678 358692
rect 197354 358680 197360 358692
rect 188672 358652 197360 358680
rect 188672 358640 188678 358652
rect 197354 358640 197360 358652
rect 197412 358640 197418 358692
rect 132034 358096 132040 358148
rect 132092 358136 132098 358148
rect 184934 358136 184940 358148
rect 132092 358108 184940 358136
rect 132092 358096 132098 358108
rect 184934 358096 184940 358108
rect 184992 358096 184998 358148
rect 63402 358028 63408 358080
rect 63460 358068 63466 358080
rect 166258 358068 166264 358080
rect 63460 358040 166264 358068
rect 63460 358028 63466 358040
rect 166258 358028 166264 358040
rect 166316 358028 166322 358080
rect 173802 358028 173808 358080
rect 173860 358068 173866 358080
rect 187878 358068 187884 358080
rect 173860 358040 187884 358068
rect 173860 358028 173866 358040
rect 187878 358028 187884 358040
rect 187936 358028 187942 358080
rect 184658 357348 184664 357400
rect 184716 357388 184722 357400
rect 197354 357388 197360 357400
rect 184716 357360 197360 357388
rect 184716 357348 184722 357360
rect 197354 357348 197360 357360
rect 197412 357348 197418 357400
rect 132954 356872 132960 356924
rect 133012 356912 133018 356924
rect 181806 356912 181812 356924
rect 133012 356884 181812 356912
rect 133012 356872 133018 356884
rect 181806 356872 181812 356884
rect 181864 356872 181870 356924
rect 136450 356804 136456 356856
rect 136508 356844 136514 356856
rect 191834 356844 191840 356856
rect 136508 356816 191840 356844
rect 136508 356804 136514 356816
rect 191834 356804 191840 356816
rect 191892 356804 191898 356856
rect 119982 356736 119988 356788
rect 120040 356776 120046 356788
rect 189166 356776 189172 356788
rect 120040 356748 189172 356776
rect 120040 356736 120046 356748
rect 189166 356736 189172 356748
rect 189224 356736 189230 356788
rect 95602 356668 95608 356720
rect 95660 356708 95666 356720
rect 167822 356708 167828 356720
rect 95660 356680 167828 356708
rect 95660 356668 95666 356680
rect 167822 356668 167828 356680
rect 167880 356668 167886 356720
rect 109586 355988 109592 356040
rect 109644 356028 109650 356040
rect 169846 356028 169852 356040
rect 109644 356000 169852 356028
rect 109644 355988 109650 356000
rect 169846 355988 169852 356000
rect 169904 356028 169910 356040
rect 170214 356028 170220 356040
rect 169904 356000 170220 356028
rect 169904 355988 169910 356000
rect 170214 355988 170220 356000
rect 170272 355988 170278 356040
rect 187234 355988 187240 356040
rect 187292 356028 187298 356040
rect 197354 356028 197360 356040
rect 187292 356000 197360 356028
rect 187292 355988 187298 356000
rect 197354 355988 197360 356000
rect 197412 355988 197418 356040
rect 169846 355512 169852 355564
rect 169904 355552 169910 355564
rect 174630 355552 174636 355564
rect 169904 355524 174636 355552
rect 169904 355512 169910 355524
rect 174630 355512 174636 355524
rect 174688 355512 174694 355564
rect 128262 355444 128268 355496
rect 128320 355484 128326 355496
rect 178770 355484 178776 355496
rect 128320 355456 178776 355484
rect 128320 355444 128326 355456
rect 178770 355444 178776 355456
rect 178828 355444 178834 355496
rect 128170 355376 128176 355428
rect 128228 355416 128234 355428
rect 187142 355416 187148 355428
rect 128228 355388 187148 355416
rect 128228 355376 128234 355388
rect 187142 355376 187148 355388
rect 187200 355376 187206 355428
rect 85666 355308 85672 355360
rect 85724 355348 85730 355360
rect 185670 355348 185676 355360
rect 85724 355320 185676 355348
rect 85724 355308 85730 355320
rect 185670 355308 185676 355320
rect 185728 355308 185734 355360
rect 115750 354628 115756 354680
rect 115808 354668 115814 354680
rect 171226 354668 171232 354680
rect 115808 354640 171232 354668
rect 115808 354628 115814 354640
rect 171226 354628 171232 354640
rect 171284 354668 171290 354680
rect 172422 354668 172428 354680
rect 171284 354640 172428 354668
rect 171284 354628 171290 354640
rect 172422 354628 172428 354640
rect 172480 354628 172486 354680
rect 191466 354356 191472 354408
rect 191524 354396 191530 354408
rect 197354 354396 197360 354408
rect 191524 354368 197360 354396
rect 191524 354356 191530 354368
rect 197354 354356 197360 354368
rect 197412 354356 197418 354408
rect 172422 354152 172428 354204
rect 172480 354192 172486 354204
rect 191190 354192 191196 354204
rect 172480 354164 191196 354192
rect 172480 354152 172486 354164
rect 191190 354152 191196 354164
rect 191248 354152 191254 354204
rect 129550 354084 129556 354136
rect 129608 354124 129614 354136
rect 180058 354124 180064 354136
rect 129608 354096 180064 354124
rect 129608 354084 129614 354096
rect 180058 354084 180064 354096
rect 180116 354084 180122 354136
rect 125410 354016 125416 354068
rect 125468 354056 125474 354068
rect 195422 354056 195428 354068
rect 125468 354028 195428 354056
rect 125468 354016 125474 354028
rect 195422 354016 195428 354028
rect 195480 354016 195486 354068
rect 88242 353948 88248 354000
rect 88300 353988 88306 354000
rect 173710 353988 173716 354000
rect 88300 353960 173716 353988
rect 88300 353948 88306 353960
rect 173710 353948 173716 353960
rect 173768 353948 173774 354000
rect 180242 353200 180248 353252
rect 180300 353240 180306 353252
rect 197354 353240 197360 353252
rect 180300 353212 197360 353240
rect 180300 353200 180306 353212
rect 197354 353200 197360 353212
rect 197412 353200 197418 353252
rect 111610 352588 111616 352640
rect 111668 352628 111674 352640
rect 167730 352628 167736 352640
rect 111668 352600 167736 352628
rect 111668 352588 111674 352600
rect 167730 352588 167736 352600
rect 167788 352588 167794 352640
rect 75822 352520 75828 352572
rect 75880 352560 75886 352572
rect 174906 352560 174912 352572
rect 75880 352532 174912 352560
rect 75880 352520 75886 352532
rect 174906 352520 174912 352532
rect 174964 352520 174970 352572
rect 176286 351840 176292 351892
rect 176344 351880 176350 351892
rect 197354 351880 197360 351892
rect 176344 351852 197360 351880
rect 176344 351840 176350 351852
rect 197354 351840 197360 351852
rect 197412 351840 197418 351892
rect 559650 351840 559656 351892
rect 559708 351880 559714 351892
rect 566458 351880 566464 351892
rect 559708 351852 566464 351880
rect 559708 351840 559714 351852
rect 566458 351840 566464 351852
rect 566516 351840 566522 351892
rect 130930 351364 130936 351416
rect 130988 351404 130994 351416
rect 170858 351404 170864 351416
rect 130988 351376 170864 351404
rect 130988 351364 130994 351376
rect 170858 351364 170864 351376
rect 170916 351364 170922 351416
rect 124030 351296 124036 351348
rect 124088 351336 124094 351348
rect 172330 351336 172336 351348
rect 124088 351308 172336 351336
rect 124088 351296 124094 351308
rect 172330 351296 172336 351308
rect 172388 351296 172394 351348
rect 118510 351228 118516 351280
rect 118568 351268 118574 351280
rect 195330 351268 195336 351280
rect 118568 351240 195336 351268
rect 118568 351228 118574 351240
rect 195330 351228 195336 351240
rect 195388 351268 195394 351280
rect 198826 351268 198832 351280
rect 195388 351240 198832 351268
rect 195388 351228 195394 351240
rect 198826 351228 198832 351240
rect 198884 351228 198890 351280
rect 99282 351160 99288 351212
rect 99340 351200 99346 351212
rect 181898 351200 181904 351212
rect 99340 351172 181904 351200
rect 99340 351160 99346 351172
rect 181898 351160 181904 351172
rect 181956 351160 181962 351212
rect 112990 350480 112996 350532
rect 113048 350520 113054 350532
rect 173986 350520 173992 350532
rect 113048 350492 173992 350520
rect 113048 350480 113054 350492
rect 173986 350480 173992 350492
rect 174044 350520 174050 350532
rect 175182 350520 175188 350532
rect 174044 350492 175188 350520
rect 174044 350480 174050 350492
rect 175182 350480 175188 350492
rect 175240 350480 175246 350532
rect 185762 350480 185768 350532
rect 185820 350520 185826 350532
rect 197354 350520 197360 350532
rect 185820 350492 197360 350520
rect 185820 350480 185826 350492
rect 197354 350480 197360 350492
rect 197412 350480 197418 350532
rect 175182 350004 175188 350056
rect 175240 350044 175246 350056
rect 183554 350044 183560 350056
rect 175240 350016 183560 350044
rect 175240 350004 175246 350016
rect 183554 350004 183560 350016
rect 183612 350004 183618 350056
rect 137922 349936 137928 349988
rect 137980 349976 137986 349988
rect 190454 349976 190460 349988
rect 137980 349948 190460 349976
rect 137980 349936 137986 349948
rect 190454 349936 190460 349948
rect 190512 349936 190518 349988
rect 115842 349868 115848 349920
rect 115900 349908 115906 349920
rect 176286 349908 176292 349920
rect 115900 349880 176292 349908
rect 115900 349868 115906 349880
rect 176286 349868 176292 349880
rect 176344 349868 176350 349920
rect 93762 349800 93768 349852
rect 93820 349840 93826 349852
rect 182910 349840 182916 349852
rect 93820 349812 182916 349840
rect 93820 349800 93826 349812
rect 182910 349800 182916 349812
rect 182968 349800 182974 349852
rect 174814 349052 174820 349104
rect 174872 349092 174878 349104
rect 197354 349092 197360 349104
rect 174872 349064 197360 349092
rect 174872 349052 174878 349064
rect 197354 349052 197360 349064
rect 197412 349052 197418 349104
rect 192662 348984 192668 349036
rect 192720 349024 192726 349036
rect 197446 349024 197452 349036
rect 192720 348996 197452 349024
rect 192720 348984 192726 348996
rect 197446 348984 197452 348996
rect 197504 348984 197510 349036
rect 148962 348508 148968 348560
rect 149020 348548 149026 348560
rect 178954 348548 178960 348560
rect 149020 348520 178960 348548
rect 149020 348508 149026 348520
rect 178954 348508 178960 348520
rect 179012 348508 179018 348560
rect 113082 348440 113088 348492
rect 113140 348480 113146 348492
rect 179046 348480 179052 348492
rect 113140 348452 179052 348480
rect 113140 348440 113146 348452
rect 179046 348440 179052 348452
rect 179104 348440 179110 348492
rect 78582 348372 78588 348424
rect 78640 348412 78646 348424
rect 188338 348412 188344 348424
rect 78640 348384 188344 348412
rect 78640 348372 78646 348384
rect 188338 348372 188344 348384
rect 188396 348372 188402 348424
rect 108942 347692 108948 347744
rect 109000 347732 109006 347744
rect 169846 347732 169852 347744
rect 109000 347704 169852 347732
rect 109000 347692 109006 347704
rect 169846 347692 169852 347704
rect 169904 347692 169910 347744
rect 168282 347624 168288 347676
rect 168340 347664 168346 347676
rect 197354 347664 197360 347676
rect 168340 347636 197360 347664
rect 168340 347624 168346 347636
rect 197354 347624 197360 347636
rect 197412 347624 197418 347676
rect 169846 347216 169852 347268
rect 169904 347256 169910 347268
rect 185026 347256 185032 347268
rect 169904 347228 185032 347256
rect 169904 347216 169910 347228
rect 185026 347216 185032 347228
rect 185084 347216 185090 347268
rect 129642 347148 129648 347200
rect 129700 347188 129706 347200
rect 182174 347188 182180 347200
rect 129700 347160 182180 347188
rect 129700 347148 129706 347160
rect 182174 347148 182180 347160
rect 182232 347148 182238 347200
rect 118602 347080 118608 347132
rect 118660 347120 118666 347132
rect 174814 347120 174820 347132
rect 118660 347092 174820 347120
rect 118660 347080 118666 347092
rect 174814 347080 174820 347092
rect 174872 347080 174878 347132
rect 100662 347012 100668 347064
rect 100720 347052 100726 347064
rect 180242 347052 180248 347064
rect 100720 347024 180248 347052
rect 100720 347012 100726 347024
rect 180242 347012 180248 347024
rect 180300 347012 180306 347064
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 187510 346372 187516 346384
rect 3384 346344 187516 346372
rect 3384 346332 3390 346344
rect 187510 346332 187516 346344
rect 187568 346332 187574 346384
rect 117222 346264 117228 346316
rect 117280 346304 117286 346316
rect 172514 346304 172520 346316
rect 117280 346276 172520 346304
rect 117280 346264 117286 346276
rect 172514 346264 172520 346276
rect 172572 346304 172578 346316
rect 173802 346304 173808 346316
rect 172572 346276 173808 346304
rect 172572 346264 172578 346276
rect 173802 346264 173808 346276
rect 173860 346264 173866 346316
rect 183002 346264 183008 346316
rect 183060 346304 183066 346316
rect 197354 346304 197360 346316
rect 183060 346276 197360 346304
rect 183060 346264 183066 346276
rect 197354 346264 197360 346276
rect 197412 346264 197418 346316
rect 139210 345720 139216 345772
rect 139268 345760 139274 345772
rect 189074 345760 189080 345772
rect 139268 345732 189080 345760
rect 139268 345720 139274 345732
rect 189074 345720 189080 345732
rect 189132 345720 189138 345772
rect 84102 345652 84108 345704
rect 84160 345692 84166 345704
rect 172422 345692 172428 345704
rect 84160 345664 172428 345692
rect 84160 345652 84166 345664
rect 172422 345652 172428 345664
rect 172480 345652 172486 345704
rect 173802 345652 173808 345704
rect 173860 345692 173866 345704
rect 198734 345692 198740 345704
rect 173860 345664 198740 345692
rect 173860 345652 173866 345664
rect 198734 345652 198740 345664
rect 198792 345652 198798 345704
rect 143442 344972 143448 345024
rect 143500 345012 143506 345024
rect 179230 345012 179236 345024
rect 143500 344984 179236 345012
rect 143500 344972 143506 344984
rect 179230 344972 179236 344984
rect 179288 344972 179294 345024
rect 189902 344972 189908 345024
rect 189960 345012 189966 345024
rect 197354 345012 197360 345024
rect 189960 344984 197360 345012
rect 189960 344972 189966 344984
rect 197354 344972 197360 344984
rect 197412 344972 197418 345024
rect 121270 344428 121276 344480
rect 121328 344468 121334 344480
rect 173618 344468 173624 344480
rect 121328 344440 173624 344468
rect 121328 344428 121334 344440
rect 173618 344428 173624 344440
rect 173676 344428 173682 344480
rect 125502 344360 125508 344412
rect 125560 344400 125566 344412
rect 186314 344400 186320 344412
rect 125560 344372 186320 344400
rect 125560 344360 125566 344372
rect 186314 344360 186320 344372
rect 186372 344360 186378 344412
rect 106182 344292 106188 344344
rect 106240 344332 106246 344344
rect 167914 344332 167920 344344
rect 106240 344304 167920 344332
rect 106240 344292 106246 344304
rect 167914 344292 167920 344304
rect 167972 344292 167978 344344
rect 179230 344292 179236 344344
rect 179288 344332 179294 344344
rect 186958 344332 186964 344344
rect 179288 344304 186964 344332
rect 179288 344292 179294 344304
rect 186958 344292 186964 344304
rect 187016 344292 187022 344344
rect 191374 343544 191380 343596
rect 191432 343584 191438 343596
rect 197354 343584 197360 343596
rect 191432 343556 197360 343584
rect 191432 343544 191438 343556
rect 197354 343544 197360 343556
rect 197412 343544 197418 343596
rect 560202 343544 560208 343596
rect 560260 343584 560266 343596
rect 570690 343584 570696 343596
rect 560260 343556 570696 343584
rect 560260 343544 560266 343556
rect 570690 343544 570696 343556
rect 570748 343544 570754 343596
rect 131022 342932 131028 342984
rect 131080 342972 131086 342984
rect 177482 342972 177488 342984
rect 131080 342944 177488 342972
rect 131080 342932 131086 342944
rect 177482 342932 177488 342944
rect 177540 342932 177546 342984
rect 91002 342864 91008 342916
rect 91060 342904 91066 342916
rect 184474 342904 184480 342916
rect 91060 342876 184480 342904
rect 91060 342864 91066 342876
rect 184474 342864 184480 342876
rect 184532 342864 184538 342916
rect 142062 342184 142068 342236
rect 142120 342224 142126 342236
rect 187326 342224 187332 342236
rect 142120 342196 187332 342224
rect 142120 342184 142126 342196
rect 187326 342184 187332 342196
rect 187384 342184 187390 342236
rect 192570 342184 192576 342236
rect 192628 342224 192634 342236
rect 197354 342224 197360 342236
rect 192628 342196 197360 342224
rect 192628 342184 192634 342196
rect 197354 342184 197360 342196
rect 197412 342184 197418 342236
rect 122742 341504 122748 341556
rect 122800 341544 122806 341556
rect 176194 341544 176200 341556
rect 122800 341516 176200 341544
rect 122800 341504 122806 341516
rect 176194 341504 176200 341516
rect 176252 341504 176258 341556
rect 29822 340892 29828 340944
rect 29880 340932 29886 340944
rect 46934 340932 46940 340944
rect 29880 340904 46940 340932
rect 29880 340892 29886 340904
rect 46934 340892 46940 340904
rect 46992 340892 46998 340944
rect 187326 340892 187332 340944
rect 187384 340932 187390 340944
rect 187786 340932 187792 340944
rect 187384 340904 187792 340932
rect 187384 340892 187390 340904
rect 187786 340892 187792 340904
rect 187844 340892 187850 340944
rect 114462 340824 114468 340876
rect 114520 340864 114526 340876
rect 171134 340864 171140 340876
rect 114520 340836 171140 340864
rect 114520 340824 114526 340836
rect 171134 340824 171140 340836
rect 171192 340864 171198 340876
rect 171686 340864 171692 340876
rect 171192 340836 171692 340864
rect 171192 340824 171198 340836
rect 171686 340824 171692 340836
rect 171744 340824 171750 340876
rect 181714 340824 181720 340876
rect 181772 340864 181778 340876
rect 197354 340864 197360 340876
rect 181772 340836 197360 340864
rect 181772 340824 181778 340836
rect 197354 340824 197360 340836
rect 197412 340824 197418 340876
rect 171686 340416 171692 340468
rect 171744 340456 171750 340468
rect 181622 340456 181628 340468
rect 171744 340428 181628 340456
rect 171744 340416 171750 340428
rect 181622 340416 181628 340428
rect 181680 340416 181686 340468
rect 135162 340348 135168 340400
rect 135220 340388 135226 340400
rect 181530 340388 181536 340400
rect 135220 340360 181536 340388
rect 135220 340348 135226 340360
rect 181530 340348 181536 340360
rect 181588 340348 181594 340400
rect 68922 340280 68928 340332
rect 68980 340320 68986 340332
rect 176838 340320 176844 340332
rect 68980 340292 176844 340320
rect 68980 340280 68986 340292
rect 176838 340280 176844 340292
rect 176896 340280 176902 340332
rect 29546 340212 29552 340264
rect 29604 340252 29610 340264
rect 46198 340252 46204 340264
rect 29604 340224 46204 340252
rect 29604 340212 29610 340224
rect 46198 340212 46204 340224
rect 46256 340212 46262 340264
rect 66162 340212 66168 340264
rect 66220 340252 66226 340264
rect 194870 340252 194876 340264
rect 66220 340224 194876 340252
rect 66220 340212 66226 340224
rect 194870 340212 194876 340224
rect 194928 340212 194934 340264
rect 3970 340144 3976 340196
rect 4028 340184 4034 340196
rect 197078 340184 197084 340196
rect 4028 340156 197084 340184
rect 4028 340144 4034 340156
rect 197078 340144 197084 340156
rect 197136 340144 197142 340196
rect 28534 339532 28540 339584
rect 28592 339572 28598 339584
rect 35158 339572 35164 339584
rect 28592 339544 35164 339572
rect 28592 339532 28598 339544
rect 35158 339532 35164 339544
rect 35216 339532 35222 339584
rect 60642 339396 60648 339448
rect 60700 339436 60706 339448
rect 197354 339436 197360 339448
rect 60700 339408 197360 339436
rect 60700 339396 60706 339408
rect 197354 339396 197360 339408
rect 197412 339396 197418 339448
rect 121178 339328 121184 339380
rect 121236 339368 121242 339380
rect 184566 339368 184572 339380
rect 121236 339340 184572 339368
rect 121236 339328 121242 339340
rect 184566 339328 184572 339340
rect 184624 339368 184630 339380
rect 184842 339368 184848 339380
rect 184624 339340 184848 339368
rect 184624 339328 184630 339340
rect 184842 339328 184848 339340
rect 184900 339328 184906 339380
rect 71682 338988 71688 339040
rect 71740 339028 71746 339040
rect 168006 339028 168012 339040
rect 71740 339000 168012 339028
rect 71740 338988 71746 339000
rect 168006 338988 168012 339000
rect 168064 338988 168070 339040
rect 81342 338920 81348 338972
rect 81400 338960 81406 338972
rect 187234 338960 187240 338972
rect 81400 338932 187240 338960
rect 81400 338920 81406 338932
rect 187234 338920 187240 338932
rect 187292 338920 187298 338972
rect 4062 338852 4068 338904
rect 4120 338892 4126 338904
rect 172238 338892 172244 338904
rect 4120 338864 172244 338892
rect 4120 338852 4126 338864
rect 172238 338852 172244 338864
rect 172296 338852 172302 338904
rect 3878 338784 3884 338836
rect 3936 338824 3942 338836
rect 173526 338824 173532 338836
rect 3936 338796 173532 338824
rect 3936 338784 3942 338796
rect 173526 338784 173532 338796
rect 173584 338784 173590 338836
rect 184842 338784 184848 338836
rect 184900 338824 184906 338836
rect 196802 338824 196808 338836
rect 184900 338796 196808 338824
rect 184900 338784 184906 338796
rect 196802 338784 196808 338796
rect 196860 338784 196866 338836
rect 3786 338716 3792 338768
rect 3844 338756 3850 338768
rect 196986 338756 196992 338768
rect 3844 338728 196992 338756
rect 3844 338716 3850 338728
rect 196986 338716 196992 338728
rect 197044 338716 197050 338768
rect 166258 338036 166264 338088
rect 166316 338076 166322 338088
rect 197354 338076 197360 338088
rect 166316 338048 197360 338076
rect 166316 338036 166322 338048
rect 197354 338036 197360 338048
rect 197412 338036 197418 338088
rect 176838 336676 176844 336728
rect 176896 336716 176902 336728
rect 197354 336716 197360 336728
rect 176896 336688 197360 336716
rect 176896 336676 176902 336688
rect 197354 336676 197360 336688
rect 197412 336676 197418 336728
rect 194870 336608 194876 336660
rect 194928 336648 194934 336660
rect 197446 336648 197452 336660
rect 194928 336620 197452 336648
rect 194928 336608 194934 336620
rect 197446 336608 197452 336620
rect 197504 336608 197510 336660
rect 168006 335248 168012 335300
rect 168064 335288 168070 335300
rect 197354 335288 197360 335300
rect 168064 335260 197360 335288
rect 168064 335248 168070 335260
rect 197354 335248 197360 335260
rect 197412 335248 197418 335300
rect 560202 335248 560208 335300
rect 560260 335288 560266 335300
rect 578970 335288 578976 335300
rect 560260 335260 578976 335288
rect 560260 335248 560266 335260
rect 578970 335248 578976 335260
rect 579028 335248 579034 335300
rect 176378 333888 176384 333940
rect 176436 333928 176442 333940
rect 197354 333928 197360 333940
rect 176436 333900 197360 333928
rect 176436 333888 176442 333900
rect 197354 333888 197360 333900
rect 197412 333888 197418 333940
rect 174906 332528 174912 332580
rect 174964 332568 174970 332580
rect 197354 332568 197360 332580
rect 174964 332540 197360 332568
rect 174964 332528 174970 332540
rect 197354 332528 197360 332540
rect 197412 332528 197418 332580
rect 188338 331168 188344 331220
rect 188396 331208 188402 331220
rect 197354 331208 197360 331220
rect 188396 331180 197360 331208
rect 188396 331168 188402 331180
rect 197354 331168 197360 331180
rect 197412 331168 197418 331220
rect 187234 329740 187240 329792
rect 187292 329780 187298 329792
rect 197354 329780 197360 329792
rect 187292 329752 197360 329780
rect 187292 329740 187298 329752
rect 197354 329740 197360 329752
rect 197412 329740 197418 329792
rect 172422 328380 172428 328432
rect 172480 328420 172486 328432
rect 197354 328420 197360 328432
rect 172480 328392 197360 328420
rect 172480 328380 172486 328392
rect 197354 328380 197360 328392
rect 197412 328380 197418 328432
rect 559926 328380 559932 328432
rect 559984 328420 559990 328432
rect 565170 328420 565176 328432
rect 559984 328392 565176 328420
rect 559984 328380 559990 328392
rect 565170 328380 565176 328392
rect 565228 328380 565234 328432
rect 185670 327020 185676 327072
rect 185728 327060 185734 327072
rect 197354 327060 197360 327072
rect 185728 327032 197360 327060
rect 185728 327020 185734 327032
rect 197354 327020 197360 327032
rect 197412 327020 197418 327072
rect 173710 325592 173716 325644
rect 173768 325632 173774 325644
rect 197354 325632 197360 325644
rect 173768 325604 197360 325632
rect 173768 325592 173774 325604
rect 197354 325592 197360 325604
rect 197412 325592 197418 325644
rect 565078 324300 565084 324352
rect 565136 324340 565142 324352
rect 580074 324340 580080 324352
rect 565136 324312 580080 324340
rect 565136 324300 565142 324312
rect 580074 324300 580080 324312
rect 580132 324300 580138 324352
rect 182910 324232 182916 324284
rect 182968 324272 182974 324284
rect 197446 324272 197452 324284
rect 182968 324244 197452 324272
rect 182968 324232 182974 324244
rect 197446 324232 197452 324244
rect 197504 324232 197510 324284
rect 184474 324164 184480 324216
rect 184532 324204 184538 324216
rect 197354 324204 197360 324216
rect 184532 324176 197360 324204
rect 184532 324164 184538 324176
rect 197354 324164 197360 324176
rect 197412 324164 197418 324216
rect 167822 322872 167828 322924
rect 167880 322912 167886 322924
rect 197354 322912 197360 322924
rect 167880 322884 197360 322912
rect 167880 322872 167886 322884
rect 197354 322872 197360 322884
rect 197412 322872 197418 322924
rect 181898 321512 181904 321564
rect 181956 321552 181962 321564
rect 197354 321552 197360 321564
rect 181956 321524 197360 321552
rect 181956 321512 181962 321524
rect 197354 321512 197360 321524
rect 197412 321512 197418 321564
rect 180242 320084 180248 320136
rect 180300 320124 180306 320136
rect 197354 320124 197360 320136
rect 180300 320096 197360 320124
rect 180300 320084 180306 320096
rect 197354 320084 197360 320096
rect 197412 320084 197418 320136
rect 559374 320084 559380 320136
rect 559432 320124 559438 320136
rect 566550 320124 566556 320136
rect 559432 320096 566556 320124
rect 559432 320084 559438 320096
rect 566550 320084 566556 320096
rect 566608 320084 566614 320136
rect 167638 318724 167644 318776
rect 167696 318764 167702 318776
rect 197354 318764 197360 318776
rect 167696 318736 197360 318764
rect 167696 318724 167702 318736
rect 197354 318724 197360 318736
rect 197412 318724 197418 318776
rect 167914 317364 167920 317416
rect 167972 317404 167978 317416
rect 197354 317404 197360 317416
rect 167972 317376 197360 317404
rect 167972 317364 167978 317376
rect 197354 317364 197360 317376
rect 197412 317364 197418 317416
rect 177298 315936 177304 315988
rect 177356 315976 177362 315988
rect 197354 315976 197360 315988
rect 177356 315948 197360 315976
rect 177356 315936 177362 315948
rect 197354 315936 197360 315948
rect 197412 315936 197418 315988
rect 167730 314576 167736 314628
rect 167788 314616 167794 314628
rect 197354 314616 197360 314628
rect 167788 314588 197360 314616
rect 167788 314576 167794 314588
rect 197354 314576 197360 314588
rect 197412 314576 197418 314628
rect 176286 313216 176292 313268
rect 176344 313256 176350 313268
rect 197446 313256 197452 313268
rect 176344 313228 197452 313256
rect 176344 313216 176350 313228
rect 197446 313216 197452 313228
rect 197504 313216 197510 313268
rect 179046 313148 179052 313200
rect 179104 313188 179110 313200
rect 197354 313188 197360 313200
rect 179104 313160 197360 313188
rect 179104 313148 179110 313160
rect 197354 313148 197360 313160
rect 197412 313148 197418 313200
rect 577498 311856 577504 311908
rect 577556 311896 577562 311908
rect 580442 311896 580448 311908
rect 577556 311868 580448 311896
rect 577556 311856 577562 311868
rect 580442 311856 580448 311868
rect 580500 311856 580506 311908
rect 174814 311788 174820 311840
rect 174872 311828 174878 311840
rect 197354 311828 197360 311840
rect 174872 311800 197360 311828
rect 174872 311788 174878 311800
rect 197354 311788 197360 311800
rect 197412 311788 197418 311840
rect 560202 311788 560208 311840
rect 560260 311828 560266 311840
rect 577590 311828 577596 311840
rect 560260 311800 577596 311828
rect 560260 311788 560266 311800
rect 577590 311788 577596 311800
rect 577648 311788 577654 311840
rect 173618 310428 173624 310480
rect 173676 310468 173682 310480
rect 197354 310468 197360 310480
rect 173676 310440 197360 310468
rect 173676 310428 173682 310440
rect 197354 310428 197360 310440
rect 197412 310428 197418 310480
rect 172330 309068 172336 309120
rect 172388 309108 172394 309120
rect 197354 309108 197360 309120
rect 172388 309080 197360 309108
rect 172388 309068 172394 309080
rect 197354 309068 197360 309080
rect 197412 309068 197418 309120
rect 195422 307708 195428 307760
rect 195480 307748 195486 307760
rect 197722 307748 197728 307760
rect 195480 307720 197728 307748
rect 195480 307708 195486 307720
rect 197722 307708 197728 307720
rect 197780 307708 197786 307760
rect 187142 306280 187148 306332
rect 187200 306320 187206 306332
rect 197354 306320 197360 306332
rect 187200 306292 197360 306320
rect 187200 306280 187206 306292
rect 197354 306280 197360 306292
rect 197412 306280 197418 306332
rect 177482 304920 177488 304972
rect 177540 304960 177546 304972
rect 197354 304960 197360 304972
rect 177540 304932 197360 304960
rect 177540 304920 177546 304932
rect 197354 304920 197360 304932
rect 197412 304920 197418 304972
rect 181806 303560 181812 303612
rect 181864 303600 181870 303612
rect 197354 303600 197360 303612
rect 181864 303572 197360 303600
rect 181864 303560 181870 303572
rect 197354 303560 197360 303572
rect 197412 303560 197418 303612
rect 559282 303424 559288 303476
rect 559340 303464 559346 303476
rect 561030 303464 561036 303476
rect 559340 303436 561036 303464
rect 559340 303424 559346 303436
rect 561030 303424 561036 303436
rect 561088 303424 561094 303476
rect 174722 302132 174728 302184
rect 174780 302172 174786 302184
rect 197354 302172 197360 302184
rect 174780 302144 197360 302172
rect 174780 302132 174786 302144
rect 197354 302132 197360 302144
rect 197412 302132 197418 302184
rect 180334 300772 180340 300824
rect 180392 300812 180398 300824
rect 197354 300812 197360 300824
rect 180392 300784 197360 300812
rect 180392 300772 180398 300784
rect 197354 300772 197360 300784
rect 197412 300772 197418 300824
rect 173526 299480 173532 299532
rect 173584 299520 173590 299532
rect 197354 299520 197360 299532
rect 173584 299492 197360 299520
rect 173584 299480 173590 299492
rect 197354 299480 197360 299492
rect 197412 299480 197418 299532
rect 174722 298120 174728 298172
rect 174780 298160 174786 298172
rect 197354 298160 197360 298172
rect 174780 298132 197360 298160
rect 174780 298120 174786 298132
rect 197354 298120 197360 298132
rect 197412 298120 197418 298172
rect 560938 298120 560944 298172
rect 560996 298160 561002 298172
rect 580166 298160 580172 298172
rect 560996 298132 580172 298160
rect 560996 298120 561002 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 167638 296692 167644 296744
rect 167696 296732 167702 296744
rect 197354 296732 197360 296744
rect 167696 296704 197360 296732
rect 167696 296692 167702 296704
rect 197354 296692 197360 296704
rect 197412 296692 197418 296744
rect 559006 296624 559012 296676
rect 559064 296664 559070 296676
rect 580350 296664 580356 296676
rect 559064 296636 580356 296664
rect 559064 296624 559070 296636
rect 580350 296624 580356 296636
rect 580408 296624 580414 296676
rect 177298 295332 177304 295384
rect 177356 295372 177362 295384
rect 197354 295372 197360 295384
rect 177356 295344 197360 295372
rect 177356 295332 177362 295344
rect 197354 295332 197360 295344
rect 197412 295332 197418 295384
rect 172238 293972 172244 294024
rect 172296 294012 172302 294024
rect 197354 294012 197360 294024
rect 172296 293984 197360 294012
rect 172296 293972 172302 293984
rect 197354 293972 197360 293984
rect 197412 293972 197418 294024
rect 173618 292544 173624 292596
rect 173676 292584 173682 292596
rect 197354 292584 197360 292596
rect 173676 292556 197360 292584
rect 173676 292544 173682 292556
rect 197354 292544 197360 292556
rect 197412 292544 197418 292596
rect 167730 291184 167736 291236
rect 167788 291224 167794 291236
rect 197354 291224 197360 291236
rect 167788 291196 197360 291224
rect 167788 291184 167794 291196
rect 197354 291184 197360 291196
rect 197412 291184 197418 291236
rect 180242 289824 180248 289876
rect 180300 289864 180306 289876
rect 197354 289864 197360 289876
rect 180300 289836 197360 289864
rect 180300 289824 180306 289836
rect 197354 289824 197360 289836
rect 197412 289824 197418 289876
rect 174814 288396 174820 288448
rect 174872 288436 174878 288448
rect 197354 288436 197360 288448
rect 174872 288408 197360 288436
rect 174872 288396 174878 288408
rect 197354 288396 197360 288408
rect 197412 288396 197418 288448
rect 560202 288328 560208 288380
rect 560260 288368 560266 288380
rect 567930 288368 567936 288380
rect 560260 288340 567936 288368
rect 560260 288328 560266 288340
rect 567930 288328 567936 288340
rect 567988 288328 567994 288380
rect 176286 287104 176292 287156
rect 176344 287144 176350 287156
rect 197446 287144 197452 287156
rect 176344 287116 197452 287144
rect 176344 287104 176350 287116
rect 197446 287104 197452 287116
rect 197504 287104 197510 287156
rect 167914 287036 167920 287088
rect 167972 287076 167978 287088
rect 197354 287076 197360 287088
rect 167972 287048 197360 287076
rect 167972 287036 167978 287048
rect 197354 287036 197360 287048
rect 197412 287036 197418 287088
rect 172330 285676 172336 285728
rect 172388 285716 172394 285728
rect 197354 285716 197360 285728
rect 172388 285688 197360 285716
rect 172388 285676 172394 285688
rect 197354 285676 197360 285688
rect 197412 285676 197418 285728
rect 168006 284316 168012 284368
rect 168064 284356 168070 284368
rect 197354 284356 197360 284368
rect 168064 284328 197360 284356
rect 168064 284316 168070 284328
rect 197354 284316 197360 284328
rect 197412 284316 197418 284368
rect 168098 282888 168104 282940
rect 168156 282928 168162 282940
rect 197354 282928 197360 282940
rect 168156 282900 197360 282928
rect 168156 282888 168162 282900
rect 197354 282888 197360 282900
rect 197412 282888 197418 282940
rect 181714 281528 181720 281580
rect 181772 281568 181778 281580
rect 197354 281568 197360 281580
rect 181772 281540 197360 281568
rect 181772 281528 181778 281540
rect 197354 281528 197360 281540
rect 197412 281528 197418 281580
rect 167822 280168 167828 280220
rect 167880 280208 167886 280220
rect 197354 280208 197360 280220
rect 167880 280180 197360 280208
rect 167880 280168 167886 280180
rect 197354 280168 197360 280180
rect 197412 280168 197418 280220
rect 559926 280100 559932 280152
rect 559984 280140 559990 280152
rect 574830 280140 574836 280152
rect 559984 280112 574836 280140
rect 559984 280100 559990 280112
rect 574830 280100 574836 280112
rect 574888 280100 574894 280152
rect 168190 278740 168196 278792
rect 168248 278780 168254 278792
rect 197354 278780 197360 278792
rect 168248 278752 197360 278780
rect 168248 278740 168254 278752
rect 197354 278740 197360 278752
rect 197412 278740 197418 278792
rect 177482 277380 177488 277432
rect 177540 277420 177546 277432
rect 197354 277420 197360 277432
rect 177540 277392 197360 277420
rect 177540 277380 177546 277392
rect 197354 277380 197360 277392
rect 197412 277380 197418 277432
rect 174906 276088 174912 276140
rect 174964 276128 174970 276140
rect 197354 276128 197360 276140
rect 174964 276100 197360 276128
rect 174964 276088 174970 276100
rect 197354 276088 197360 276100
rect 197412 276088 197418 276140
rect 173710 276020 173716 276072
rect 173768 276060 173774 276072
rect 197446 276060 197452 276072
rect 173768 276032 197452 276060
rect 173768 276020 173774 276032
rect 197446 276020 197452 276032
rect 197504 276020 197510 276072
rect 172422 274660 172428 274712
rect 172480 274700 172486 274712
rect 197354 274700 197360 274712
rect 172480 274672 197360 274700
rect 172480 274660 172486 274672
rect 197354 274660 197360 274672
rect 197412 274660 197418 274712
rect 180334 273232 180340 273284
rect 180392 273272 180398 273284
rect 197354 273272 197360 273284
rect 180392 273244 197360 273272
rect 180392 273232 180398 273244
rect 197354 273232 197360 273244
rect 197412 273232 197418 273284
rect 171042 271872 171048 271924
rect 171100 271912 171106 271924
rect 197354 271912 197360 271924
rect 171100 271884 197360 271912
rect 171100 271872 171106 271884
rect 197354 271872 197360 271884
rect 197412 271872 197418 271924
rect 566458 271872 566464 271924
rect 566516 271912 566522 271924
rect 579798 271912 579804 271924
rect 566516 271884 579804 271912
rect 566516 271872 566522 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 187142 270512 187148 270564
rect 187200 270552 187206 270564
rect 197354 270552 197360 270564
rect 187200 270524 197360 270552
rect 187200 270512 187206 270524
rect 197354 270512 197360 270524
rect 197412 270512 197418 270564
rect 183002 267724 183008 267776
rect 183060 267764 183066 267776
rect 197354 267764 197360 267776
rect 183060 267736 197360 267764
rect 183060 267724 183066 267736
rect 197354 267724 197360 267736
rect 197412 267724 197418 267776
rect 181806 266364 181812 266416
rect 181864 266404 181870 266416
rect 197354 266404 197360 266416
rect 181864 266376 197360 266404
rect 181864 266364 181870 266376
rect 197354 266364 197360 266376
rect 197412 266364 197418 266416
rect 179046 264936 179052 264988
rect 179104 264976 179110 264988
rect 197354 264976 197360 264988
rect 179104 264948 197360 264976
rect 179104 264936 179110 264948
rect 197354 264936 197360 264948
rect 197412 264936 197418 264988
rect 169202 264188 169208 264240
rect 169260 264228 169266 264240
rect 182910 264228 182916 264240
rect 169260 264200 182916 264228
rect 169260 264188 169266 264200
rect 182910 264188 182916 264200
rect 182968 264188 182974 264240
rect 176378 263644 176384 263696
rect 176436 263684 176442 263696
rect 197446 263684 197452 263696
rect 176436 263656 197452 263684
rect 176436 263644 176442 263656
rect 197446 263644 197452 263656
rect 197504 263644 197510 263696
rect 171686 263576 171692 263628
rect 171744 263616 171750 263628
rect 197354 263616 197360 263628
rect 171744 263588 197360 263616
rect 171744 263576 171750 263588
rect 197354 263576 197360 263588
rect 197412 263576 197418 263628
rect 560202 263508 560208 263560
rect 560260 263548 560266 263560
rect 570598 263548 570604 263560
rect 560260 263520 570604 263548
rect 560260 263508 560266 263520
rect 570598 263508 570604 263520
rect 570656 263508 570662 263560
rect 168282 262216 168288 262268
rect 168340 262256 168346 262268
rect 197354 262256 197360 262268
rect 168340 262228 197360 262256
rect 168340 262216 168346 262228
rect 197354 262216 197360 262228
rect 197412 262216 197418 262268
rect 168558 261468 168564 261520
rect 168616 261508 168622 261520
rect 195422 261508 195428 261520
rect 168616 261480 195428 261508
rect 168616 261468 168622 261480
rect 195422 261468 195428 261480
rect 195480 261468 195486 261520
rect 187234 260856 187240 260908
rect 187292 260896 187298 260908
rect 197354 260896 197360 260908
rect 187292 260868 197360 260896
rect 187292 260856 187298 260868
rect 197354 260856 197360 260868
rect 197412 260856 197418 260908
rect 169846 258068 169852 258120
rect 169904 258108 169910 258120
rect 197354 258108 197360 258120
rect 169904 258080 197360 258108
rect 169904 258068 169910 258080
rect 197354 258068 197360 258080
rect 197412 258068 197418 258120
rect 567838 258068 567844 258120
rect 567896 258108 567902 258120
rect 580166 258108 580172 258120
rect 567896 258080 580172 258108
rect 567896 258068 567902 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 560018 256640 560024 256692
rect 560076 256680 560082 256692
rect 578878 256680 578884 256692
rect 560076 256652 578884 256680
rect 560076 256640 560082 256652
rect 578878 256640 578884 256652
rect 578936 256640 578942 256692
rect 166718 254532 166724 254584
rect 166776 254572 166782 254584
rect 197814 254572 197820 254584
rect 166776 254544 197820 254572
rect 166776 254532 166782 254544
rect 197814 254532 197820 254544
rect 197872 254532 197878 254584
rect 27522 253852 27528 253904
rect 27580 253892 27586 253904
rect 197906 253892 197912 253904
rect 27580 253864 197912 253892
rect 27580 253852 27586 253864
rect 197906 253852 197912 253864
rect 197964 253852 197970 253904
rect 128078 253784 128084 253836
rect 128136 253824 128142 253836
rect 179046 253824 179052 253836
rect 128136 253796 179052 253824
rect 128136 253784 128142 253796
rect 179046 253784 179052 253796
rect 179104 253784 179110 253836
rect 115658 253716 115664 253768
rect 115716 253756 115722 253768
rect 171042 253756 171048 253768
rect 115716 253728 171048 253756
rect 115716 253716 115722 253728
rect 171042 253716 171048 253728
rect 171100 253716 171106 253768
rect 125502 253648 125508 253700
rect 125560 253688 125566 253700
rect 181806 253688 181812 253700
rect 125560 253660 181812 253688
rect 125560 253648 125566 253660
rect 181806 253648 181812 253660
rect 181864 253648 181870 253700
rect 123018 253580 123024 253632
rect 123076 253620 123082 253632
rect 183002 253620 183008 253632
rect 123076 253592 183008 253620
rect 123076 253580 123082 253592
rect 183002 253580 183008 253592
rect 183060 253580 183066 253632
rect 118326 253512 118332 253564
rect 118384 253552 118390 253564
rect 187142 253552 187148 253564
rect 118384 253524 187148 253552
rect 118384 253512 118390 253524
rect 187142 253512 187148 253524
rect 187200 253512 187206 253564
rect 98270 253444 98276 253496
rect 98328 253484 98334 253496
rect 167822 253484 167828 253496
rect 98328 253456 167828 253484
rect 98328 253444 98334 253456
rect 167822 253444 167828 253456
rect 167880 253444 167886 253496
rect 75546 253376 75552 253428
rect 75604 253416 75610 253428
rect 167730 253416 167736 253428
rect 75604 253388 167736 253416
rect 75604 253376 75610 253388
rect 167730 253376 167736 253388
rect 167788 253376 167794 253428
rect 70670 253308 70676 253360
rect 70728 253348 70734 253360
rect 172238 253348 172244 253360
rect 70728 253320 172244 253348
rect 70728 253308 70734 253320
rect 172238 253308 172244 253320
rect 172296 253308 172302 253360
rect 65702 253240 65708 253292
rect 65760 253280 65766 253292
rect 167638 253280 167644 253292
rect 65760 253252 167644 253280
rect 65760 253240 65766 253252
rect 167638 253240 167644 253252
rect 167696 253240 167702 253292
rect 28350 253172 28356 253224
rect 28408 253212 28414 253224
rect 29454 253212 29460 253224
rect 28408 253184 29460 253212
rect 28408 253172 28414 253184
rect 29454 253172 29460 253184
rect 29512 253212 29518 253224
rect 43346 253212 43352 253224
rect 29512 253184 43352 253212
rect 29512 253172 29518 253184
rect 43346 253172 43352 253184
rect 43404 253172 43410 253224
rect 60642 253172 60648 253224
rect 60700 253212 60706 253224
rect 173526 253212 173532 253224
rect 60700 253184 173532 253212
rect 60700 253172 60706 253184
rect 173526 253172 173532 253184
rect 173584 253172 173590 253224
rect 130562 253104 130568 253156
rect 130620 253144 130626 253156
rect 176378 253144 176384 253156
rect 130620 253116 176384 253144
rect 130620 253104 130626 253116
rect 176378 253104 176384 253116
rect 176436 253104 176442 253156
rect 132954 253036 132960 253088
rect 133012 253076 133018 253088
rect 171686 253076 171692 253088
rect 133012 253048 171692 253076
rect 133012 253036 133018 253048
rect 171686 253036 171692 253048
rect 171744 253036 171750 253088
rect 27062 252492 27068 252544
rect 27120 252532 27126 252544
rect 27246 252532 27252 252544
rect 27120 252504 27252 252532
rect 27120 252492 27126 252504
rect 27246 252492 27252 252504
rect 27304 252492 27310 252544
rect 28442 252492 28448 252544
rect 28500 252532 28506 252544
rect 34514 252532 34520 252544
rect 28500 252504 34520 252532
rect 28500 252492 28506 252504
rect 34514 252492 34520 252504
rect 34572 252492 34578 252544
rect 197998 252532 198004 252544
rect 35866 252504 198004 252532
rect 27264 252464 27292 252492
rect 35866 252464 35894 252504
rect 197998 252492 198004 252504
rect 198056 252492 198062 252544
rect 27264 252436 35894 252464
rect 166994 252424 167000 252476
rect 167052 252464 167058 252476
rect 197446 252464 197452 252476
rect 167052 252436 197452 252464
rect 167052 252424 167058 252436
rect 197446 252424 197452 252436
rect 197504 252424 197510 252476
rect 68186 252356 68192 252408
rect 68244 252396 68250 252408
rect 177298 252396 177304 252408
rect 68244 252368 177304 252396
rect 68244 252356 68250 252368
rect 177298 252356 177304 252368
rect 177356 252356 177362 252408
rect 189258 252356 189264 252408
rect 189316 252396 189322 252408
rect 190362 252396 190368 252408
rect 189316 252368 190368 252396
rect 189316 252356 189322 252368
rect 190362 252356 190368 252368
rect 190420 252396 190426 252408
rect 197354 252396 197360 252408
rect 190420 252368 197360 252396
rect 190420 252356 190426 252368
rect 197354 252356 197360 252368
rect 197412 252356 197418 252408
rect 78122 252288 78128 252340
rect 78180 252328 78186 252340
rect 180242 252328 180248 252340
rect 78180 252300 180248 252328
rect 78180 252288 78186 252300
rect 180242 252288 180248 252300
rect 180300 252288 180306 252340
rect 73154 252220 73160 252272
rect 73212 252260 73218 252272
rect 173618 252260 173624 252272
rect 73212 252232 173624 252260
rect 73212 252220 73218 252232
rect 173618 252220 173624 252232
rect 173676 252220 173682 252272
rect 83550 252152 83556 252204
rect 83608 252192 83614 252204
rect 176286 252192 176292 252204
rect 83608 252164 176292 252192
rect 83608 252152 83614 252164
rect 176286 252152 176292 252164
rect 176344 252152 176350 252204
rect 95602 252084 95608 252136
rect 95660 252124 95666 252136
rect 181714 252124 181720 252136
rect 95660 252096 181720 252124
rect 95660 252084 95666 252096
rect 181714 252084 181720 252096
rect 181772 252084 181778 252136
rect 85666 252016 85672 252068
rect 85724 252056 85730 252068
rect 167914 252056 167920 252068
rect 85724 252028 167920 252056
rect 85724 252016 85730 252028
rect 167914 252016 167920 252028
rect 167972 252016 167978 252068
rect 90818 251948 90824 252000
rect 90876 251988 90882 252000
rect 168006 251988 168012 252000
rect 90876 251960 168012 251988
rect 90876 251948 90882 251960
rect 168006 251948 168012 251960
rect 168064 251948 168070 252000
rect 93210 251880 93216 251932
rect 93268 251920 93274 251932
rect 168098 251920 168104 251932
rect 93268 251892 168104 251920
rect 93268 251880 93274 251892
rect 168098 251880 168104 251892
rect 168156 251880 168162 251932
rect 100570 251812 100576 251864
rect 100628 251852 100634 251864
rect 168190 251852 168196 251864
rect 100628 251824 168196 251852
rect 100628 251812 100634 251824
rect 168190 251812 168196 251824
rect 168248 251812 168254 251864
rect 174998 251812 175004 251864
rect 175056 251852 175062 251864
rect 189258 251852 189264 251864
rect 175056 251824 189264 251852
rect 175056 251812 175062 251824
rect 189258 251812 189264 251824
rect 189316 251812 189322 251864
rect 120902 251744 120908 251796
rect 120960 251784 120966 251796
rect 166718 251784 166724 251796
rect 120960 251756 166724 251784
rect 120960 251744 120966 251756
rect 166718 251744 166724 251756
rect 166776 251744 166782 251796
rect 166994 251744 167000 251796
rect 167052 251784 167058 251796
rect 167822 251784 167828 251796
rect 167052 251756 167828 251784
rect 167052 251744 167058 251756
rect 167822 251744 167828 251756
rect 167880 251744 167886 251796
rect 135990 251676 135996 251728
rect 136048 251716 136054 251728
rect 168282 251716 168288 251728
rect 136048 251688 168288 251716
rect 136048 251676 136054 251688
rect 168282 251676 168288 251688
rect 168340 251676 168346 251728
rect 151078 251608 151084 251660
rect 151136 251648 151142 251660
rect 166994 251648 167000 251660
rect 151136 251620 167000 251648
rect 151136 251608 151142 251620
rect 166994 251608 167000 251620
rect 167052 251608 167058 251660
rect 63402 251540 63408 251592
rect 63460 251580 63466 251592
rect 174722 251580 174728 251592
rect 63460 251552 174728 251580
rect 63460 251540 63466 251552
rect 174722 251540 174728 251552
rect 174780 251540 174786 251592
rect 81250 251132 81256 251184
rect 81308 251172 81314 251184
rect 174814 251172 174820 251184
rect 81308 251144 174820 251172
rect 81308 251132 81314 251144
rect 174814 251132 174820 251144
rect 174872 251132 174878 251184
rect 88242 251064 88248 251116
rect 88300 251104 88306 251116
rect 172330 251104 172336 251116
rect 88300 251076 172336 251104
rect 88300 251064 88306 251076
rect 172330 251064 172336 251076
rect 172388 251064 172394 251116
rect 103146 250996 103152 251048
rect 103204 251036 103210 251048
rect 177482 251036 177488 251048
rect 103204 251008 177488 251036
rect 103204 250996 103210 251008
rect 177482 250996 177488 251008
rect 177540 250996 177546 251048
rect 106090 250928 106096 250980
rect 106148 250968 106154 250980
rect 173710 250968 173716 250980
rect 106148 250940 173716 250968
rect 106148 250928 106154 250940
rect 173710 250928 173716 250940
rect 173768 250928 173774 250980
rect 113082 250860 113088 250912
rect 113140 250900 113146 250912
rect 180334 250900 180340 250912
rect 113140 250872 180340 250900
rect 113140 250860 113146 250872
rect 180334 250860 180340 250872
rect 180392 250860 180398 250912
rect 108482 250792 108488 250844
rect 108540 250832 108546 250844
rect 174906 250832 174912 250844
rect 108540 250804 174912 250832
rect 108540 250792 108546 250804
rect 174906 250792 174912 250804
rect 174964 250792 174970 250844
rect 110506 250724 110512 250776
rect 110564 250764 110570 250776
rect 172422 250764 172428 250776
rect 110564 250736 172428 250764
rect 110564 250724 110570 250736
rect 172422 250724 172428 250736
rect 172480 250724 172486 250776
rect 138290 250656 138296 250708
rect 138348 250696 138354 250708
rect 187234 250696 187240 250708
rect 138348 250668 187240 250696
rect 138348 250656 138354 250668
rect 187234 250656 187240 250668
rect 187292 250656 187298 250708
rect 129550 249704 129556 249756
rect 129608 249744 129614 249756
rect 193582 249744 193588 249756
rect 129608 249716 193588 249744
rect 129608 249704 129614 249716
rect 193582 249704 193588 249716
rect 193640 249704 193646 249756
rect 114370 249636 114376 249688
rect 114428 249676 114434 249688
rect 174538 249676 174544 249688
rect 114428 249648 174544 249676
rect 114428 249636 114434 249648
rect 174538 249636 174544 249648
rect 174596 249676 174602 249688
rect 175182 249676 175188 249688
rect 174596 249648 175188 249676
rect 174596 249636 174602 249648
rect 175182 249636 175188 249648
rect 175240 249636 175246 249688
rect 143350 249568 143356 249620
rect 143408 249608 143414 249620
rect 176838 249608 176844 249620
rect 143408 249580 176844 249608
rect 143408 249568 143414 249580
rect 176838 249568 176844 249580
rect 176896 249568 176902 249620
rect 193582 249160 193588 249212
rect 193640 249200 193646 249212
rect 194686 249200 194692 249212
rect 193640 249172 194692 249200
rect 193640 249160 193646 249172
rect 194686 249160 194692 249172
rect 194744 249160 194750 249212
rect 176838 249092 176844 249144
rect 176896 249132 176902 249144
rect 177390 249132 177396 249144
rect 176896 249104 177396 249132
rect 176896 249092 176902 249104
rect 177390 249092 177396 249104
rect 177448 249132 177454 249144
rect 186406 249132 186412 249144
rect 177448 249104 186412 249132
rect 177448 249092 177454 249104
rect 186406 249092 186412 249104
rect 186464 249092 186470 249144
rect 175182 249024 175188 249076
rect 175240 249064 175246 249076
rect 192018 249064 192024 249076
rect 175240 249036 192024 249064
rect 175240 249024 175246 249036
rect 192018 249024 192024 249036
rect 192076 249024 192082 249076
rect 114462 248344 114468 248396
rect 114520 248384 114526 248396
rect 176102 248384 176108 248396
rect 114520 248356 176108 248384
rect 114520 248344 114526 248356
rect 176102 248344 176108 248356
rect 176160 248344 176166 248396
rect 560202 248344 560208 248396
rect 560260 248384 560266 248396
rect 577498 248384 577504 248396
rect 560260 248356 577504 248384
rect 560260 248344 560266 248356
rect 577498 248344 577504 248356
rect 577556 248344 577562 248396
rect 132034 248276 132040 248328
rect 132092 248316 132098 248328
rect 191098 248316 191104 248328
rect 132092 248288 191104 248316
rect 132092 248276 132098 248288
rect 191098 248276 191104 248288
rect 191156 248276 191162 248328
rect 126882 248208 126888 248260
rect 126940 248248 126946 248260
rect 176654 248248 176660 248260
rect 126940 248220 176660 248248
rect 126940 248208 126946 248220
rect 176654 248208 176660 248220
rect 176712 248208 176718 248260
rect 176654 247120 176660 247172
rect 176712 247160 176718 247172
rect 177390 247160 177396 247172
rect 176712 247132 177396 247160
rect 176712 247120 176718 247132
rect 177390 247120 177396 247132
rect 177448 247120 177454 247172
rect 176102 247052 176108 247104
rect 176160 247092 176166 247104
rect 177298 247092 177304 247104
rect 176160 247064 177304 247092
rect 176160 247052 176166 247064
rect 177298 247052 177304 247064
rect 177356 247052 177362 247104
rect 191098 247052 191104 247104
rect 191156 247092 191162 247104
rect 193398 247092 193404 247104
rect 191156 247064 193404 247092
rect 191156 247052 191162 247064
rect 193398 247052 193404 247064
rect 193456 247052 193462 247104
rect 28810 246984 28816 247036
rect 28868 247024 28874 247036
rect 197354 247024 197360 247036
rect 28868 246996 197360 247024
rect 28868 246984 28874 246996
rect 197354 246984 197360 246996
rect 197412 246984 197418 247036
rect 124122 246916 124128 246968
rect 124180 246956 124186 246968
rect 179414 246956 179420 246968
rect 124180 246928 179420 246956
rect 124180 246916 124186 246928
rect 179414 246916 179420 246928
rect 179472 246916 179478 246968
rect 140682 246304 140688 246356
rect 140740 246344 140746 246356
rect 167638 246344 167644 246356
rect 140740 246316 167644 246344
rect 140740 246304 140746 246316
rect 167638 246304 167644 246316
rect 167696 246304 167702 246356
rect 179414 245624 179420 245676
rect 179472 245664 179478 245676
rect 180242 245664 180248 245676
rect 179472 245636 180248 245664
rect 179472 245624 179478 245636
rect 180242 245624 180248 245636
rect 180300 245624 180306 245676
rect 28166 245556 28172 245608
rect 28224 245596 28230 245608
rect 197354 245596 197360 245608
rect 28224 245568 197360 245596
rect 28224 245556 28230 245568
rect 197354 245556 197360 245568
rect 197412 245556 197418 245608
rect 122742 245488 122748 245540
rect 122800 245528 122806 245540
rect 169846 245528 169852 245540
rect 122800 245500 169852 245528
rect 122800 245488 122806 245500
rect 169846 245488 169852 245500
rect 169904 245488 169910 245540
rect 169846 244876 169852 244928
rect 169904 244916 169910 244928
rect 170674 244916 170680 244928
rect 169904 244888 170680 244916
rect 169904 244876 169910 244888
rect 170674 244876 170680 244888
rect 170732 244916 170738 244928
rect 180794 244916 180800 244928
rect 170732 244888 180800 244916
rect 170732 244876 170738 244888
rect 180794 244876 180800 244888
rect 180852 244876 180858 244928
rect 28534 244196 28540 244248
rect 28592 244236 28598 244248
rect 197354 244236 197360 244248
rect 28592 244208 197360 244236
rect 28592 244196 28598 244208
rect 197354 244196 197360 244208
rect 197412 244196 197418 244248
rect 112990 244128 112996 244180
rect 113048 244168 113054 244180
rect 172054 244168 172060 244180
rect 113048 244140 172060 244168
rect 113048 244128 113054 244140
rect 172054 244128 172060 244140
rect 172112 244168 172118 244180
rect 179138 244168 179144 244180
rect 172112 244140 179144 244168
rect 172112 244128 172118 244140
rect 179138 244128 179144 244140
rect 179196 244128 179202 244180
rect 143442 244060 143448 244112
rect 143500 244100 143506 244112
rect 176010 244100 176016 244112
rect 143500 244072 176016 244100
rect 143500 244060 143506 244072
rect 176010 244060 176016 244072
rect 176068 244060 176074 244112
rect 176010 243516 176016 243568
rect 176068 243556 176074 243568
rect 183646 243556 183652 243568
rect 176068 243528 183652 243556
rect 176068 243516 176074 243528
rect 183646 243516 183652 243528
rect 183704 243516 183710 243568
rect 28718 242836 28724 242888
rect 28776 242876 28782 242888
rect 197354 242876 197360 242888
rect 28776 242848 197360 242876
rect 28776 242836 28782 242848
rect 197354 242836 197360 242848
rect 197412 242836 197418 242888
rect 119982 242768 119988 242820
rect 120040 242808 120046 242820
rect 189718 242808 189724 242820
rect 120040 242780 189724 242808
rect 120040 242768 120046 242780
rect 189718 242768 189724 242780
rect 189776 242808 189782 242820
rect 189994 242808 190000 242820
rect 189776 242780 190000 242808
rect 189776 242768 189782 242780
rect 189994 242768 190000 242780
rect 190052 242768 190058 242820
rect 189994 242156 190000 242208
rect 190052 242196 190058 242208
rect 196894 242196 196900 242208
rect 190052 242168 196900 242196
rect 190052 242156 190058 242168
rect 196894 242156 196900 242168
rect 196952 242156 196958 242208
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 184382 241448 184388 241460
rect 3292 241420 184388 241448
rect 3292 241408 3298 241420
rect 184382 241408 184388 241420
rect 184440 241408 184446 241460
rect 121270 241340 121276 241392
rect 121328 241380 121334 241392
rect 173434 241380 173440 241392
rect 121328 241352 173440 241380
rect 121328 241340 121334 241352
rect 173434 241340 173440 241352
rect 173492 241380 173498 241392
rect 173802 241380 173808 241392
rect 173492 241352 173808 241380
rect 173492 241340 173498 241352
rect 173802 241340 173808 241352
rect 173860 241340 173866 241392
rect 173802 240728 173808 240780
rect 173860 240768 173866 240780
rect 191098 240768 191104 240780
rect 173860 240740 191104 240768
rect 173860 240728 173866 240740
rect 191098 240728 191104 240740
rect 191156 240728 191162 240780
rect 115842 240048 115848 240100
rect 115900 240088 115906 240100
rect 175274 240088 175280 240100
rect 115900 240060 175280 240088
rect 115900 240048 115906 240060
rect 175274 240048 175280 240060
rect 175332 240048 175338 240100
rect 129642 239980 129648 240032
rect 129700 240020 129706 240032
rect 173894 240020 173900 240032
rect 129700 239992 173900 240020
rect 129700 239980 129706 239992
rect 173894 239980 173900 239992
rect 173952 239980 173958 240032
rect 560202 239572 560208 239624
rect 560260 239612 560266 239624
rect 565078 239612 565084 239624
rect 560260 239584 565084 239612
rect 560260 239572 560266 239584
rect 565078 239572 565084 239584
rect 565136 239572 565142 239624
rect 182910 239368 182916 239420
rect 182968 239408 182974 239420
rect 195974 239408 195980 239420
rect 182968 239380 195980 239408
rect 182968 239368 182974 239380
rect 195974 239368 195980 239380
rect 196032 239368 196038 239420
rect 173894 239232 173900 239284
rect 173952 239272 173958 239284
rect 174722 239272 174728 239284
rect 173952 239244 174728 239272
rect 173952 239232 173958 239244
rect 174722 239232 174728 239244
rect 174780 239232 174786 239284
rect 195974 238892 195980 238944
rect 196032 238932 196038 238944
rect 197354 238932 197360 238944
rect 196032 238904 197360 238932
rect 196032 238892 196038 238904
rect 197354 238892 197360 238904
rect 197412 238892 197418 238944
rect 107562 238688 107568 238740
rect 107620 238728 107626 238740
rect 168190 238728 168196 238740
rect 107620 238700 168196 238728
rect 107620 238688 107626 238700
rect 168190 238688 168196 238700
rect 168248 238688 168254 238740
rect 128262 238620 128268 238672
rect 128320 238660 128326 238672
rect 187694 238660 187700 238672
rect 128320 238632 187700 238660
rect 128320 238620 128326 238632
rect 187694 238620 187700 238632
rect 187752 238620 187758 238672
rect 47578 238008 47584 238060
rect 47636 238048 47642 238060
rect 174998 238048 175004 238060
rect 47636 238020 175004 238048
rect 47636 238008 47642 238020
rect 174998 238008 175004 238020
rect 175056 238008 175062 238060
rect 178678 238008 178684 238060
rect 178736 238048 178742 238060
rect 197354 238048 197360 238060
rect 178736 238020 197360 238048
rect 178736 238008 178742 238020
rect 197354 238008 197360 238020
rect 197412 238008 197418 238060
rect 168190 237396 168196 237448
rect 168248 237436 168254 237448
rect 185578 237436 185584 237448
rect 168248 237408 185584 237436
rect 168248 237396 168254 237408
rect 185578 237396 185584 237408
rect 185636 237396 185642 237448
rect 117222 237328 117228 237380
rect 117280 237368 117286 237380
rect 174078 237368 174084 237380
rect 117280 237340 174084 237368
rect 117280 237328 117286 237340
rect 174078 237328 174084 237340
rect 174136 237328 174142 237380
rect 142062 237260 142068 237312
rect 142120 237300 142126 237312
rect 175918 237300 175924 237312
rect 142120 237272 175924 237300
rect 142120 237260 142126 237272
rect 175918 237260 175924 237272
rect 175976 237260 175982 237312
rect 175918 236716 175924 236768
rect 175976 236756 175982 236768
rect 189258 236756 189264 236768
rect 175976 236728 189264 236756
rect 175976 236716 175982 236728
rect 189258 236716 189264 236728
rect 189316 236716 189322 236768
rect 28442 236648 28448 236700
rect 28500 236688 28506 236700
rect 197446 236688 197452 236700
rect 28500 236660 197452 236688
rect 28500 236648 28506 236660
rect 197446 236648 197452 236660
rect 197504 236648 197510 236700
rect 174078 235968 174084 236020
rect 174136 236008 174142 236020
rect 174538 236008 174544 236020
rect 174136 235980 174544 236008
rect 174136 235968 174142 235980
rect 174538 235968 174544 235980
rect 174596 235968 174602 236020
rect 118602 235900 118608 235952
rect 118660 235940 118666 235952
rect 185946 235940 185952 235952
rect 118660 235912 185952 235940
rect 118660 235900 118666 235912
rect 185946 235900 185952 235912
rect 186004 235900 186010 235952
rect 195422 235900 195428 235952
rect 195480 235940 195486 235952
rect 197722 235940 197728 235952
rect 195480 235912 197728 235940
rect 195480 235900 195486 235912
rect 197722 235900 197728 235912
rect 197780 235900 197786 235952
rect 139210 235832 139216 235884
rect 139268 235872 139274 235884
rect 171962 235872 171968 235884
rect 139268 235844 171968 235872
rect 139268 235832 139274 235844
rect 171962 235832 171968 235844
rect 172020 235872 172026 235884
rect 172422 235872 172428 235884
rect 172020 235844 172428 235872
rect 172020 235832 172026 235844
rect 172422 235832 172428 235844
rect 172480 235832 172486 235884
rect 185946 235356 185952 235408
rect 186004 235396 186010 235408
rect 195422 235396 195428 235408
rect 186004 235368 195428 235396
rect 186004 235356 186010 235368
rect 195422 235356 195428 235368
rect 195480 235356 195486 235408
rect 172422 235288 172428 235340
rect 172480 235328 172486 235340
rect 188430 235328 188436 235340
rect 172480 235300 188436 235328
rect 172480 235288 172486 235300
rect 188430 235288 188436 235300
rect 188488 235288 188494 235340
rect 28902 235220 28908 235272
rect 28960 235260 28966 235272
rect 197538 235260 197544 235272
rect 28960 235232 197544 235260
rect 28960 235220 28966 235232
rect 197538 235220 197544 235232
rect 197596 235220 197602 235272
rect 108942 234540 108948 234592
rect 109000 234580 109006 234592
rect 169846 234580 169852 234592
rect 109000 234552 169852 234580
rect 109000 234540 109006 234552
rect 169846 234540 169852 234552
rect 169904 234540 169910 234592
rect 121178 234472 121184 234524
rect 121236 234512 121242 234524
rect 172698 234512 172704 234524
rect 121236 234484 172704 234512
rect 121236 234472 121242 234484
rect 172698 234472 172704 234484
rect 172756 234512 172762 234524
rect 173342 234512 173348 234524
rect 172756 234484 173348 234512
rect 172756 234472 172762 234484
rect 173342 234472 173348 234484
rect 173400 234472 173406 234524
rect 131022 234404 131028 234456
rect 131080 234444 131086 234456
rect 182082 234444 182088 234456
rect 131080 234416 182088 234444
rect 131080 234404 131086 234416
rect 182082 234404 182088 234416
rect 182140 234444 182146 234456
rect 183738 234444 183744 234456
rect 182140 234416 183744 234444
rect 182140 234404 182146 234416
rect 183738 234404 183744 234416
rect 183796 234404 183802 234456
rect 169846 233860 169852 233912
rect 169904 233900 169910 233912
rect 170582 233900 170588 233912
rect 169904 233872 170588 233900
rect 169904 233860 169910 233872
rect 170582 233860 170588 233872
rect 170640 233900 170646 233912
rect 182818 233900 182824 233912
rect 170640 233872 182824 233900
rect 170640 233860 170646 233872
rect 182818 233860 182824 233872
rect 182876 233860 182882 233912
rect 179046 233248 179052 233300
rect 179104 233288 179110 233300
rect 197354 233288 197360 233300
rect 179104 233260 197360 233288
rect 179104 233248 179110 233260
rect 197354 233248 197360 233260
rect 197412 233248 197418 233300
rect 110322 233180 110328 233232
rect 110380 233220 110386 233232
rect 171778 233220 171784 233232
rect 110380 233192 171784 233220
rect 110380 233180 110386 233192
rect 171778 233180 171784 233192
rect 171836 233220 171842 233232
rect 172422 233220 172428 233232
rect 171836 233192 172428 233220
rect 171836 233180 171842 233192
rect 172422 233180 172428 233192
rect 172480 233180 172486 233232
rect 178034 233180 178040 233232
rect 178092 233220 178098 233232
rect 178862 233220 178868 233232
rect 178092 233192 178868 233220
rect 178092 233180 178098 233192
rect 178862 233180 178868 233192
rect 178920 233180 178926 233232
rect 125502 233112 125508 233164
rect 125560 233152 125566 233164
rect 178052 233152 178080 233180
rect 125560 233124 178080 233152
rect 125560 233112 125566 233124
rect 172422 232568 172428 232620
rect 172480 232608 172486 232620
rect 181714 232608 181720 232620
rect 172480 232580 181720 232608
rect 172480 232568 172486 232580
rect 181714 232568 181720 232580
rect 181772 232568 181778 232620
rect 178954 232500 178960 232552
rect 179012 232540 179018 232552
rect 197354 232540 197360 232552
rect 179012 232512 197360 232540
rect 179012 232500 179018 232512
rect 197354 232500 197360 232512
rect 197412 232500 197418 232552
rect 565078 231820 565084 231872
rect 565136 231860 565142 231872
rect 579798 231860 579804 231872
rect 565136 231832 579804 231860
rect 565136 231820 565142 231832
rect 579798 231820 579804 231832
rect 579856 231820 579862 231872
rect 111702 231752 111708 231804
rect 111760 231792 111766 231804
rect 173066 231792 173072 231804
rect 111760 231764 173072 231792
rect 111760 231752 111766 231764
rect 173066 231752 173072 231764
rect 173124 231792 173130 231804
rect 180334 231792 180340 231804
rect 173124 231764 180340 231792
rect 173124 231752 173130 231764
rect 180334 231752 180340 231764
rect 180392 231752 180398 231804
rect 183002 231752 183008 231804
rect 183060 231792 183066 231804
rect 183186 231792 183192 231804
rect 183060 231764 183192 231792
rect 183060 231752 183066 231764
rect 183186 231752 183192 231764
rect 183244 231792 183250 231804
rect 197354 231792 197360 231804
rect 183244 231764 197360 231792
rect 183244 231752 183250 231764
rect 197354 231752 197360 231764
rect 197412 231752 197418 231804
rect 559190 231684 559196 231736
rect 559248 231724 559254 231736
rect 560938 231724 560944 231736
rect 559248 231696 560944 231724
rect 559248 231684 559254 231696
rect 560938 231684 560944 231696
rect 560996 231684 561002 231736
rect 148318 231072 148324 231124
rect 148376 231112 148382 231124
rect 171134 231112 171140 231124
rect 148376 231084 171140 231112
rect 148376 231072 148382 231084
rect 171134 231072 171140 231084
rect 171192 231112 171198 231124
rect 183002 231112 183008 231124
rect 171192 231084 183008 231112
rect 171192 231072 171198 231084
rect 183002 231072 183008 231084
rect 183060 231072 183066 231124
rect 29822 230392 29828 230444
rect 29880 230432 29886 230444
rect 47578 230432 47584 230444
rect 29880 230404 47584 230432
rect 29880 230392 29886 230404
rect 47578 230392 47584 230404
rect 47636 230392 47642 230444
rect 180150 229712 180156 229764
rect 180208 229752 180214 229764
rect 197538 229752 197544 229764
rect 180208 229724 197544 229752
rect 180208 229712 180214 229724
rect 197538 229712 197544 229724
rect 197596 229712 197602 229764
rect 28718 229576 28724 229628
rect 28776 229616 28782 229628
rect 29822 229616 29828 229628
rect 28776 229588 29828 229616
rect 28776 229576 28782 229588
rect 29822 229576 29828 229588
rect 29880 229576 29886 229628
rect 28534 229100 28540 229152
rect 28592 229140 28598 229152
rect 28592 229112 28994 229140
rect 28592 229100 28598 229112
rect 28966 229072 28994 229112
rect 29638 229072 29644 229084
rect 28966 229044 29644 229072
rect 29638 229032 29644 229044
rect 29696 229072 29702 229084
rect 46750 229072 46756 229084
rect 29696 229044 46756 229072
rect 29696 229032 29702 229044
rect 46750 229032 46756 229044
rect 46808 229072 46814 229084
rect 50338 229072 50344 229084
rect 46808 229044 50344 229072
rect 46808 229032 46814 229044
rect 50338 229032 50344 229044
rect 50396 229032 50402 229084
rect 135162 229032 135168 229084
rect 135220 229072 135226 229084
rect 168558 229072 168564 229084
rect 135220 229044 168564 229072
rect 135220 229032 135226 229044
rect 168558 229032 168564 229044
rect 168616 229032 168622 229084
rect 185026 229032 185032 229084
rect 185084 229072 185090 229084
rect 198366 229072 198372 229084
rect 185084 229044 198372 229072
rect 185084 229032 185090 229044
rect 198366 229032 198372 229044
rect 198424 229032 198430 229084
rect 136450 228964 136456 229016
rect 136508 229004 136514 229016
rect 170490 229004 170496 229016
rect 136508 228976 170496 229004
rect 136508 228964 136514 228976
rect 170490 228964 170496 228976
rect 170548 228964 170554 229016
rect 191190 228964 191196 229016
rect 191248 229004 191254 229016
rect 198918 229004 198924 229016
rect 191248 228976 198924 229004
rect 191248 228964 191254 228976
rect 198918 228964 198924 228976
rect 198976 228964 198982 229016
rect 170490 228556 170496 228608
rect 170548 228596 170554 228608
rect 177574 228596 177580 228608
rect 170548 228568 177580 228596
rect 170548 228556 170554 228568
rect 177574 228556 177580 228568
rect 177632 228556 177638 228608
rect 176102 228488 176108 228540
rect 176160 228528 176166 228540
rect 185026 228528 185032 228540
rect 176160 228500 185032 228528
rect 176160 228488 176166 228500
rect 185026 228488 185032 228500
rect 185084 228488 185090 228540
rect 174630 228420 174636 228472
rect 174688 228460 174694 228472
rect 191926 228460 191932 228472
rect 174688 228432 191932 228460
rect 174688 228420 174694 228432
rect 191926 228420 191932 228432
rect 191984 228460 191990 228472
rect 199102 228460 199108 228472
rect 191984 228432 199108 228460
rect 191984 228420 191990 228432
rect 199102 228420 199108 228432
rect 199160 228420 199166 228472
rect 3694 228352 3700 228404
rect 3752 228392 3758 228404
rect 195238 228392 195244 228404
rect 3752 228364 195244 228392
rect 3752 228352 3758 228364
rect 195238 228352 195244 228364
rect 195296 228352 195302 228404
rect 29822 227740 29828 227792
rect 29880 227780 29886 227792
rect 34514 227780 34520 227792
rect 29880 227752 34520 227780
rect 29880 227740 29886 227752
rect 34514 227740 34520 227752
rect 34572 227780 34578 227792
rect 35158 227780 35164 227792
rect 34572 227752 35164 227780
rect 34572 227740 34578 227752
rect 35158 227740 35164 227752
rect 35216 227740 35222 227792
rect 168558 227740 168564 227792
rect 168616 227780 168622 227792
rect 187142 227780 187148 227792
rect 168616 227752 187148 227780
rect 168616 227740 168622 227752
rect 187142 227740 187148 227752
rect 187200 227740 187206 227792
rect 133782 227672 133788 227724
rect 133840 227712 133846 227724
rect 187050 227712 187056 227724
rect 133840 227684 187056 227712
rect 133840 227672 133846 227684
rect 187050 227672 187056 227684
rect 187108 227672 187114 227724
rect 192478 227672 192484 227724
rect 192536 227712 192542 227724
rect 198550 227712 198556 227724
rect 192536 227684 198556 227712
rect 192536 227672 192542 227684
rect 198550 227672 198556 227684
rect 198608 227672 198614 227724
rect 137922 227604 137928 227656
rect 137980 227644 137986 227656
rect 171870 227644 171876 227656
rect 137980 227616 171876 227644
rect 137980 227604 137986 227616
rect 171870 227604 171876 227616
rect 171928 227644 171934 227656
rect 172422 227644 172428 227656
rect 171928 227616 172428 227644
rect 171928 227604 171934 227616
rect 172422 227604 172428 227616
rect 172480 227604 172486 227656
rect 136358 227536 136364 227588
rect 136416 227576 136422 227588
rect 170214 227576 170220 227588
rect 136416 227548 170220 227576
rect 136416 227536 136422 227548
rect 170214 227536 170220 227548
rect 170272 227536 170278 227588
rect 170214 227128 170220 227180
rect 170272 227168 170278 227180
rect 180886 227168 180892 227180
rect 170272 227140 180892 227168
rect 170272 227128 170278 227140
rect 180886 227128 180892 227140
rect 180944 227128 180950 227180
rect 172422 227060 172428 227112
rect 172480 227100 172486 227112
rect 193950 227100 193956 227112
rect 172480 227072 193956 227100
rect 172480 227060 172486 227072
rect 193950 227060 193956 227072
rect 194008 227060 194014 227112
rect 3878 226992 3884 227044
rect 3936 227032 3942 227044
rect 172146 227032 172152 227044
rect 3936 227004 172152 227032
rect 3936 226992 3942 227004
rect 172146 226992 172152 227004
rect 172204 226992 172210 227044
rect 187050 226312 187056 226364
rect 187108 226352 187114 226364
rect 189350 226352 189356 226364
rect 187108 226324 189356 226352
rect 187108 226312 187114 226324
rect 189350 226312 189356 226324
rect 189408 226312 189414 226364
rect 183554 226244 183560 226296
rect 183612 226284 183618 226296
rect 198458 226284 198464 226296
rect 183612 226256 198464 226284
rect 183612 226244 183618 226256
rect 198458 226244 198464 226256
rect 198516 226244 198522 226296
rect 171778 225564 171784 225616
rect 171836 225604 171842 225616
rect 183554 225604 183560 225616
rect 171836 225576 183560 225604
rect 171836 225564 171842 225576
rect 183554 225564 183560 225576
rect 183612 225564 183618 225616
rect 181622 224204 181628 224256
rect 181680 224244 181686 224256
rect 185026 224244 185032 224256
rect 181680 224216 185032 224244
rect 181680 224204 181686 224216
rect 185026 224204 185032 224216
rect 185084 224244 185090 224256
rect 197354 224244 197360 224256
rect 185084 224216 197360 224244
rect 185084 224204 185090 224216
rect 197354 224204 197360 224216
rect 197412 224204 197418 224256
rect 187878 223524 187884 223576
rect 187936 223564 187942 223576
rect 199010 223564 199016 223576
rect 187936 223536 199016 223564
rect 187936 223524 187942 223536
rect 199010 223524 199016 223536
rect 199068 223564 199074 223576
rect 199562 223564 199568 223576
rect 199068 223536 199568 223564
rect 199068 223524 199074 223536
rect 199562 223524 199568 223536
rect 199620 223524 199626 223576
rect 560202 223524 560208 223576
rect 560260 223564 560266 223576
rect 567838 223564 567844 223576
rect 560260 223536 567844 223564
rect 560260 223524 560266 223536
rect 567838 223524 567844 223536
rect 567896 223524 567902 223576
rect 171870 222844 171876 222896
rect 171928 222884 171934 222896
rect 187878 222884 187884 222896
rect 171928 222856 187884 222884
rect 171928 222844 171934 222856
rect 187878 222844 187884 222856
rect 187936 222844 187942 222896
rect 193490 220804 193496 220856
rect 193548 220844 193554 220856
rect 198918 220844 198924 220856
rect 193548 220816 198924 220844
rect 193548 220804 193554 220816
rect 198918 220804 198924 220816
rect 198976 220804 198982 220856
rect 184382 220056 184388 220108
rect 184440 220096 184446 220108
rect 197354 220096 197360 220108
rect 184440 220068 197360 220096
rect 184440 220056 184446 220068
rect 197354 220056 197360 220068
rect 197412 220056 197418 220108
rect 195330 218764 195336 218816
rect 195388 218804 195394 218816
rect 197906 218804 197912 218816
rect 195388 218776 197912 218804
rect 195388 218764 195394 218776
rect 197906 218764 197912 218776
rect 197964 218764 197970 218816
rect 174814 218696 174820 218748
rect 174872 218736 174878 218748
rect 193490 218736 193496 218748
rect 174872 218708 193496 218736
rect 174872 218696 174878 218708
rect 193490 218696 193496 218708
rect 193548 218696 193554 218748
rect 559558 218016 559564 218068
rect 559616 218056 559622 218068
rect 579890 218056 579896 218068
rect 559616 218028 579896 218056
rect 559616 218016 559622 218028
rect 579890 218016 579896 218028
rect 579948 218016 579954 218068
rect 189166 217948 189172 218000
rect 189224 217988 189230 218000
rect 197354 217988 197360 218000
rect 189224 217960 197360 217988
rect 189224 217948 189230 217960
rect 197354 217948 197360 217960
rect 197412 217948 197418 218000
rect 171042 217268 171048 217320
rect 171100 217308 171106 217320
rect 189166 217308 189172 217320
rect 171100 217280 189172 217308
rect 171100 217268 171106 217280
rect 189166 217268 189172 217280
rect 189224 217268 189230 217320
rect 170950 215908 170956 215960
rect 171008 215948 171014 215960
rect 197354 215948 197360 215960
rect 171008 215920 197360 215948
rect 171008 215908 171014 215920
rect 197354 215908 197360 215920
rect 197412 215948 197418 215960
rect 197998 215948 198004 215960
rect 197412 215920 198004 215948
rect 197412 215908 197418 215920
rect 197998 215908 198004 215920
rect 198056 215908 198062 215960
rect 559190 215772 559196 215824
rect 559248 215812 559254 215824
rect 566458 215812 566464 215824
rect 559248 215784 566464 215812
rect 559248 215772 559254 215784
rect 566458 215772 566464 215784
rect 566516 215772 566522 215824
rect 196802 215364 196808 215416
rect 196860 215404 196866 215416
rect 197722 215404 197728 215416
rect 196860 215376 197728 215404
rect 196860 215364 196866 215376
rect 197722 215364 197728 215376
rect 197780 215404 197786 215416
rect 198090 215404 198096 215416
rect 197780 215376 198096 215404
rect 197780 215364 197786 215376
rect 198090 215364 198096 215376
rect 198148 215364 198154 215416
rect 176194 213936 176200 213988
rect 176252 213976 176258 213988
rect 179414 213976 179420 213988
rect 176252 213948 179420 213976
rect 176252 213936 176258 213948
rect 179414 213936 179420 213948
rect 179472 213976 179478 213988
rect 197354 213976 197360 213988
rect 179472 213948 197360 213976
rect 179472 213936 179478 213948
rect 197354 213936 197360 213948
rect 197412 213936 197418 213988
rect 170766 213188 170772 213240
rect 170824 213228 170830 213240
rect 178126 213228 178132 213240
rect 170824 213200 178132 213228
rect 170824 213188 170830 213200
rect 178126 213188 178132 213200
rect 178184 213188 178190 213240
rect 178126 212508 178132 212560
rect 178184 212548 178190 212560
rect 197354 212548 197360 212560
rect 178184 212520 197360 212548
rect 178184 212508 178190 212520
rect 197354 212508 197360 212520
rect 197412 212508 197418 212560
rect 186314 212440 186320 212492
rect 186372 212480 186378 212492
rect 197630 212480 197636 212492
rect 186372 212452 197636 212480
rect 186372 212440 186378 212452
rect 197630 212440 197636 212452
rect 197688 212440 197694 212492
rect 167914 211760 167920 211812
rect 167972 211800 167978 211812
rect 186314 211800 186320 211812
rect 167972 211772 186320 211800
rect 167972 211760 167978 211772
rect 186314 211760 186320 211772
rect 186372 211760 186378 211812
rect 197630 211556 197636 211608
rect 197688 211596 197694 211608
rect 197906 211596 197912 211608
rect 197688 211568 197912 211596
rect 197688 211556 197694 211568
rect 197906 211556 197912 211568
rect 197964 211556 197970 211608
rect 176654 211080 176660 211132
rect 176712 211120 176718 211132
rect 197354 211120 197360 211132
rect 176712 211092 197360 211120
rect 176712 211080 176718 211092
rect 197354 211080 197360 211092
rect 197412 211080 197418 211132
rect 170766 210400 170772 210452
rect 170824 210440 170830 210452
rect 176654 210440 176660 210452
rect 170824 210412 176660 210440
rect 170824 210400 170830 210412
rect 176654 210400 176660 210412
rect 176712 210400 176718 210452
rect 197354 210196 197360 210248
rect 197412 210236 197418 210248
rect 197722 210236 197728 210248
rect 197412 210208 197728 210236
rect 197412 210196 197418 210208
rect 197722 210196 197728 210208
rect 197780 210196 197786 210248
rect 197722 210060 197728 210112
rect 197780 210100 197786 210112
rect 197998 210100 198004 210112
rect 197780 210072 198004 210100
rect 197780 210060 197786 210072
rect 197998 210060 198004 210072
rect 198056 210060 198062 210112
rect 182910 209176 182916 209228
rect 182968 209216 182974 209228
rect 197354 209216 197360 209228
rect 182968 209188 197360 209216
rect 182968 209176 182974 209188
rect 197354 209176 197360 209188
rect 197412 209176 197418 209228
rect 197722 209176 197728 209228
rect 197780 209216 197786 209228
rect 197906 209216 197912 209228
rect 197780 209188 197912 209216
rect 197780 209176 197786 209188
rect 197906 209176 197912 209188
rect 197964 209176 197970 209228
rect 178770 209040 178776 209092
rect 178828 209080 178834 209092
rect 180978 209080 180984 209092
rect 178828 209052 180984 209080
rect 178828 209040 178834 209052
rect 180978 209040 180984 209052
rect 181036 209040 181042 209092
rect 176194 208292 176200 208344
rect 176252 208332 176258 208344
rect 182174 208332 182180 208344
rect 176252 208304 182180 208332
rect 176252 208292 176258 208304
rect 182174 208292 182180 208304
rect 182232 208332 182238 208344
rect 197354 208332 197360 208344
rect 182232 208304 197360 208332
rect 182232 208292 182238 208304
rect 197354 208292 197360 208304
rect 197412 208292 197418 208344
rect 560202 208292 560208 208344
rect 560260 208332 560266 208344
rect 580258 208332 580264 208344
rect 560260 208304 580264 208332
rect 560260 208292 560266 208304
rect 580258 208292 580264 208304
rect 580316 208292 580322 208344
rect 180058 206320 180064 206372
rect 180116 206360 180122 206372
rect 196066 206360 196072 206372
rect 180116 206332 196072 206360
rect 180116 206320 180122 206332
rect 196066 206320 196072 206332
rect 196124 206360 196130 206372
rect 197354 206360 197360 206372
rect 196124 206332 197360 206360
rect 196124 206320 196130 206332
rect 197354 206320 197360 206332
rect 197412 206320 197418 206372
rect 170950 206252 170956 206304
rect 171008 206292 171014 206304
rect 180978 206292 180984 206304
rect 171008 206264 180984 206292
rect 171008 206252 171014 206264
rect 180978 206252 180984 206264
rect 181036 206292 181042 206304
rect 197722 206292 197728 206304
rect 181036 206264 197728 206292
rect 181036 206252 181042 206264
rect 197722 206252 197728 206264
rect 197780 206252 197786 206304
rect 170858 204892 170864 204944
rect 170916 204932 170922 204944
rect 186314 204932 186320 204944
rect 170916 204904 186320 204932
rect 170916 204892 170922 204904
rect 186314 204892 186320 204904
rect 186372 204892 186378 204944
rect 186314 204280 186320 204332
rect 186372 204320 186378 204332
rect 186498 204320 186504 204332
rect 186372 204292 186504 204320
rect 186372 204280 186378 204292
rect 186498 204280 186504 204292
rect 186556 204320 186562 204332
rect 197354 204320 197360 204332
rect 186556 204292 197360 204320
rect 186556 204280 186562 204292
rect 197354 204280 197360 204292
rect 197412 204280 197418 204332
rect 168098 204212 168104 204264
rect 168156 204252 168162 204264
rect 169754 204252 169760 204264
rect 168156 204224 169760 204252
rect 168156 204212 168162 204224
rect 169754 204212 169760 204224
rect 169812 204252 169818 204264
rect 197722 204252 197728 204264
rect 169812 204224 197728 204252
rect 169812 204212 169818 204224
rect 197722 204212 197728 204224
rect 197780 204212 197786 204264
rect 184934 204144 184940 204196
rect 184992 204184 184998 204196
rect 185394 204184 185400 204196
rect 184992 204156 185400 204184
rect 184992 204144 184998 204156
rect 185394 204144 185400 204156
rect 185452 204184 185458 204196
rect 197354 204184 197360 204196
rect 185452 204156 197360 204184
rect 185452 204144 185458 204156
rect 197354 204144 197360 204156
rect 197412 204144 197418 204196
rect 168006 203532 168012 203584
rect 168064 203572 168070 203584
rect 185394 203572 185400 203584
rect 168064 203544 185400 203572
rect 168064 203532 168070 203544
rect 185394 203532 185400 203544
rect 185452 203532 185458 203584
rect 181530 202784 181536 202836
rect 181588 202824 181594 202836
rect 187878 202824 187884 202836
rect 181588 202796 187884 202824
rect 181588 202784 181594 202796
rect 187878 202784 187884 202796
rect 187936 202784 187942 202836
rect 191282 202784 191288 202836
rect 191340 202824 191346 202836
rect 197906 202824 197912 202836
rect 191340 202796 197912 202824
rect 191340 202784 191346 202796
rect 197906 202784 197912 202796
rect 197964 202784 197970 202836
rect 187878 201492 187884 201544
rect 187936 201532 187942 201544
rect 197354 201532 197360 201544
rect 187936 201504 197360 201532
rect 187936 201492 187942 201504
rect 197354 201492 197360 201504
rect 197412 201492 197418 201544
rect 168190 200744 168196 200796
rect 168248 200784 168254 200796
rect 191834 200784 191840 200796
rect 168248 200756 191840 200784
rect 168248 200744 168254 200756
rect 191834 200744 191840 200756
rect 191892 200784 191898 200796
rect 197354 200784 197360 200796
rect 191892 200756 197360 200784
rect 191892 200744 191898 200756
rect 197354 200744 197360 200756
rect 197412 200744 197418 200796
rect 184290 199384 184296 199436
rect 184348 199424 184354 199436
rect 193306 199424 193312 199436
rect 184348 199396 193312 199424
rect 184348 199384 184354 199396
rect 193306 199384 193312 199396
rect 193364 199424 193370 199436
rect 197354 199424 197360 199436
rect 193364 199396 197360 199424
rect 193364 199384 193370 199396
rect 197354 199384 197360 199396
rect 197412 199384 197418 199436
rect 168282 197956 168288 198008
rect 168340 197996 168346 198008
rect 190454 197996 190460 198008
rect 168340 197968 190460 197996
rect 168340 197956 168346 197968
rect 190454 197956 190460 197968
rect 190512 197996 190518 198008
rect 197354 197996 197360 198008
rect 190512 197968 197360 197996
rect 190512 197956 190518 197968
rect 197354 197956 197360 197968
rect 197412 197956 197418 198008
rect 189074 197276 189080 197328
rect 189132 197316 189138 197328
rect 197354 197316 197360 197328
rect 189132 197288 197360 197316
rect 189132 197276 189138 197288
rect 197354 197276 197360 197288
rect 197412 197276 197418 197328
rect 173434 196596 173440 196648
rect 173492 196636 173498 196648
rect 189074 196636 189080 196648
rect 173492 196608 189080 196636
rect 173492 196596 173498 196608
rect 189074 196596 189080 196608
rect 189132 196596 189138 196648
rect 194594 195916 194600 195968
rect 194652 195956 194658 195968
rect 197354 195956 197360 195968
rect 194652 195928 197360 195956
rect 194652 195916 194658 195928
rect 197354 195916 197360 195928
rect 197412 195916 197418 195968
rect 181622 195236 181628 195288
rect 181680 195276 181686 195288
rect 194594 195276 194600 195288
rect 181680 195248 194600 195276
rect 181680 195236 181686 195248
rect 194594 195236 194600 195248
rect 194652 195236 194658 195288
rect 187786 194488 187792 194540
rect 187844 194528 187850 194540
rect 197354 194528 197360 194540
rect 187844 194500 197360 194528
rect 187844 194488 187850 194500
rect 197354 194488 197360 194500
rect 197412 194488 197418 194540
rect 174906 193808 174912 193860
rect 174964 193848 174970 193860
rect 187786 193848 187792 193860
rect 174964 193820 187792 193848
rect 174964 193808 174970 193820
rect 187786 193808 187792 193820
rect 187844 193808 187850 193860
rect 177758 192448 177764 192500
rect 177816 192488 177822 192500
rect 193214 192488 193220 192500
rect 177816 192460 193220 192488
rect 177816 192448 177822 192460
rect 193214 192448 193220 192460
rect 193272 192488 193278 192500
rect 197722 192488 197728 192500
rect 193272 192460 197728 192488
rect 193272 192448 193278 192460
rect 197722 192448 197728 192460
rect 197780 192448 197786 192500
rect 186958 191836 186964 191888
rect 187016 191876 187022 191888
rect 190454 191876 190460 191888
rect 187016 191848 190460 191876
rect 187016 191836 187022 191848
rect 190454 191836 190460 191848
rect 190512 191876 190518 191888
rect 197354 191876 197360 191888
rect 190512 191848 197360 191876
rect 190512 191836 190518 191848
rect 197354 191836 197360 191848
rect 197412 191836 197418 191888
rect 560938 191836 560944 191888
rect 560996 191876 561002 191888
rect 580166 191876 580172 191888
rect 560996 191848 580172 191876
rect 560996 191836 561002 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 560202 191700 560208 191752
rect 560260 191740 560266 191752
rect 565078 191740 565084 191752
rect 560260 191712 565084 191740
rect 560260 191700 560266 191712
rect 565078 191700 565084 191712
rect 565136 191700 565142 191752
rect 185578 191088 185584 191140
rect 185636 191128 185642 191140
rect 197354 191128 197360 191140
rect 185636 191100 197360 191128
rect 185636 191088 185642 191100
rect 197354 191088 197360 191100
rect 197412 191088 197418 191140
rect 182818 189728 182824 189780
rect 182876 189768 182882 189780
rect 197354 189768 197360 189780
rect 182876 189740 197360 189768
rect 182876 189728 182882 189740
rect 197354 189728 197360 189740
rect 197412 189728 197418 189780
rect 181714 188300 181720 188352
rect 181772 188340 181778 188352
rect 197354 188340 197360 188352
rect 181772 188312 197360 188340
rect 181772 188300 181778 188312
rect 197354 188300 197360 188312
rect 197412 188300 197418 188352
rect 181530 187688 181536 187740
rect 181588 187728 181594 187740
rect 181714 187728 181720 187740
rect 181588 187700 181720 187728
rect 181588 187688 181594 187700
rect 181714 187688 181720 187700
rect 181772 187688 181778 187740
rect 180058 186940 180064 186992
rect 180116 186980 180122 186992
rect 180334 186980 180340 186992
rect 180116 186952 180340 186980
rect 180116 186940 180122 186952
rect 180334 186940 180340 186952
rect 180392 186980 180398 186992
rect 197354 186980 197360 186992
rect 180392 186952 197360 186980
rect 180392 186940 180398 186952
rect 197354 186940 197360 186952
rect 197412 186940 197418 186992
rect 178678 185580 178684 185632
rect 178736 185620 178742 185632
rect 179138 185620 179144 185632
rect 178736 185592 179144 185620
rect 178736 185580 178742 185592
rect 179138 185580 179144 185592
rect 179196 185620 179202 185632
rect 197354 185620 197360 185632
rect 179196 185592 197360 185620
rect 179196 185580 179202 185592
rect 197354 185580 197360 185592
rect 197412 185580 197418 185632
rect 560018 184832 560024 184884
rect 560076 184872 560082 184884
rect 580258 184872 580264 184884
rect 560076 184844 580264 184872
rect 560076 184832 560082 184844
rect 580258 184832 580264 184844
rect 580316 184832 580322 184884
rect 177298 184152 177304 184204
rect 177356 184192 177362 184204
rect 197354 184192 197360 184204
rect 177356 184164 197360 184192
rect 177356 184152 177362 184164
rect 197354 184152 197360 184164
rect 197412 184152 197418 184204
rect 170490 182792 170496 182844
rect 170548 182832 170554 182844
rect 192018 182832 192024 182844
rect 170548 182804 192024 182832
rect 170548 182792 170554 182804
rect 192018 182792 192024 182804
rect 192076 182832 192082 182844
rect 197354 182832 197360 182844
rect 192076 182804 197360 182832
rect 192076 182792 192082 182804
rect 197354 182792 197360 182804
rect 197412 182792 197418 182844
rect 175274 182112 175280 182164
rect 175332 182152 175338 182164
rect 175734 182152 175740 182164
rect 175332 182124 175740 182152
rect 175332 182112 175338 182124
rect 175734 182112 175740 182124
rect 175792 182152 175798 182164
rect 197354 182152 197360 182164
rect 175792 182124 197360 182152
rect 175792 182112 175798 182124
rect 197354 182112 197360 182124
rect 197412 182112 197418 182164
rect 170398 181432 170404 181484
rect 170456 181472 170462 181484
rect 175734 181472 175740 181484
rect 170456 181444 175740 181472
rect 170456 181432 170462 181444
rect 175734 181432 175740 181444
rect 175792 181432 175798 181484
rect 174538 180072 174544 180124
rect 174596 180112 174602 180124
rect 197354 180112 197360 180124
rect 174596 180084 197360 180112
rect 174596 180072 174602 180084
rect 197354 180072 197360 180084
rect 197412 180072 197418 180124
rect 195238 179460 195244 179512
rect 195296 179500 195302 179512
rect 197354 179500 197360 179512
rect 195296 179472 197360 179500
rect 195296 179460 195302 179472
rect 197354 179460 197360 179472
rect 197412 179460 197418 179512
rect 168926 178644 168932 178696
rect 168984 178684 168990 178696
rect 181714 178684 181720 178696
rect 168984 178656 181720 178684
rect 168984 178644 168990 178656
rect 181714 178644 181720 178656
rect 181772 178644 181778 178696
rect 196802 178236 196808 178288
rect 196860 178276 196866 178288
rect 197906 178276 197912 178288
rect 196860 178248 197912 178276
rect 196860 178236 196866 178248
rect 197906 178236 197912 178248
rect 197964 178236 197970 178288
rect 169294 177352 169300 177404
rect 169352 177392 169358 177404
rect 180334 177392 180340 177404
rect 169352 177364 180340 177392
rect 169352 177352 169358 177364
rect 180334 177352 180340 177364
rect 180392 177352 180398 177404
rect 173342 177284 173348 177336
rect 173400 177324 173406 177336
rect 197354 177324 197360 177336
rect 173400 177296 197360 177324
rect 173400 177284 173406 177296
rect 197354 177284 197360 177296
rect 197412 177284 197418 177336
rect 560202 176604 560208 176656
rect 560260 176644 560266 176656
rect 580166 176644 580172 176656
rect 560260 176616 580172 176644
rect 560260 176604 560266 176616
rect 580166 176604 580172 176616
rect 580224 176604 580230 176656
rect 168926 175992 168932 176044
rect 168984 176032 168990 176044
rect 178218 176032 178224 176044
rect 168984 176004 178224 176032
rect 168984 175992 168990 176004
rect 178218 175992 178224 176004
rect 178276 175992 178282 176044
rect 169202 175924 169208 175976
rect 169260 175964 169266 175976
rect 197630 175964 197636 175976
rect 169260 175936 197636 175964
rect 169260 175924 169266 175936
rect 197630 175924 197636 175936
rect 197688 175924 197694 175976
rect 191098 175652 191104 175704
rect 191156 175692 191162 175704
rect 197354 175692 197360 175704
rect 191156 175664 197360 175692
rect 191156 175652 191162 175664
rect 197354 175652 197360 175664
rect 197412 175652 197418 175704
rect 182082 175176 182088 175228
rect 182140 175216 182146 175228
rect 197354 175216 197360 175228
rect 182140 175188 197360 175216
rect 182140 175176 182146 175188
rect 197354 175176 197360 175188
rect 197412 175176 197418 175228
rect 168834 174564 168840 174616
rect 168892 174604 168898 174616
rect 174998 174604 175004 174616
rect 168892 174576 175004 174604
rect 168892 174564 168898 174576
rect 174998 174564 175004 174576
rect 175056 174564 175062 174616
rect 170674 174496 170680 174548
rect 170732 174536 170738 174548
rect 180794 174536 180800 174548
rect 170732 174508 180800 174536
rect 170732 174496 170738 174508
rect 180794 174496 180800 174508
rect 180852 174536 180858 174548
rect 182082 174536 182088 174548
rect 180852 174508 182088 174536
rect 180852 174496 180858 174508
rect 182082 174496 182088 174508
rect 182140 174496 182146 174548
rect 180242 173204 180248 173256
rect 180300 173244 180306 173256
rect 197354 173244 197360 173256
rect 180300 173216 197360 173244
rect 180300 173204 180306 173216
rect 197354 173204 197360 173216
rect 197412 173204 197418 173256
rect 168742 173136 168748 173188
rect 168800 173176 168806 173188
rect 194594 173176 194600 173188
rect 168800 173148 194600 173176
rect 168800 173136 168806 173148
rect 194594 173136 194600 173148
rect 194652 173136 194658 173188
rect 174630 172456 174636 172508
rect 174688 172496 174694 172508
rect 178034 172496 178040 172508
rect 174688 172468 178040 172496
rect 174688 172456 174694 172468
rect 178034 172456 178040 172468
rect 178092 172496 178098 172508
rect 197354 172496 197360 172508
rect 178092 172468 197360 172496
rect 178092 172456 178098 172468
rect 197354 172456 197360 172468
rect 197412 172456 197418 172508
rect 168926 171776 168932 171828
rect 168984 171816 168990 171828
rect 177850 171816 177856 171828
rect 168984 171788 177856 171816
rect 168984 171776 168990 171788
rect 177850 171776 177856 171788
rect 177908 171776 177914 171828
rect 169110 170484 169116 170536
rect 169168 170524 169174 170536
rect 178954 170524 178960 170536
rect 169168 170496 178960 170524
rect 169168 170484 169174 170496
rect 178954 170484 178960 170496
rect 179012 170484 179018 170536
rect 177390 170416 177396 170468
rect 177448 170456 177454 170468
rect 197354 170456 197360 170468
rect 177448 170428 197360 170456
rect 177448 170416 177454 170428
rect 197354 170416 197360 170428
rect 197412 170416 197418 170468
rect 169018 170348 169024 170400
rect 169076 170388 169082 170400
rect 197538 170388 197544 170400
rect 169076 170360 197544 170388
rect 169076 170348 169082 170360
rect 197538 170348 197544 170360
rect 197596 170348 197602 170400
rect 187694 169668 187700 169720
rect 187752 169708 187758 169720
rect 197354 169708 197360 169720
rect 187752 169680 197360 169708
rect 187752 169668 187758 169680
rect 197354 169668 197360 169680
rect 197412 169668 197418 169720
rect 178770 168988 178776 169040
rect 178828 169028 178834 169040
rect 187694 169028 187700 169040
rect 178828 169000 187700 169028
rect 178828 168988 178834 169000
rect 187694 168988 187700 169000
rect 187752 168988 187758 169040
rect 194686 168308 194692 168360
rect 194744 168348 194750 168360
rect 197538 168348 197544 168360
rect 194744 168320 197544 168348
rect 194744 168308 194750 168320
rect 197538 168308 197544 168320
rect 197596 168308 197602 168360
rect 559006 168240 559012 168292
rect 559064 168280 559070 168292
rect 560938 168280 560944 168292
rect 559064 168252 560944 168280
rect 559064 168240 559070 168252
rect 560938 168240 560944 168252
rect 560996 168240 561002 168292
rect 184290 167696 184296 167748
rect 184348 167736 184354 167748
rect 194686 167736 194692 167748
rect 184348 167708 194692 167736
rect 184348 167696 184354 167708
rect 194686 167696 194692 167708
rect 194744 167696 194750 167748
rect 174722 167628 174728 167680
rect 174780 167668 174786 167680
rect 197354 167668 197360 167680
rect 174780 167640 197360 167668
rect 174780 167628 174786 167640
rect 197354 167628 197360 167640
rect 197412 167628 197418 167680
rect 184842 166948 184848 167000
rect 184900 166988 184906 167000
rect 197354 166988 197360 167000
rect 184900 166960 197360 166988
rect 184900 166948 184906 166960
rect 197354 166948 197360 166960
rect 197412 166948 197418 167000
rect 177482 166268 177488 166320
rect 177540 166308 177546 166320
rect 183738 166308 183744 166320
rect 177540 166280 183744 166308
rect 177540 166268 177546 166280
rect 183738 166268 183744 166280
rect 183796 166308 183802 166320
rect 184842 166308 184848 166320
rect 183796 166280 184848 166308
rect 183796 166268 183802 166280
rect 184842 166268 184848 166280
rect 184900 166268 184906 166320
rect 559558 165588 559564 165640
rect 559616 165628 559622 165640
rect 580166 165628 580172 165640
rect 559616 165600 580172 165628
rect 559616 165588 559622 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 178862 164908 178868 164960
rect 178920 164948 178926 164960
rect 193398 164948 193404 164960
rect 178920 164920 193404 164948
rect 178920 164908 178926 164920
rect 193398 164908 193404 164920
rect 193456 164948 193462 164960
rect 197354 164948 197360 164960
rect 193456 164920 197360 164948
rect 193456 164908 193462 164920
rect 197354 164908 197360 164920
rect 197412 164908 197418 164960
rect 169110 164840 169116 164892
rect 169168 164880 169174 164892
rect 195974 164880 195980 164892
rect 169168 164852 195980 164880
rect 169168 164840 169174 164852
rect 195974 164840 195980 164852
rect 196032 164840 196038 164892
rect 188338 164160 188344 164212
rect 188396 164200 188402 164212
rect 189350 164200 189356 164212
rect 188396 164172 189356 164200
rect 188396 164160 188402 164172
rect 189350 164160 189356 164172
rect 189408 164200 189414 164212
rect 197354 164200 197360 164212
rect 189408 164172 197360 164200
rect 189408 164160 189414 164172
rect 197354 164160 197360 164172
rect 197412 164160 197418 164212
rect 187142 162120 187148 162172
rect 187200 162160 187206 162172
rect 197354 162160 197360 162172
rect 187200 162132 197360 162160
rect 187200 162120 187206 162132
rect 197354 162120 197360 162132
rect 197412 162120 197418 162172
rect 180794 161372 180800 161424
rect 180852 161412 180858 161424
rect 197354 161412 197360 161424
rect 180852 161384 197360 161412
rect 180852 161372 180858 161384
rect 197354 161372 197360 161384
rect 197412 161372 197418 161424
rect 170582 160692 170588 160744
rect 170640 160732 170646 160744
rect 180794 160732 180800 160744
rect 170640 160704 180800 160732
rect 170640 160692 170646 160704
rect 180794 160692 180800 160704
rect 180852 160692 180858 160744
rect 177574 159332 177580 159384
rect 177632 159372 177638 159384
rect 197354 159372 197360 159384
rect 177632 159344 197360 159372
rect 177632 159332 177638 159344
rect 197354 159332 197360 159344
rect 197412 159332 197418 159384
rect 193950 158312 193956 158364
rect 194008 158352 194014 158364
rect 197354 158352 197360 158364
rect 194008 158324 197360 158352
rect 194008 158312 194014 158324
rect 197354 158312 197360 158324
rect 197412 158312 197418 158364
rect 188430 156612 188436 156664
rect 188488 156652 188494 156664
rect 197354 156652 197360 156664
rect 188488 156624 197360 156652
rect 188488 156612 188494 156624
rect 197354 156612 197360 156624
rect 197412 156612 197418 156664
rect 189074 155864 189080 155916
rect 189132 155904 189138 155916
rect 189258 155904 189264 155916
rect 189132 155876 189264 155904
rect 189132 155864 189138 155876
rect 189258 155864 189264 155876
rect 189316 155904 189322 155916
rect 197538 155904 197544 155916
rect 189316 155876 197544 155904
rect 189316 155864 189322 155876
rect 197538 155864 197544 155876
rect 197596 155864 197602 155916
rect 167730 155252 167736 155304
rect 167788 155292 167794 155304
rect 189074 155292 189080 155304
rect 167788 155264 189080 155292
rect 167788 155252 167794 155264
rect 189074 155252 189080 155264
rect 189132 155252 189138 155304
rect 167638 155184 167644 155236
rect 167696 155224 167702 155236
rect 197354 155224 197360 155236
rect 167696 155196 197360 155224
rect 167696 155184 167702 155196
rect 197354 155184 197360 155196
rect 197412 155184 197418 155236
rect 184842 154504 184848 154556
rect 184900 154544 184906 154556
rect 197354 154544 197360 154556
rect 184900 154516 197360 154544
rect 184900 154504 184906 154516
rect 197354 154504 197360 154516
rect 197412 154504 197418 154556
rect 175918 153824 175924 153876
rect 175976 153864 175982 153876
rect 183646 153864 183652 153876
rect 175976 153836 183652 153864
rect 175976 153824 175982 153836
rect 183646 153824 183652 153836
rect 183704 153864 183710 153876
rect 184842 153864 184848 153876
rect 183704 153836 184848 153864
rect 183704 153824 183710 153836
rect 184842 153824 184848 153836
rect 184900 153824 184906 153876
rect 186314 153144 186320 153196
rect 186372 153184 186378 153196
rect 197354 153184 197360 153196
rect 186372 153156 197360 153184
rect 186372 153144 186378 153156
rect 197354 153144 197360 153156
rect 197412 153144 197418 153196
rect 176010 152464 176016 152516
rect 176068 152504 176074 152516
rect 186314 152504 186320 152516
rect 176068 152476 186320 152504
rect 176068 152464 176074 152476
rect 186314 152464 186320 152476
rect 186372 152464 186378 152516
rect 168742 151036 168748 151088
rect 168800 151076 168806 151088
rect 179046 151076 179052 151088
rect 168800 151048 179052 151076
rect 168800 151036 168806 151048
rect 179046 151036 179052 151048
rect 179104 151036 179110 151088
rect 197354 150464 197360 150476
rect 173544 150436 197360 150464
rect 168558 150356 168564 150408
rect 168616 150396 168622 150408
rect 173544 150396 173572 150436
rect 197354 150424 197360 150436
rect 197412 150424 197418 150476
rect 168616 150368 173572 150396
rect 168616 150356 168622 150368
rect 181714 149064 181720 149116
rect 181772 149104 181778 149116
rect 187694 149104 187700 149116
rect 181772 149076 187700 149104
rect 181772 149064 181778 149076
rect 187694 149064 187700 149076
rect 187752 149104 187758 149116
rect 197354 149104 197360 149116
rect 187752 149076 197360 149104
rect 187752 149064 187758 149076
rect 197354 149064 197360 149076
rect 197412 149064 197418 149116
rect 180334 148996 180340 149048
rect 180392 149036 180398 149048
rect 181898 149036 181904 149048
rect 180392 149008 181904 149036
rect 180392 148996 180398 149008
rect 181898 148996 181904 149008
rect 181956 148996 181962 149048
rect 180794 147636 180800 147688
rect 180852 147676 180858 147688
rect 181898 147676 181904 147688
rect 180852 147648 181904 147676
rect 180852 147636 180858 147648
rect 181898 147636 181904 147648
rect 181956 147676 181962 147688
rect 197538 147676 197544 147688
rect 181956 147648 197544 147676
rect 181956 147636 181962 147648
rect 197538 147636 197544 147648
rect 197596 147636 197602 147688
rect 177666 147568 177672 147620
rect 177724 147608 177730 147620
rect 178218 147608 178224 147620
rect 177724 147580 178224 147608
rect 177724 147568 177730 147580
rect 178218 147568 178224 147580
rect 178276 147608 178282 147620
rect 197354 147608 197360 147620
rect 178276 147580 197360 147608
rect 178276 147568 178282 147580
rect 197354 147568 197360 147580
rect 197412 147568 197418 147620
rect 174998 146208 175004 146260
rect 175056 146248 175062 146260
rect 178034 146248 178040 146260
rect 175056 146220 178040 146248
rect 175056 146208 175062 146220
rect 178034 146208 178040 146220
rect 178092 146208 178098 146260
rect 178034 144916 178040 144968
rect 178092 144956 178098 144968
rect 197354 144956 197360 144968
rect 178092 144928 197360 144956
rect 178092 144916 178098 144928
rect 197354 144916 197360 144928
rect 197412 144916 197418 144968
rect 560018 144848 560024 144900
rect 560076 144888 560082 144900
rect 580258 144888 580264 144900
rect 560076 144860 580264 144888
rect 560076 144848 560082 144860
rect 580258 144848 580264 144860
rect 580316 144848 580322 144900
rect 191190 144712 191196 144764
rect 191248 144752 191254 144764
rect 194594 144752 194600 144764
rect 191248 144724 194600 144752
rect 191248 144712 191254 144724
rect 194594 144712 194600 144724
rect 194652 144752 194658 144764
rect 197354 144752 197360 144764
rect 194652 144724 197360 144752
rect 194652 144712 194658 144724
rect 197354 144712 197360 144724
rect 197412 144712 197418 144764
rect 177850 144168 177856 144220
rect 177908 144208 177914 144220
rect 194594 144208 194600 144220
rect 177908 144180 194600 144208
rect 177908 144168 177914 144180
rect 194594 144168 194600 144180
rect 194652 144168 194658 144220
rect 194594 143556 194600 143608
rect 194652 143596 194658 143608
rect 197354 143596 197360 143608
rect 194652 143568 197360 143596
rect 194652 143556 194658 143568
rect 197354 143556 197360 143568
rect 197412 143556 197418 143608
rect 178954 142808 178960 142860
rect 179012 142848 179018 142860
rect 186314 142848 186320 142860
rect 179012 142820 186320 142848
rect 179012 142808 179018 142820
rect 186314 142808 186320 142820
rect 186372 142808 186378 142860
rect 186314 142128 186320 142180
rect 186372 142168 186378 142180
rect 197354 142168 197360 142180
rect 186372 142140 197360 142168
rect 186372 142128 186378 142140
rect 197354 142128 197360 142140
rect 197412 142128 197418 142180
rect 166166 141448 166172 141500
rect 166224 141488 166230 141500
rect 197814 141488 197820 141500
rect 166224 141460 197820 141488
rect 166224 141448 166230 141460
rect 197814 141448 197820 141460
rect 197872 141448 197878 141500
rect 166258 141380 166264 141432
rect 166316 141420 166322 141432
rect 197446 141420 197452 141432
rect 166316 141392 197452 141420
rect 166316 141380 166322 141392
rect 197446 141380 197452 141392
rect 197504 141380 197510 141432
rect 133138 141312 133144 141364
rect 133196 141352 133202 141364
rect 168098 141352 168104 141364
rect 133196 141324 168104 141352
rect 133196 141312 133202 141324
rect 168098 141312 168104 141324
rect 168156 141312 168162 141364
rect 140038 141244 140044 141296
rect 140096 141284 140102 141296
rect 181622 141284 181628 141296
rect 140096 141256 181628 141284
rect 140096 141244 140102 141256
rect 181622 141244 181628 141256
rect 181680 141244 181686 141296
rect 128538 141176 128544 141228
rect 128596 141216 128602 141228
rect 176194 141216 176200 141228
rect 128596 141188 176200 141216
rect 128596 141176 128602 141188
rect 176194 141176 176200 141188
rect 176252 141176 176258 141228
rect 142338 141108 142344 141160
rect 142396 141148 142402 141160
rect 190454 141148 190460 141160
rect 142396 141120 190460 141148
rect 142396 141108 142402 141120
rect 190454 141108 190460 141120
rect 190512 141108 190518 141160
rect 134242 141040 134248 141092
rect 134300 141080 134306 141092
rect 187878 141080 187884 141092
rect 134300 141052 187884 141080
rect 134300 141040 134306 141052
rect 187878 141040 187884 141052
rect 187936 141040 187942 141092
rect 123754 140972 123760 141024
rect 123812 141012 123818 141024
rect 178126 141012 178132 141024
rect 123812 140984 178132 141012
rect 123812 140972 123818 140984
rect 178126 140972 178132 140984
rect 178184 140972 178190 141024
rect 136542 140904 136548 140956
rect 136600 140944 136606 140956
rect 193306 140944 193312 140956
rect 136600 140916 193312 140944
rect 136600 140904 136606 140916
rect 193306 140904 193312 140916
rect 193364 140904 193370 140956
rect 112162 140836 112168 140888
rect 112220 140876 112226 140888
rect 171778 140876 171784 140888
rect 112220 140848 171784 140876
rect 112220 140836 112226 140848
rect 171778 140836 171784 140848
rect 171836 140836 171842 140888
rect 108482 140768 108488 140820
rect 108540 140808 108546 140820
rect 176102 140808 176108 140820
rect 108540 140780 176108 140808
rect 108540 140768 108546 140780
rect 176102 140768 176108 140780
rect 176160 140768 176166 140820
rect 137922 140700 137928 140752
rect 137980 140740 137986 140752
rect 168282 140740 168288 140752
rect 137980 140712 168288 140740
rect 137980 140700 137986 140712
rect 168282 140700 168288 140712
rect 168340 140700 168346 140752
rect 135346 140632 135352 140684
rect 135404 140672 135410 140684
rect 168190 140672 168196 140684
rect 135404 140644 168196 140672
rect 135404 140632 135410 140644
rect 168190 140632 168196 140644
rect 168248 140632 168254 140684
rect 141234 140564 141240 140616
rect 141292 140604 141298 140616
rect 174906 140604 174912 140616
rect 141292 140576 174912 140604
rect 141292 140564 141298 140576
rect 174906 140564 174912 140576
rect 174964 140564 174970 140616
rect 139026 140496 139032 140548
rect 139084 140536 139090 140548
rect 173434 140536 173440 140548
rect 139084 140508 173440 140536
rect 139084 140496 139090 140508
rect 173434 140496 173440 140508
rect 173492 140496 173498 140548
rect 143442 140428 143448 140480
rect 143500 140468 143506 140480
rect 177758 140468 177764 140480
rect 143500 140440 177764 140468
rect 143500 140428 143506 140440
rect 177758 140428 177764 140440
rect 177816 140428 177822 140480
rect 132034 140360 132040 140412
rect 132092 140400 132098 140412
rect 168006 140400 168012 140412
rect 132092 140372 168012 140400
rect 132092 140360 132098 140372
rect 168006 140360 168012 140372
rect 168064 140360 168070 140412
rect 125962 140292 125968 140344
rect 126020 140332 126026 140344
rect 170766 140332 170772 140344
rect 126020 140304 170772 140332
rect 126020 140292 126026 140304
rect 170766 140292 170772 140304
rect 170824 140292 170830 140344
rect 118970 140224 118976 140276
rect 119028 140264 119034 140276
rect 171042 140264 171048 140276
rect 119028 140236 171048 140264
rect 119028 140224 119034 140236
rect 171042 140224 171048 140236
rect 171100 140224 171106 140276
rect 116762 140156 116768 140208
rect 116820 140196 116826 140208
rect 184382 140196 184388 140208
rect 116820 140168 184388 140196
rect 116820 140156 116826 140168
rect 184382 140156 184388 140168
rect 184440 140156 184446 140208
rect 29822 140088 29828 140140
rect 29880 140128 29886 140140
rect 35894 140128 35900 140140
rect 29880 140100 35900 140128
rect 29880 140088 29886 140100
rect 35894 140088 35900 140100
rect 35952 140088 35958 140140
rect 113266 140088 113272 140140
rect 113324 140128 113330 140140
rect 185026 140128 185032 140140
rect 113324 140100 185032 140128
rect 113324 140088 113330 140100
rect 185026 140088 185032 140100
rect 185084 140088 185090 140140
rect 109586 140020 109592 140072
rect 109644 140060 109650 140072
rect 191926 140060 191932 140072
rect 109644 140032 191932 140060
rect 109644 140020 109650 140032
rect 191926 140020 191932 140032
rect 191984 140020 191990 140072
rect 167822 139952 167828 140004
rect 167880 139992 167886 140004
rect 197354 139992 197360 140004
rect 167880 139964 197360 139992
rect 167880 139952 167886 139964
rect 197354 139952 197360 139964
rect 197412 139952 197418 140004
rect 166994 139884 167000 139936
rect 167052 139924 167058 139936
rect 197262 139924 197268 139936
rect 167052 139896 197268 139924
rect 167052 139884 167058 139896
rect 197262 139884 197268 139896
rect 197320 139884 197326 139936
rect 149514 139408 149520 139460
rect 149572 139448 149578 139460
rect 166994 139448 167000 139460
rect 149572 139420 167000 139448
rect 149572 139408 149578 139420
rect 166994 139408 167000 139420
rect 167052 139408 167058 139460
rect 120350 139340 120356 139392
rect 120408 139380 120414 139392
rect 191282 139380 191288 139392
rect 120408 139352 191288 139380
rect 120408 139340 120414 139352
rect 191282 139340 191288 139352
rect 191340 139340 191346 139392
rect 559558 139340 559564 139392
rect 559616 139380 559622 139392
rect 580166 139380 580172 139392
rect 559616 139352 580172 139380
rect 559616 139340 559622 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 129642 139272 129648 139324
rect 129700 139312 129706 139324
rect 196066 139312 196072 139324
rect 129700 139284 196072 139312
rect 129700 139272 129706 139284
rect 196066 139272 196072 139284
rect 196124 139272 196130 139324
rect 121362 139204 121368 139256
rect 121420 139244 121426 139256
rect 182910 139244 182916 139256
rect 121420 139216 182916 139244
rect 121420 139204 121426 139216
rect 182910 139204 182916 139216
rect 182968 139204 182974 139256
rect 115474 139136 115480 139188
rect 115532 139176 115538 139188
rect 174814 139176 174820 139188
rect 115532 139148 174820 139176
rect 115532 139136 115538 139148
rect 174814 139136 174820 139148
rect 174872 139136 174878 139188
rect 107378 139068 107384 139120
rect 107436 139108 107442 139120
rect 166258 139108 166264 139120
rect 107436 139080 166264 139108
rect 107436 139068 107442 139080
rect 166258 139068 166264 139080
rect 166316 139068 166322 139120
rect 114370 139000 114376 139052
rect 114428 139040 114434 139052
rect 171870 139040 171876 139052
rect 114428 139012 171876 139040
rect 114428 139000 114434 139012
rect 171870 139000 171876 139012
rect 171928 139000 171934 139052
rect 110874 138932 110880 138984
rect 110932 138972 110938 138984
rect 169018 138972 169024 138984
rect 110932 138944 169024 138972
rect 110932 138932 110938 138944
rect 169018 138932 169024 138944
rect 169076 138932 169082 138984
rect 122650 138864 122656 138916
rect 122708 138904 122714 138916
rect 179414 138904 179420 138916
rect 122708 138876 179420 138904
rect 122708 138864 122714 138876
rect 179414 138864 179420 138876
rect 179472 138864 179478 138916
rect 28810 138796 28816 138848
rect 28868 138836 28874 138848
rect 43438 138836 43444 138848
rect 28868 138808 43444 138836
rect 28868 138796 28874 138808
rect 43438 138796 43444 138808
rect 43496 138796 43502 138848
rect 130746 138796 130752 138848
rect 130804 138836 130810 138848
rect 186498 138836 186504 138848
rect 130804 138808 186504 138836
rect 130804 138796 130810 138808
rect 186498 138796 186504 138808
rect 186556 138796 186562 138848
rect 117866 138728 117872 138780
rect 117924 138768 117930 138780
rect 169202 138768 169208 138780
rect 117924 138740 169208 138768
rect 117924 138728 117930 138740
rect 169202 138728 169208 138740
rect 169260 138728 169266 138780
rect 28626 138660 28632 138712
rect 28684 138700 28690 138712
rect 43070 138700 43076 138712
rect 28684 138672 43076 138700
rect 28684 138660 28690 138672
rect 43070 138660 43076 138672
rect 43128 138660 43134 138712
rect 127710 138660 127716 138712
rect 127768 138700 127774 138712
rect 170950 138700 170956 138712
rect 127768 138672 170956 138700
rect 127768 138660 127774 138672
rect 170950 138660 170956 138672
rect 171008 138660 171014 138712
rect 125226 138592 125232 138644
rect 125284 138632 125290 138644
rect 167914 138632 167920 138644
rect 125284 138604 167920 138632
rect 125284 138592 125290 138604
rect 167914 138592 167920 138604
rect 167972 138592 167978 138644
rect 28350 138524 28356 138576
rect 28408 138564 28414 138576
rect 28810 138564 28816 138576
rect 28408 138536 28816 138564
rect 28408 138524 28414 138536
rect 28810 138524 28816 138536
rect 28868 138524 28874 138576
rect 148410 138524 148416 138576
rect 148468 138564 148474 138576
rect 166166 138564 166172 138576
rect 148468 138536 166172 138564
rect 148468 138524 148474 138536
rect 166166 138524 166172 138536
rect 166224 138524 166230 138576
rect 151078 138456 151084 138508
rect 151136 138496 151142 138508
rect 167086 138496 167092 138508
rect 151136 138468 167092 138496
rect 151136 138456 151142 138468
rect 167086 138456 167092 138468
rect 167144 138456 167150 138508
rect 167086 138252 167092 138304
rect 167144 138292 167150 138304
rect 167822 138292 167828 138304
rect 167144 138264 167828 138292
rect 167144 138252 167150 138264
rect 167822 138252 167828 138264
rect 167880 138252 167886 138304
rect 60642 137980 60648 138032
rect 60700 138020 60706 138032
rect 117222 138020 117228 138032
rect 60700 137992 117228 138020
rect 60700 137980 60706 137992
rect 117222 137980 117228 137992
rect 117280 137980 117286 138032
rect 3326 137912 3332 137964
rect 3384 137952 3390 137964
rect 181438 137952 181444 137964
rect 3384 137924 181444 137952
rect 3384 137912 3390 137924
rect 181438 137912 181444 137924
rect 181496 137912 181502 137964
rect 63218 137844 63224 137896
rect 63276 137884 63282 137896
rect 197354 137884 197360 137896
rect 63276 137856 197360 137884
rect 63276 137844 63282 137856
rect 197354 137844 197360 137856
rect 197412 137844 197418 137896
rect 117222 137776 117228 137828
rect 117280 137816 117286 137828
rect 197446 137816 197452 137828
rect 117280 137788 197452 137816
rect 117280 137776 117286 137788
rect 197446 137776 197452 137788
rect 197504 137776 197510 137828
rect 164878 136824 164884 136876
rect 164936 136864 164942 136876
rect 168558 136864 168564 136876
rect 164936 136836 168564 136864
rect 164936 136824 164942 136836
rect 168558 136824 168564 136836
rect 168616 136824 168622 136876
rect 65794 136552 65800 136604
rect 65852 136592 65858 136604
rect 197354 136592 197360 136604
rect 65852 136564 197360 136592
rect 65852 136552 65858 136564
rect 197354 136552 197360 136564
rect 197412 136552 197418 136604
rect 136450 135872 136456 135924
rect 136508 135912 136514 135924
rect 194042 135912 194048 135924
rect 136508 135884 194048 135912
rect 136508 135872 136514 135884
rect 194042 135872 194048 135884
rect 194100 135872 194106 135924
rect 559282 135328 559288 135380
rect 559340 135368 559346 135380
rect 560938 135368 560944 135380
rect 559340 135340 560944 135368
rect 559340 135328 559346 135340
rect 560938 135328 560944 135340
rect 560996 135328 561002 135380
rect 68922 135192 68928 135244
rect 68980 135232 68986 135244
rect 197354 135232 197360 135244
rect 68980 135204 197360 135232
rect 68980 135192 68986 135204
rect 197354 135192 197360 135204
rect 197412 135192 197418 135244
rect 124122 134512 124128 134564
rect 124180 134552 124186 134564
rect 178954 134552 178960 134564
rect 124180 134524 178960 134552
rect 124180 134512 124186 134524
rect 178954 134512 178960 134524
rect 179012 134512 179018 134564
rect 71038 133832 71044 133884
rect 71096 133872 71102 133884
rect 197354 133872 197360 133884
rect 71096 133844 197360 133872
rect 71096 133832 71102 133844
rect 197354 133832 197360 133844
rect 197412 133832 197418 133884
rect 118418 133152 118424 133204
rect 118476 133192 118482 133204
rect 180242 133192 180248 133204
rect 118476 133164 180248 133192
rect 118476 133152 118482 133164
rect 180242 133152 180248 133164
rect 180300 133152 180306 133204
rect 74442 132404 74448 132456
rect 74500 132444 74506 132456
rect 197354 132444 197360 132456
rect 74500 132416 197360 132444
rect 74500 132404 74506 132416
rect 197354 132404 197360 132416
rect 197412 132404 197418 132456
rect 75822 132336 75828 132388
rect 75880 132376 75886 132388
rect 197446 132376 197452 132388
rect 75880 132348 197452 132376
rect 75880 132336 75886 132348
rect 197446 132336 197452 132348
rect 197504 132336 197510 132388
rect 78582 131044 78588 131096
rect 78640 131084 78646 131096
rect 197354 131084 197360 131096
rect 78640 131056 197360 131084
rect 78640 131044 78646 131056
rect 197354 131044 197360 131056
rect 197412 131044 197418 131096
rect 121362 130364 121368 130416
rect 121420 130404 121426 130416
rect 181438 130404 181444 130416
rect 121420 130376 181444 130404
rect 121420 130364 121426 130376
rect 181438 130364 181444 130376
rect 181496 130364 181502 130416
rect 81342 129684 81348 129736
rect 81400 129724 81406 129736
rect 197354 129724 197360 129736
rect 81400 129696 197360 129724
rect 81400 129684 81406 129696
rect 197354 129684 197360 129696
rect 197412 129684 197418 129736
rect 125410 129004 125416 129056
rect 125468 129044 125474 129056
rect 174814 129044 174820 129056
rect 125468 129016 174820 129044
rect 125468 129004 125474 129016
rect 174814 129004 174820 129016
rect 174872 129004 174878 129056
rect 84102 128256 84108 128308
rect 84160 128296 84166 128308
rect 197354 128296 197360 128308
rect 84160 128268 197360 128296
rect 84160 128256 84166 128268
rect 197354 128256 197360 128268
rect 197412 128256 197418 128308
rect 128262 127576 128268 127628
rect 128320 127616 128326 127628
rect 177758 127616 177764 127628
rect 128320 127588 177764 127616
rect 128320 127576 128326 127588
rect 177758 127576 177764 127588
rect 177816 127576 177822 127628
rect 86862 126896 86868 126948
rect 86920 126936 86926 126948
rect 197354 126936 197360 126948
rect 86920 126908 197360 126936
rect 86920 126896 86926 126908
rect 197354 126896 197360 126908
rect 197412 126896 197418 126948
rect 560938 126896 560944 126948
rect 560996 126936 561002 126948
rect 580166 126936 580172 126948
rect 560996 126908 580172 126936
rect 560996 126896 561002 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 133782 126284 133788 126336
rect 133840 126324 133846 126336
rect 167822 126324 167828 126336
rect 133840 126296 167828 126324
rect 133840 126284 133846 126296
rect 167822 126284 167828 126296
rect 167880 126284 167886 126336
rect 115842 126216 115848 126268
rect 115900 126256 115906 126268
rect 184382 126256 184388 126268
rect 115900 126228 184388 126256
rect 115900 126216 115906 126228
rect 184382 126216 184388 126228
rect 184440 126216 184446 126268
rect 88242 125536 88248 125588
rect 88300 125576 88306 125588
rect 197354 125576 197360 125588
rect 88300 125548 197360 125576
rect 88300 125536 88306 125548
rect 197354 125536 197360 125548
rect 197412 125536 197418 125588
rect 131022 124856 131028 124908
rect 131080 124896 131086 124908
rect 174906 124896 174912 124908
rect 131080 124868 174912 124896
rect 131080 124856 131086 124868
rect 174906 124856 174912 124868
rect 174964 124856 174970 124908
rect 91002 124108 91008 124160
rect 91060 124148 91066 124160
rect 197354 124148 197360 124160
rect 91060 124120 197360 124148
rect 91060 124108 91066 124120
rect 197354 124108 197360 124120
rect 197412 124108 197418 124160
rect 139302 123496 139308 123548
rect 139360 123536 139366 123548
rect 180334 123536 180340 123548
rect 139360 123508 180340 123536
rect 139360 123496 139366 123508
rect 180334 123496 180340 123508
rect 180392 123496 180398 123548
rect 113082 123428 113088 123480
rect 113140 123468 113146 123480
rect 171778 123468 171784 123480
rect 113140 123440 171784 123468
rect 113140 123428 113146 123440
rect 171778 123428 171784 123440
rect 171836 123428 171842 123480
rect 93762 122748 93768 122800
rect 93820 122788 93826 122800
rect 197354 122788 197360 122800
rect 93820 122760 197360 122788
rect 93820 122748 93826 122760
rect 197354 122748 197360 122760
rect 197412 122748 197418 122800
rect 96522 121388 96528 121440
rect 96580 121428 96586 121440
rect 197354 121428 197360 121440
rect 96580 121400 197360 121428
rect 96580 121388 96586 121400
rect 197354 121388 197360 121400
rect 197412 121388 197418 121440
rect 99282 120028 99288 120080
rect 99340 120068 99346 120080
rect 197354 120068 197360 120080
rect 99340 120040 197360 120068
rect 99340 120028 99346 120040
rect 197354 120028 197360 120040
rect 197412 120028 197418 120080
rect 100662 119960 100668 120012
rect 100720 120000 100726 120012
rect 197446 120000 197452 120012
rect 100720 119972 197452 120000
rect 100720 119960 100726 119972
rect 197446 119960 197452 119972
rect 197504 119960 197510 120012
rect 558914 118668 558920 118720
rect 558972 118708 558978 118720
rect 561030 118708 561036 118720
rect 558972 118680 561036 118708
rect 558972 118668 558978 118680
rect 561030 118668 561036 118680
rect 561088 118668 561094 118720
rect 103422 118600 103428 118652
rect 103480 118640 103486 118652
rect 197354 118640 197360 118652
rect 103480 118612 197360 118640
rect 103480 118600 103486 118612
rect 197354 118600 197360 118612
rect 197412 118600 197418 118652
rect 35894 117240 35900 117292
rect 35952 117280 35958 117292
rect 164878 117280 164884 117292
rect 35952 117252 164884 117280
rect 35952 117240 35958 117252
rect 164878 117240 164884 117252
rect 164936 117280 164942 117292
rect 168558 117280 168564 117292
rect 164936 117252 168564 117280
rect 164936 117240 164942 117252
rect 168558 117240 168564 117252
rect 168616 117240 168622 117292
rect 28718 117172 28724 117224
rect 28776 117212 28782 117224
rect 46934 117212 46940 117224
rect 28776 117184 46940 117212
rect 28776 117172 28782 117184
rect 46934 117172 46940 117184
rect 46992 117172 46998 117224
rect 106182 117172 106188 117224
rect 106240 117212 106246 117224
rect 197354 117212 197360 117224
rect 106240 117184 197360 117212
rect 106240 117172 106246 117184
rect 197354 117172 197360 117184
rect 197412 117172 197418 117224
rect 28534 117104 28540 117156
rect 28592 117144 28598 117156
rect 45830 117144 45836 117156
rect 28592 117116 45836 117144
rect 28592 117104 28598 117116
rect 45830 117104 45836 117116
rect 45888 117104 45894 117156
rect 108942 115880 108948 115932
rect 109000 115920 109006 115932
rect 197354 115920 197360 115932
rect 109000 115892 197360 115920
rect 109000 115880 109006 115892
rect 197354 115880 197360 115892
rect 197412 115880 197418 115932
rect 3786 115336 3792 115388
rect 3844 115376 3850 115388
rect 173250 115376 173256 115388
rect 3844 115348 173256 115376
rect 3844 115336 3850 115348
rect 173250 115336 173256 115348
rect 173308 115336 173314 115388
rect 3878 115268 3884 115320
rect 3936 115308 3942 115320
rect 193858 115308 193864 115320
rect 3936 115280 193864 115308
rect 3936 115268 3942 115280
rect 193858 115268 193864 115280
rect 193916 115268 193922 115320
rect 3602 115200 3608 115252
rect 3660 115240 3666 115252
rect 196710 115240 196716 115252
rect 3660 115212 196716 115240
rect 3660 115200 3666 115212
rect 196710 115200 196716 115212
rect 196768 115200 196774 115252
rect 111702 114452 111708 114504
rect 111760 114492 111766 114504
rect 197354 114492 197360 114504
rect 111760 114464 197360 114492
rect 111760 114452 111766 114464
rect 197354 114452 197360 114464
rect 197412 114452 197418 114504
rect 3694 113840 3700 113892
rect 3752 113880 3758 113892
rect 173158 113880 173164 113892
rect 3752 113852 173164 113880
rect 3752 113840 3758 113852
rect 173158 113840 173164 113852
rect 173216 113840 173222 113892
rect 4062 113772 4068 113824
rect 4120 113812 4126 113824
rect 196618 113812 196624 113824
rect 4120 113784 196624 113812
rect 4120 113772 4126 113784
rect 196618 113772 196624 113784
rect 196676 113772 196682 113824
rect 171778 113092 171784 113144
rect 171836 113132 171842 113144
rect 197354 113132 197360 113144
rect 171836 113104 197360 113132
rect 171836 113092 171842 113104
rect 197354 113092 197360 113104
rect 197412 113092 197418 113144
rect 561030 113092 561036 113144
rect 561088 113132 561094 113144
rect 579798 113132 579804 113144
rect 561088 113104 579804 113132
rect 561088 113092 561094 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 559190 111800 559196 111852
rect 559248 111840 559254 111852
rect 560938 111840 560944 111852
rect 559248 111812 560944 111840
rect 559248 111800 559254 111812
rect 560938 111800 560944 111812
rect 560996 111800 561002 111852
rect 184382 111732 184388 111784
rect 184440 111772 184446 111784
rect 197354 111772 197360 111784
rect 184440 111744 197360 111772
rect 184440 111732 184446 111744
rect 197354 111732 197360 111744
rect 197412 111732 197418 111784
rect 180242 110372 180248 110424
rect 180300 110412 180306 110424
rect 197354 110412 197360 110424
rect 180300 110384 197360 110412
rect 180300 110372 180306 110384
rect 197354 110372 197360 110384
rect 197412 110372 197418 110424
rect 178954 108944 178960 108996
rect 179012 108984 179018 108996
rect 197538 108984 197544 108996
rect 179012 108956 197544 108984
rect 179012 108944 179018 108956
rect 197538 108944 197544 108956
rect 197596 108944 197602 108996
rect 181438 108876 181444 108928
rect 181496 108916 181502 108928
rect 197354 108916 197360 108928
rect 181496 108888 197360 108916
rect 181496 108876 181502 108888
rect 197354 108876 197360 108888
rect 197412 108876 197418 108928
rect 174814 107584 174820 107636
rect 174872 107624 174878 107636
rect 197446 107624 197452 107636
rect 174872 107596 197452 107624
rect 174872 107584 174878 107596
rect 197446 107584 197452 107596
rect 197504 107584 197510 107636
rect 177758 106224 177764 106276
rect 177816 106264 177822 106276
rect 197354 106264 197360 106276
rect 177816 106236 197360 106264
rect 177816 106224 177822 106236
rect 197354 106224 197360 106236
rect 197412 106224 197418 106276
rect 174906 104796 174912 104848
rect 174964 104836 174970 104848
rect 197354 104836 197360 104848
rect 174964 104808 197360 104836
rect 174964 104796 174970 104808
rect 197354 104796 197360 104808
rect 197412 104796 197418 104848
rect 560202 103776 560208 103828
rect 560260 103816 560266 103828
rect 566458 103816 566464 103828
rect 560260 103788 566464 103816
rect 560260 103776 560266 103788
rect 566458 103776 566464 103788
rect 566516 103776 566522 103828
rect 167822 103436 167828 103488
rect 167880 103476 167886 103488
rect 197354 103476 197360 103488
rect 167880 103448 197360 103476
rect 167880 103436 167886 103448
rect 197354 103436 197360 103448
rect 197412 103436 197418 103488
rect 194042 102076 194048 102128
rect 194100 102116 194106 102128
rect 197354 102116 197360 102128
rect 194100 102088 197360 102116
rect 194100 102076 194106 102088
rect 197354 102076 197360 102088
rect 197412 102076 197418 102128
rect 180334 100648 180340 100700
rect 180392 100688 180398 100700
rect 197354 100688 197360 100700
rect 180392 100660 197360 100688
rect 180392 100648 180398 100660
rect 197354 100648 197360 100660
rect 197412 100648 197418 100700
rect 559558 100648 559564 100700
rect 559616 100688 559622 100700
rect 580166 100688 580172 100700
rect 559616 100660 580172 100688
rect 559616 100648 559622 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 167822 97996 167828 98048
rect 167880 98036 167886 98048
rect 197354 98036 197360 98048
rect 167880 98008 197360 98036
rect 167880 97996 167886 98008
rect 197354 97996 197360 98008
rect 197412 97996 197418 98048
rect 559742 95208 559748 95260
rect 559800 95248 559806 95260
rect 565078 95248 565084 95260
rect 559800 95220 565084 95248
rect 559800 95208 559806 95220
rect 565078 95208 565084 95220
rect 565136 95208 565142 95260
rect 178954 93848 178960 93900
rect 179012 93888 179018 93900
rect 197354 93888 197360 93900
rect 179012 93860 197360 93888
rect 179012 93848 179018 93860
rect 197354 93848 197360 93860
rect 197412 93848 197418 93900
rect 167914 92488 167920 92540
rect 167972 92528 167978 92540
rect 197354 92528 197360 92540
rect 167972 92500 197360 92528
rect 167972 92488 167978 92500
rect 197354 92488 197360 92500
rect 197412 92488 197418 92540
rect 176102 91060 176108 91112
rect 176160 91100 176166 91112
rect 197354 91100 197360 91112
rect 176160 91072 197360 91100
rect 176160 91060 176166 91072
rect 197354 91060 197360 91072
rect 197412 91060 197418 91112
rect 177758 89700 177764 89752
rect 177816 89740 177822 89752
rect 197354 89740 197360 89752
rect 177816 89712 197360 89740
rect 177816 89700 177822 89712
rect 197354 89700 197360 89712
rect 197412 89700 197418 89752
rect 176194 88340 176200 88392
rect 176252 88380 176258 88392
rect 197354 88380 197360 88392
rect 176252 88352 197360 88380
rect 176252 88340 176258 88352
rect 197354 88340 197360 88352
rect 197412 88340 197418 88392
rect 174814 86980 174820 87032
rect 174872 87020 174878 87032
rect 197354 87020 197360 87032
rect 174872 86992 197360 87020
rect 174872 86980 174878 86992
rect 197354 86980 197360 86992
rect 197412 86980 197418 87032
rect 560202 86980 560208 87032
rect 560260 87020 560266 87032
rect 574830 87020 574836 87032
rect 560260 86992 574836 87020
rect 560260 86980 560266 86992
rect 574830 86980 574836 86992
rect 574888 86980 574894 87032
rect 560938 86912 560944 86964
rect 560996 86952 561002 86964
rect 580166 86952 580172 86964
rect 560996 86924 580172 86952
rect 560996 86912 561002 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 173158 85552 173164 85604
rect 173216 85592 173222 85604
rect 197354 85592 197360 85604
rect 173216 85564 197360 85592
rect 173216 85552 173222 85564
rect 197354 85552 197360 85564
rect 197412 85552 197418 85604
rect 169018 84192 169024 84244
rect 169076 84232 169082 84244
rect 197354 84232 197360 84244
rect 169076 84204 197360 84232
rect 169076 84192 169082 84204
rect 197354 84192 197360 84204
rect 197412 84192 197418 84244
rect 168006 82832 168012 82884
rect 168064 82872 168070 82884
rect 197354 82872 197360 82884
rect 168064 82844 197360 82872
rect 168064 82832 168070 82844
rect 197354 82832 197360 82844
rect 197412 82832 197418 82884
rect 174906 81472 174912 81524
rect 174964 81512 174970 81524
rect 197446 81512 197452 81524
rect 174964 81484 197452 81512
rect 174964 81472 174970 81484
rect 197446 81472 197452 81484
rect 197504 81472 197510 81524
rect 173250 81404 173256 81456
rect 173308 81444 173314 81456
rect 197354 81444 197360 81456
rect 173308 81416 197360 81444
rect 173308 81404 173314 81416
rect 197354 81404 197360 81416
rect 197412 81404 197418 81456
rect 174998 80044 175004 80096
rect 175056 80084 175062 80096
rect 197354 80084 197360 80096
rect 175056 80056 197360 80084
rect 175056 80044 175062 80056
rect 197354 80044 197360 80056
rect 197412 80044 197418 80096
rect 169110 78684 169116 78736
rect 169168 78724 169174 78736
rect 197354 78724 197360 78736
rect 169168 78696 197360 78724
rect 169168 78684 169174 78696
rect 197354 78684 197360 78696
rect 197412 78684 197418 78736
rect 560018 78684 560024 78736
rect 560076 78724 560082 78736
rect 577498 78724 577504 78736
rect 560076 78696 577504 78724
rect 560076 78684 560082 78696
rect 577498 78684 577504 78696
rect 577556 78684 577562 78736
rect 168190 77256 168196 77308
rect 168248 77296 168254 77308
rect 197354 77296 197360 77308
rect 168248 77268 197360 77296
rect 168248 77256 168254 77268
rect 197354 77256 197360 77268
rect 197412 77256 197418 77308
rect 171778 75896 171784 75948
rect 171836 75936 171842 75948
rect 197354 75936 197360 75948
rect 171836 75908 197360 75936
rect 171836 75896 171842 75908
rect 197354 75896 197360 75908
rect 197412 75896 197418 75948
rect 168098 74536 168104 74588
rect 168156 74576 168162 74588
rect 197354 74576 197360 74588
rect 168156 74548 197360 74576
rect 168156 74536 168162 74548
rect 197354 74536 197360 74548
rect 197412 74536 197418 74588
rect 169202 73176 169208 73228
rect 169260 73216 169266 73228
rect 197354 73216 197360 73228
rect 169260 73188 197360 73216
rect 169260 73176 169266 73188
rect 197354 73176 197360 73188
rect 197412 73176 197418 73228
rect 565078 73108 565084 73160
rect 565136 73148 565142 73160
rect 580166 73148 580172 73160
rect 565136 73120 580172 73148
rect 565136 73108 565142 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 559190 71816 559196 71868
rect 559248 71856 559254 71868
rect 560938 71856 560944 71868
rect 559248 71828 560944 71856
rect 559248 71816 559254 71828
rect 560938 71816 560944 71828
rect 560996 71816 561002 71868
rect 173434 71748 173440 71800
rect 173492 71788 173498 71800
rect 197354 71788 197360 71800
rect 173492 71760 197360 71788
rect 173492 71748 173498 71760
rect 197354 71748 197360 71760
rect 197412 71748 197418 71800
rect 176286 70388 176292 70440
rect 176344 70428 176350 70440
rect 197354 70428 197360 70440
rect 176344 70400 197360 70428
rect 176344 70388 176350 70400
rect 197354 70388 197360 70400
rect 197412 70388 197418 70440
rect 168834 69640 168840 69692
rect 168892 69680 168898 69692
rect 187694 69680 187700 69692
rect 168892 69652 187700 69680
rect 168892 69640 168898 69652
rect 187694 69640 187700 69652
rect 187752 69640 187758 69692
rect 168834 66172 168840 66224
rect 168892 66212 168898 66224
rect 180794 66212 180800 66224
rect 168892 66184 180800 66212
rect 168892 66172 168898 66184
rect 180794 66172 180800 66184
rect 180852 66172 180858 66224
rect 168834 64812 168840 64864
rect 168892 64852 168898 64864
rect 177666 64852 177672 64864
rect 168892 64824 177672 64852
rect 168892 64812 168898 64824
rect 177666 64812 177672 64824
rect 177724 64812 177730 64864
rect 168926 64132 168932 64184
rect 168984 64172 168990 64184
rect 191190 64172 191196 64184
rect 168984 64144 191196 64172
rect 168984 64132 168990 64144
rect 191190 64132 191196 64144
rect 191248 64132 191254 64184
rect 170950 63520 170956 63572
rect 171008 63560 171014 63572
rect 197354 63560 197360 63572
rect 171008 63532 197360 63560
rect 171008 63520 171014 63532
rect 197354 63520 197360 63532
rect 197412 63520 197418 63572
rect 560202 63520 560208 63572
rect 560260 63560 560266 63572
rect 570598 63560 570604 63572
rect 560260 63532 570604 63560
rect 560260 63520 560266 63532
rect 570598 63520 570604 63532
rect 570656 63520 570662 63572
rect 169386 63452 169392 63504
rect 169444 63492 169450 63504
rect 178034 63492 178040 63504
rect 169444 63464 178040 63492
rect 169444 63452 169450 63464
rect 178034 63452 178040 63464
rect 178092 63452 178098 63504
rect 168834 61344 168840 61396
rect 168892 61384 168898 61396
rect 194594 61384 194600 61396
rect 168892 61356 194600 61384
rect 168892 61344 168898 61356
rect 194594 61344 194600 61356
rect 194652 61344 194658 61396
rect 172054 60732 172060 60784
rect 172112 60772 172118 60784
rect 197354 60772 197360 60784
rect 172112 60744 197360 60772
rect 172112 60732 172118 60744
rect 197354 60732 197360 60744
rect 197412 60732 197418 60784
rect 566458 60664 566464 60716
rect 566516 60704 566522 60716
rect 580166 60704 580172 60716
rect 566516 60676 580172 60704
rect 566516 60664 566522 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 169294 59372 169300 59424
rect 169352 59412 169358 59424
rect 197538 59412 197544 59424
rect 169352 59384 197544 59412
rect 169352 59372 169358 59384
rect 197538 59372 197544 59384
rect 197596 59372 197602 59424
rect 168834 59304 168840 59356
rect 168892 59344 168898 59356
rect 186314 59344 186320 59356
rect 168892 59316 186320 59344
rect 168892 59304 168898 59316
rect 186314 59304 186320 59316
rect 186372 59304 186378 59356
rect 560938 58624 560944 58676
rect 560996 58664 561002 58676
rect 580350 58664 580356 58676
rect 560996 58636 580356 58664
rect 560996 58624 561002 58636
rect 580350 58624 580356 58636
rect 580408 58624 580414 58676
rect 201236 58092 202184 58120
rect 196618 57808 196624 57860
rect 196676 57848 196682 57860
rect 201236 57848 201264 58092
rect 201494 58012 201500 58064
rect 201552 58052 201558 58064
rect 202046 58052 202052 58064
rect 201552 58024 202052 58052
rect 201552 58012 201558 58024
rect 202046 58012 202052 58024
rect 202104 58012 202110 58064
rect 196676 57820 201264 57848
rect 201328 57956 201724 57984
rect 196676 57808 196682 57820
rect 181438 57740 181444 57792
rect 181496 57780 181502 57792
rect 201328 57780 201356 57956
rect 181496 57752 201356 57780
rect 201696 57780 201724 57956
rect 202156 57916 202184 58092
rect 206738 57916 206744 57928
rect 202156 57888 206744 57916
rect 206738 57876 206744 57888
rect 206796 57876 206802 57928
rect 211798 57780 211804 57792
rect 201696 57752 211804 57780
rect 181496 57740 181502 57752
rect 211798 57740 211804 57752
rect 211856 57740 211862 57792
rect 214650 57740 214656 57792
rect 214708 57780 214714 57792
rect 224126 57780 224132 57792
rect 214708 57752 224132 57780
rect 214708 57740 214714 57752
rect 224126 57740 224132 57752
rect 224184 57740 224190 57792
rect 471238 57740 471244 57792
rect 471296 57780 471302 57792
rect 477678 57780 477684 57792
rect 471296 57752 477684 57780
rect 471296 57740 471302 57752
rect 477678 57740 477684 57752
rect 477736 57740 477742 57792
rect 480898 57740 480904 57792
rect 480956 57780 480962 57792
rect 487062 57780 487068 57792
rect 480956 57752 487068 57780
rect 480956 57740 480962 57752
rect 487062 57740 487068 57752
rect 487120 57740 487126 57792
rect 502426 57740 502432 57792
rect 502484 57780 502490 57792
rect 508038 57780 508044 57792
rect 502484 57752 508044 57780
rect 502484 57740 502490 57752
rect 508038 57740 508044 57752
rect 508096 57740 508102 57792
rect 171962 57672 171968 57724
rect 172020 57712 172026 57724
rect 203150 57712 203156 57724
rect 172020 57684 203156 57712
rect 172020 57672 172026 57684
rect 203150 57672 203156 57684
rect 203208 57672 203214 57724
rect 214558 57672 214564 57724
rect 214616 57712 214622 57724
rect 214616 57684 217732 57712
rect 214616 57672 214622 57684
rect 175090 57604 175096 57656
rect 175148 57644 175154 57656
rect 217594 57644 217600 57656
rect 175148 57616 217600 57644
rect 175148 57604 175154 57616
rect 217594 57604 217600 57616
rect 217652 57604 217658 57656
rect 171870 57536 171876 57588
rect 171928 57576 171934 57588
rect 214742 57576 214748 57588
rect 171928 57548 214748 57576
rect 171928 57536 171934 57548
rect 214742 57536 214748 57548
rect 214800 57536 214806 57588
rect 217704 57576 217732 57684
rect 407206 57672 407212 57724
rect 407264 57712 407270 57724
rect 407758 57712 407764 57724
rect 407264 57684 407764 57712
rect 407264 57672 407270 57684
rect 407758 57672 407764 57684
rect 407816 57672 407822 57724
rect 419534 57672 419540 57724
rect 419592 57712 419598 57724
rect 420086 57712 420092 57724
rect 419592 57684 420092 57712
rect 419592 57672 419598 57684
rect 420086 57672 420092 57684
rect 420144 57672 420150 57724
rect 420914 57672 420920 57724
rect 420972 57712 420978 57724
rect 421558 57712 421564 57724
rect 420972 57684 421564 57712
rect 420972 57672 420978 57684
rect 421558 57672 421564 57684
rect 421616 57672 421622 57724
rect 423674 57672 423680 57724
rect 423732 57712 423738 57724
rect 424502 57712 424508 57724
rect 423732 57684 424508 57712
rect 423732 57672 423738 57684
rect 424502 57672 424508 57684
rect 424560 57672 424566 57724
rect 425054 57672 425060 57724
rect 425112 57712 425118 57724
rect 425974 57712 425980 57724
rect 425112 57684 425980 57712
rect 425112 57672 425118 57684
rect 425974 57672 425980 57684
rect 426032 57672 426038 57724
rect 438118 57672 438124 57724
rect 438176 57712 438182 57724
rect 439222 57712 439228 57724
rect 438176 57684 439228 57712
rect 438176 57672 438182 57684
rect 439222 57672 439228 57684
rect 439280 57672 439286 57724
rect 467098 57672 467104 57724
rect 467156 57712 467162 57724
rect 475470 57712 475476 57724
rect 467156 57684 475476 57712
rect 467156 57672 467162 57684
rect 475470 57672 475476 57684
rect 475528 57672 475534 57724
rect 478138 57672 478144 57724
rect 478196 57712 478202 57724
rect 484854 57712 484860 57724
rect 478196 57684 484860 57712
rect 478196 57672 478202 57684
rect 484854 57672 484860 57684
rect 484912 57672 484918 57724
rect 487798 57672 487804 57724
rect 487856 57712 487862 57724
rect 495710 57712 495716 57724
rect 487856 57684 495716 57712
rect 487856 57672 487862 57684
rect 495710 57672 495716 57684
rect 495768 57672 495774 57724
rect 503714 57672 503720 57724
rect 503772 57712 503778 57724
rect 508774 57712 508780 57724
rect 503772 57684 508780 57712
rect 503772 57672 503778 57684
rect 508774 57672 508780 57684
rect 508832 57672 508838 57724
rect 522574 57672 522580 57724
rect 522632 57712 522638 57724
rect 525886 57712 525892 57724
rect 522632 57684 525892 57712
rect 522632 57672 522638 57684
rect 525886 57672 525892 57684
rect 525944 57672 525950 57724
rect 541342 57672 541348 57724
rect 541400 57712 541406 57724
rect 556338 57712 556344 57724
rect 541400 57684 556344 57712
rect 541400 57672 541406 57684
rect 556338 57672 556344 57684
rect 556396 57672 556402 57724
rect 227714 57604 227720 57656
rect 227772 57644 227778 57656
rect 228174 57644 228180 57656
rect 227772 57616 228180 57644
rect 227772 57604 227778 57616
rect 228174 57604 228180 57616
rect 228232 57604 228238 57656
rect 229094 57604 229100 57656
rect 229152 57644 229158 57656
rect 229646 57644 229652 57656
rect 229152 57616 229652 57644
rect 229152 57604 229158 57616
rect 229646 57604 229652 57616
rect 229704 57604 229710 57656
rect 233234 57604 233240 57656
rect 233292 57644 233298 57656
rect 233878 57644 233884 57656
rect 233292 57616 233884 57644
rect 233292 57604 233298 57616
rect 233878 57604 233884 57616
rect 233936 57604 233942 57656
rect 237374 57604 237380 57656
rect 237432 57644 237438 57656
rect 238294 57644 238300 57656
rect 237432 57616 238300 57644
rect 237432 57604 237438 57616
rect 238294 57604 238300 57616
rect 238352 57604 238358 57656
rect 242894 57604 242900 57656
rect 242952 57644 242958 57656
rect 243446 57644 243452 57656
rect 242952 57616 243452 57644
rect 242952 57604 242958 57616
rect 243446 57604 243452 57616
rect 243504 57604 243510 57656
rect 244274 57604 244280 57656
rect 244332 57644 244338 57656
rect 244918 57644 244924 57656
rect 244332 57616 244924 57644
rect 244332 57604 244338 57616
rect 244918 57604 244924 57616
rect 244976 57604 244982 57656
rect 247034 57604 247040 57656
rect 247092 57644 247098 57656
rect 247678 57644 247684 57656
rect 247092 57616 247684 57644
rect 247092 57604 247098 57616
rect 247678 57604 247684 57616
rect 247736 57604 247742 57656
rect 250530 57604 250536 57656
rect 250588 57644 250594 57656
rect 253106 57644 253112 57656
rect 250588 57616 253112 57644
rect 250588 57604 250594 57616
rect 253106 57604 253112 57616
rect 253164 57604 253170 57656
rect 254854 57604 254860 57656
rect 254912 57644 254918 57656
rect 255314 57644 255320 57656
rect 254912 57616 255320 57644
rect 254912 57604 254918 57616
rect 255314 57604 255320 57616
rect 255372 57604 255378 57656
rect 259454 57604 259460 57656
rect 259512 57644 259518 57656
rect 260006 57644 260012 57656
rect 259512 57616 260012 57644
rect 259512 57604 259518 57616
rect 260006 57604 260012 57616
rect 260064 57604 260070 57656
rect 260834 57604 260840 57656
rect 260892 57644 260898 57656
rect 261478 57644 261484 57656
rect 260892 57616 261484 57644
rect 260892 57604 260898 57616
rect 261478 57604 261484 57616
rect 261536 57604 261542 57656
rect 276014 57604 276020 57656
rect 276072 57644 276078 57656
rect 276750 57644 276756 57656
rect 276072 57616 276756 57644
rect 276072 57604 276078 57616
rect 276750 57604 276756 57616
rect 276808 57604 276814 57656
rect 278038 57604 278044 57656
rect 278096 57644 278102 57656
rect 279234 57644 279240 57656
rect 278096 57616 279240 57644
rect 278096 57604 278102 57616
rect 279234 57604 279240 57616
rect 279292 57604 279298 57656
rect 289814 57604 289820 57656
rect 289872 57644 289878 57656
rect 290550 57644 290556 57656
rect 289872 57616 290556 57644
rect 289872 57604 289878 57616
rect 290550 57604 290556 57616
rect 290608 57604 290614 57656
rect 296714 57604 296720 57656
rect 296772 57644 296778 57656
rect 297726 57644 297732 57656
rect 296772 57616 297732 57644
rect 296772 57604 296778 57616
rect 297726 57604 297732 57616
rect 297784 57604 297790 57656
rect 302234 57604 302240 57656
rect 302292 57644 302298 57656
rect 302694 57644 302700 57656
rect 302292 57616 302700 57644
rect 302292 57604 302298 57616
rect 302694 57604 302700 57616
rect 302752 57604 302758 57656
rect 303614 57604 303620 57656
rect 303672 57644 303678 57656
rect 304166 57644 304172 57656
rect 303672 57616 304172 57644
rect 303672 57604 303678 57616
rect 304166 57604 304172 57616
rect 304224 57604 304230 57656
rect 307754 57604 307760 57656
rect 307812 57644 307818 57656
rect 308582 57644 308588 57656
rect 307812 57616 308588 57644
rect 307812 57604 307818 57616
rect 308582 57604 308588 57616
rect 308640 57604 308646 57656
rect 318794 57604 318800 57656
rect 318852 57644 318858 57656
rect 319438 57644 319444 57656
rect 318852 57616 319444 57644
rect 318852 57604 318858 57616
rect 319438 57604 319444 57616
rect 319496 57604 319502 57656
rect 320174 57604 320180 57656
rect 320232 57644 320238 57656
rect 320910 57644 320916 57656
rect 320232 57616 320916 57644
rect 320232 57604 320238 57616
rect 320910 57604 320916 57616
rect 320968 57604 320974 57656
rect 324314 57604 324320 57656
rect 324372 57644 324378 57656
rect 325142 57644 325148 57656
rect 324372 57616 325148 57644
rect 324372 57604 324378 57616
rect 325142 57604 325148 57616
rect 325200 57604 325206 57656
rect 325694 57604 325700 57656
rect 325752 57644 325758 57656
rect 326614 57644 326620 57656
rect 325752 57616 326620 57644
rect 325752 57604 325758 57616
rect 326614 57604 326620 57616
rect 326672 57604 326678 57656
rect 329834 57604 329840 57656
rect 329892 57644 329898 57656
rect 330294 57644 330300 57656
rect 329892 57616 330300 57644
rect 329892 57604 329898 57616
rect 330294 57604 330300 57616
rect 330352 57604 330358 57656
rect 331214 57604 331220 57656
rect 331272 57644 331278 57656
rect 331766 57644 331772 57656
rect 331272 57616 331772 57644
rect 331272 57604 331278 57616
rect 331766 57604 331772 57616
rect 331824 57604 331830 57656
rect 333974 57604 333980 57656
rect 334032 57644 334038 57656
rect 334710 57644 334716 57656
rect 334032 57616 334716 57644
rect 334032 57604 334038 57616
rect 334710 57604 334716 57616
rect 334768 57604 334774 57656
rect 345014 57604 345020 57656
rect 345072 57644 345078 57656
rect 345566 57644 345572 57656
rect 345072 57616 345572 57644
rect 345072 57604 345078 57616
rect 345566 57604 345572 57616
rect 345624 57604 345630 57656
rect 346486 57604 346492 57656
rect 346544 57644 346550 57656
rect 347038 57644 347044 57656
rect 346544 57616 347044 57644
rect 346544 57604 346550 57616
rect 347038 57604 347044 57616
rect 347096 57604 347102 57656
rect 349154 57604 349160 57656
rect 349212 57644 349218 57656
rect 349798 57644 349804 57656
rect 349212 57616 349804 57644
rect 349212 57604 349218 57616
rect 349798 57604 349804 57616
rect 349856 57604 349862 57656
rect 350626 57604 350632 57656
rect 350684 57644 350690 57656
rect 351270 57644 351276 57656
rect 350684 57616 351276 57644
rect 350684 57604 350690 57616
rect 351270 57604 351276 57616
rect 351328 57604 351334 57656
rect 362954 57604 362960 57656
rect 363012 57644 363018 57656
rect 363598 57644 363604 57656
rect 363012 57616 363604 57644
rect 363012 57604 363018 57616
rect 363598 57604 363604 57616
rect 363656 57604 363662 57656
rect 367094 57604 367100 57656
rect 367152 57644 367158 57656
rect 368014 57644 368020 57656
rect 367152 57616 368020 57644
rect 367152 57604 367158 57616
rect 368014 57604 368020 57616
rect 368072 57604 368078 57656
rect 373994 57604 374000 57656
rect 374052 57644 374058 57656
rect 374454 57644 374460 57656
rect 374052 57616 374460 57644
rect 374052 57604 374058 57616
rect 374454 57604 374460 57616
rect 374512 57604 374518 57656
rect 378134 57604 378140 57656
rect 378192 57644 378198 57656
rect 378870 57644 378876 57656
rect 378192 57616 378876 57644
rect 378192 57604 378198 57616
rect 378870 57604 378876 57616
rect 378928 57604 378934 57656
rect 389174 57604 389180 57656
rect 389232 57644 389238 57656
rect 389726 57644 389732 57656
rect 389232 57616 389732 57644
rect 389232 57604 389238 57616
rect 389726 57604 389732 57616
rect 389784 57604 389790 57656
rect 391934 57604 391940 57656
rect 391992 57644 391998 57656
rect 392670 57644 392676 57656
rect 391992 57616 392676 57644
rect 391992 57604 391998 57616
rect 392670 57604 392676 57616
rect 392728 57604 392734 57656
rect 393406 57604 393412 57656
rect 393464 57644 393470 57656
rect 393958 57644 393964 57656
rect 393464 57616 393964 57644
rect 393464 57604 393470 57616
rect 393958 57604 393964 57616
rect 394016 57604 394022 57656
rect 394694 57604 394700 57656
rect 394752 57644 394758 57656
rect 395430 57644 395436 57656
rect 394752 57616 395436 57644
rect 394752 57604 394758 57616
rect 395430 57604 395436 57616
rect 395488 57604 395494 57656
rect 396074 57604 396080 57656
rect 396132 57644 396138 57656
rect 396902 57644 396908 57656
rect 396132 57616 396908 57644
rect 396132 57604 396138 57616
rect 396902 57604 396908 57616
rect 396960 57604 396966 57656
rect 400214 57604 400220 57656
rect 400272 57644 400278 57656
rect 445754 57644 445760 57656
rect 400272 57616 445760 57644
rect 400272 57604 400278 57616
rect 445754 57604 445760 57616
rect 445812 57604 445818 57656
rect 446398 57604 446404 57656
rect 446456 57644 446462 57656
rect 447962 57644 447968 57656
rect 446456 57616 447968 57644
rect 446456 57604 446462 57616
rect 447962 57604 447968 57616
rect 448020 57604 448026 57656
rect 452654 57604 452660 57656
rect 452712 57644 452718 57656
rect 453390 57644 453396 57656
rect 452712 57616 453396 57644
rect 452712 57604 452718 57616
rect 453390 57604 453396 57616
rect 453448 57604 453454 57656
rect 458910 57604 458916 57656
rect 458968 57644 458974 57656
rect 460290 57644 460296 57656
rect 458968 57616 460296 57644
rect 458968 57604 458974 57616
rect 460290 57604 460296 57616
rect 460348 57604 460354 57656
rect 462314 57604 462320 57656
rect 462372 57644 462378 57656
rect 462774 57644 462780 57656
rect 462372 57616 462780 57644
rect 462372 57604 462378 57616
rect 462774 57604 462780 57616
rect 462832 57604 462838 57656
rect 463694 57604 463700 57656
rect 463752 57644 463758 57656
rect 464246 57644 464252 57656
rect 463752 57616 464252 57644
rect 463752 57604 463758 57616
rect 464246 57604 464252 57616
rect 464304 57604 464310 57656
rect 464338 57604 464344 57656
rect 464396 57644 464402 57656
rect 464396 57616 473952 57644
rect 464396 57604 464402 57616
rect 250254 57576 250260 57588
rect 217704 57548 250260 57576
rect 250254 57536 250260 57548
rect 250312 57536 250318 57588
rect 254578 57536 254584 57588
rect 254636 57576 254642 57588
rect 263226 57576 263232 57588
rect 254636 57548 263232 57576
rect 254636 57536 254642 57548
rect 263226 57536 263232 57548
rect 263284 57536 263290 57588
rect 393314 57536 393320 57588
rect 393372 57576 393378 57588
rect 441430 57576 441436 57588
rect 393372 57548 441436 57576
rect 393372 57536 393378 57548
rect 441430 57536 441436 57548
rect 441488 57536 441494 57588
rect 441614 57536 441620 57588
rect 441672 57576 441678 57588
rect 442534 57576 442540 57588
rect 441672 57548 442540 57576
rect 441672 57536 441678 57548
rect 442534 57536 442540 57548
rect 442592 57536 442598 57588
rect 458818 57536 458824 57588
rect 458876 57576 458882 57588
rect 471882 57576 471888 57588
rect 458876 57548 471888 57576
rect 458876 57536 458882 57548
rect 471882 57536 471888 57548
rect 471940 57536 471946 57588
rect 473924 57576 473952 57616
rect 473998 57604 474004 57656
rect 474056 57644 474062 57656
rect 476206 57644 476212 57656
rect 474056 57616 476212 57644
rect 474056 57604 474062 57616
rect 476206 57604 476212 57616
rect 476264 57604 476270 57656
rect 479794 57644 479800 57656
rect 476316 57616 479800 57644
rect 476316 57576 476344 57616
rect 479794 57604 479800 57616
rect 479852 57604 479858 57656
rect 486418 57604 486424 57656
rect 486476 57644 486482 57656
rect 489270 57644 489276 57656
rect 486476 57616 489276 57644
rect 486476 57604 486482 57616
rect 489270 57604 489276 57616
rect 489328 57604 489334 57656
rect 489362 57604 489368 57656
rect 489420 57644 489426 57656
rect 494974 57644 494980 57656
rect 489420 57616 494980 57644
rect 489420 57604 489426 57616
rect 494974 57604 494980 57616
rect 495032 57604 495038 57656
rect 499390 57644 499396 57656
rect 495084 57616 499396 57644
rect 473924 57548 476344 57576
rect 477494 57536 477500 57588
rect 477552 57576 477558 57588
rect 492858 57576 492864 57588
rect 477552 57548 492864 57576
rect 477552 57536 477558 57548
rect 492858 57536 492864 57548
rect 492916 57536 492922 57588
rect 177666 57468 177672 57520
rect 177724 57508 177730 57520
rect 222010 57508 222016 57520
rect 177724 57480 222016 57508
rect 177724 57468 177730 57480
rect 222010 57468 222016 57480
rect 222068 57468 222074 57520
rect 224218 57468 224224 57520
rect 224276 57508 224282 57520
rect 241514 57508 241520 57520
rect 224276 57480 241520 57508
rect 224276 57468 224282 57480
rect 241514 57468 241520 57480
rect 241572 57468 241578 57520
rect 247678 57468 247684 57520
rect 247736 57508 247742 57520
rect 273438 57508 273444 57520
rect 247736 57480 273444 57508
rect 247736 57468 247742 57480
rect 273438 57468 273444 57480
rect 273496 57468 273502 57520
rect 386414 57468 386420 57520
rect 386472 57508 386478 57520
rect 437106 57508 437112 57520
rect 386472 57480 437112 57508
rect 386472 57468 386478 57480
rect 437106 57468 437112 57480
rect 437164 57468 437170 57520
rect 467190 57468 467196 57520
rect 467248 57508 467254 57520
rect 484118 57508 484124 57520
rect 467248 57480 484124 57508
rect 467248 57468 467254 57480
rect 484118 57468 484124 57480
rect 484176 57468 484182 57520
rect 488534 57468 488540 57520
rect 488592 57508 488598 57520
rect 495084 57508 495112 57616
rect 499390 57604 499396 57616
rect 499448 57604 499454 57656
rect 505278 57604 505284 57656
rect 505336 57644 505342 57656
rect 509510 57644 509516 57656
rect 505336 57616 509516 57644
rect 505336 57604 505342 57616
rect 509510 57604 509516 57616
rect 509568 57604 509574 57656
rect 513374 57604 513380 57656
rect 513432 57644 513438 57656
rect 514294 57644 514300 57656
rect 513432 57616 514300 57644
rect 513432 57604 513438 57616
rect 514294 57604 514300 57616
rect 514352 57604 514358 57656
rect 514754 57604 514760 57656
rect 514812 57644 514818 57656
rect 515766 57644 515772 57656
rect 514812 57616 515772 57644
rect 514812 57604 514818 57616
rect 515766 57604 515772 57616
rect 515824 57604 515830 57656
rect 524414 57604 524420 57656
rect 524472 57644 524478 57656
rect 525150 57644 525156 57656
rect 524472 57616 525156 57644
rect 524472 57604 524478 57616
rect 525150 57604 525156 57616
rect 525208 57604 525214 57656
rect 534074 57604 534080 57656
rect 534132 57644 534138 57656
rect 534534 57644 534540 57656
rect 534132 57616 534540 57644
rect 534132 57604 534138 57616
rect 534534 57604 534540 57616
rect 534592 57604 534598 57656
rect 536282 57604 536288 57656
rect 536340 57644 536346 57656
rect 537478 57644 537484 57656
rect 536340 57616 537484 57644
rect 536340 57604 536346 57616
rect 537478 57604 537484 57616
rect 537536 57604 537542 57656
rect 538214 57604 538220 57656
rect 538272 57644 538278 57656
rect 538950 57644 538956 57656
rect 538272 57616 538956 57644
rect 538272 57604 538278 57616
rect 538950 57604 538956 57616
rect 539008 57604 539014 57656
rect 539594 57604 539600 57656
rect 539652 57644 539658 57656
rect 540238 57644 540244 57656
rect 539652 57616 540244 57644
rect 539652 57604 539658 57616
rect 540238 57604 540244 57616
rect 540296 57604 540302 57656
rect 543734 57604 543740 57656
rect 543792 57644 543798 57656
rect 544654 57644 544660 57656
rect 543792 57616 544660 57644
rect 543792 57604 543798 57616
rect 544654 57604 544660 57616
rect 544712 57604 544718 57656
rect 550634 57604 550640 57656
rect 550692 57644 550698 57656
rect 551278 57644 551284 57656
rect 550692 57616 551284 57644
rect 550692 57604 550698 57616
rect 551278 57604 551284 57616
rect 551336 57604 551342 57656
rect 554774 57604 554780 57656
rect 554832 57644 554838 57656
rect 555510 57644 555516 57656
rect 554832 57616 555516 57644
rect 554832 57604 554838 57616
rect 555510 57604 555516 57616
rect 555568 57604 555574 57656
rect 504450 57576 504456 57588
rect 497016 57548 504456 57576
rect 497016 57520 497044 57548
rect 504450 57536 504456 57548
rect 504508 57536 504514 57588
rect 509326 57536 509332 57588
rect 509384 57576 509390 57588
rect 512362 57576 512368 57588
rect 509384 57548 512368 57576
rect 509384 57536 509390 57548
rect 512362 57536 512368 57548
rect 512420 57536 512426 57588
rect 529750 57536 529756 57588
rect 529808 57576 529814 57588
rect 534718 57576 534724 57588
rect 529808 57548 534724 57576
rect 529808 57536 529814 57548
rect 534718 57536 534724 57548
rect 534776 57536 534782 57588
rect 552198 57536 552204 57588
rect 552256 57576 552262 57588
rect 567838 57576 567844 57588
rect 552256 57548 567844 57576
rect 552256 57536 552262 57548
rect 567838 57536 567844 57548
rect 567896 57536 567902 57588
rect 488592 57480 495112 57508
rect 488592 57468 488598 57480
rect 496998 57468 497004 57520
rect 497056 57468 497062 57520
rect 498286 57468 498292 57520
rect 498344 57508 498350 57520
rect 505922 57508 505928 57520
rect 498344 57480 505928 57508
rect 498344 57468 498350 57480
rect 505922 57468 505928 57480
rect 505980 57468 505986 57520
rect 510798 57468 510804 57520
rect 510856 57508 510862 57520
rect 513098 57508 513104 57520
rect 510856 57480 513104 57508
rect 510856 57468 510862 57480
rect 513098 57468 513104 57480
rect 513156 57468 513162 57520
rect 542814 57468 542820 57520
rect 542872 57508 542878 57520
rect 558178 57508 558184 57520
rect 542872 57480 558184 57508
rect 542872 57468 542878 57480
rect 558178 57468 558184 57480
rect 558236 57468 558242 57520
rect 170766 57400 170772 57452
rect 170824 57440 170830 57452
rect 245838 57440 245844 57452
rect 170824 57412 245844 57440
rect 170824 57400 170830 57412
rect 245838 57400 245844 57412
rect 245896 57400 245902 57452
rect 246298 57400 246304 57452
rect 246356 57440 246362 57452
rect 251634 57440 251640 57452
rect 246356 57412 251640 57440
rect 246356 57400 246362 57412
rect 251634 57400 251640 57412
rect 251692 57400 251698 57452
rect 254670 57400 254676 57452
rect 254728 57440 254734 57452
rect 284662 57440 284668 57452
rect 254728 57412 284668 57440
rect 254728 57400 254734 57412
rect 284662 57400 284668 57412
rect 284720 57400 284726 57452
rect 284938 57400 284944 57452
rect 284996 57440 285002 57452
rect 295886 57440 295892 57452
rect 284996 57412 295892 57440
rect 284996 57400 285002 57412
rect 295886 57400 295892 57412
rect 295944 57400 295950 57452
rect 377398 57400 377404 57452
rect 377456 57440 377462 57452
rect 430574 57440 430580 57452
rect 377456 57412 430580 57440
rect 377456 57400 377462 57412
rect 430574 57400 430580 57412
rect 430632 57400 430638 57452
rect 459554 57400 459560 57452
rect 459612 57440 459618 57452
rect 482002 57440 482008 57452
rect 459612 57412 482008 57440
rect 459612 57400 459618 57412
rect 482002 57400 482008 57412
rect 482060 57400 482066 57452
rect 485038 57400 485044 57452
rect 485096 57440 485102 57452
rect 489362 57440 489368 57452
rect 485096 57412 489368 57440
rect 485096 57400 485102 57412
rect 489362 57400 489368 57412
rect 489420 57400 489426 57452
rect 494054 57400 494060 57452
rect 494112 57440 494118 57452
rect 502978 57440 502984 57452
rect 494112 57412 502984 57440
rect 494112 57400 494118 57412
rect 502978 57400 502984 57412
rect 503036 57400 503042 57452
rect 535546 57400 535552 57452
rect 535604 57440 535610 57452
rect 547138 57440 547144 57452
rect 535604 57412 547144 57440
rect 535604 57400 535610 57412
rect 547138 57400 547144 57412
rect 547196 57400 547202 57452
rect 549346 57400 549352 57452
rect 549404 57440 549410 57452
rect 566458 57440 566464 57452
rect 549404 57412 566464 57440
rect 549404 57400 549410 57412
rect 566458 57400 566464 57412
rect 566516 57400 566522 57452
rect 188522 57332 188528 57384
rect 188580 57372 188586 57384
rect 269758 57372 269764 57384
rect 188580 57344 269764 57372
rect 188580 57332 188586 57344
rect 269758 57332 269764 57344
rect 269816 57332 269822 57384
rect 271138 57332 271144 57384
rect 271196 57372 271202 57384
rect 287146 57372 287152 57384
rect 271196 57344 287152 57372
rect 271196 57332 271202 57344
rect 287146 57332 287152 57344
rect 287204 57332 287210 57384
rect 287698 57332 287704 57384
rect 287756 57372 287762 57384
rect 289354 57372 289360 57384
rect 287756 57344 289360 57372
rect 287756 57332 287762 57344
rect 289354 57332 289360 57344
rect 289412 57332 289418 57384
rect 350534 57332 350540 57384
rect 350592 57372 350598 57384
rect 415394 57372 415400 57384
rect 350592 57344 415400 57372
rect 350592 57332 350598 57344
rect 415394 57332 415400 57344
rect 415452 57332 415458 57384
rect 440878 57332 440884 57384
rect 440936 57372 440942 57384
rect 440936 57344 467604 57372
rect 440936 57332 440942 57344
rect 175182 57264 175188 57316
rect 175240 57304 175246 57316
rect 258902 57304 258908 57316
rect 175240 57276 258908 57304
rect 175240 57264 175246 57276
rect 258902 57264 258908 57276
rect 258960 57264 258966 57316
rect 266998 57264 267004 57316
rect 267056 57304 267062 57316
rect 272702 57304 272708 57316
rect 267056 57276 272708 57304
rect 267056 57264 267062 57276
rect 272702 57264 272708 57276
rect 272760 57264 272766 57316
rect 273898 57264 273904 57316
rect 273956 57304 273962 57316
rect 293678 57304 293684 57316
rect 273956 57276 293684 57304
rect 273956 57264 273962 57276
rect 293678 57264 293684 57276
rect 293736 57264 293742 57316
rect 343634 57264 343640 57316
rect 343692 57304 343698 57316
rect 410978 57304 410984 57316
rect 343692 57276 410984 57304
rect 343692 57264 343698 57276
rect 410978 57264 410984 57276
rect 411036 57264 411042 57316
rect 436094 57264 436100 57316
rect 436152 57304 436158 57316
rect 467466 57304 467472 57316
rect 436152 57276 467472 57304
rect 436152 57264 436158 57276
rect 467466 57264 467472 57276
rect 467524 57264 467530 57316
rect 467576 57304 467604 57344
rect 468478 57332 468484 57384
rect 468536 57372 468542 57384
rect 468536 57344 482232 57372
rect 468536 57332 468542 57344
rect 468938 57304 468944 57316
rect 467576 57276 468944 57304
rect 468938 57264 468944 57276
rect 468996 57264 469002 57316
rect 470594 57264 470600 57316
rect 470652 57304 470658 57316
rect 482204 57304 482232 57344
rect 482278 57332 482284 57384
rect 482336 57372 482342 57384
rect 493594 57372 493600 57384
rect 482336 57344 493600 57372
rect 482336 57332 482342 57344
rect 493594 57332 493600 57344
rect 493652 57332 493658 57384
rect 500218 57332 500224 57384
rect 500276 57372 500282 57384
rect 502242 57372 502248 57384
rect 500276 57344 502248 57372
rect 500276 57332 500282 57344
rect 502242 57332 502248 57344
rect 502300 57332 502306 57384
rect 529014 57332 529020 57384
rect 529072 57372 529078 57384
rect 530578 57372 530584 57384
rect 529072 57344 530584 57372
rect 529072 57332 529078 57344
rect 530578 57332 530584 57344
rect 530636 57332 530642 57384
rect 543550 57332 543556 57384
rect 543608 57372 543614 57384
rect 560294 57372 560300 57384
rect 543608 57344 560300 57372
rect 543608 57332 543614 57344
rect 560294 57332 560300 57344
rect 560352 57332 560358 57384
rect 486326 57304 486332 57316
rect 470652 57276 482140 57304
rect 482204 57276 486332 57304
rect 470652 57264 470658 57276
rect 170858 57196 170864 57248
rect 170916 57236 170922 57248
rect 254302 57236 254308 57248
rect 170916 57208 254308 57236
rect 170916 57196 170922 57208
rect 254302 57196 254308 57208
rect 254360 57196 254366 57248
rect 258810 57196 258816 57248
rect 258868 57236 258874 57248
rect 291470 57236 291476 57248
rect 258868 57208 291476 57236
rect 258868 57196 258874 57208
rect 291470 57196 291476 57208
rect 291528 57196 291534 57248
rect 338758 57196 338764 57248
rect 338816 57236 338822 57248
rect 406654 57236 406660 57248
rect 338816 57208 406660 57236
rect 338816 57196 338822 57208
rect 406654 57196 406660 57208
rect 406712 57196 406718 57248
rect 407114 57196 407120 57248
rect 407172 57236 407178 57248
rect 450078 57236 450084 57248
rect 407172 57208 450084 57236
rect 407172 57196 407178 57208
rect 450078 57196 450084 57208
rect 450136 57196 450142 57248
rect 454678 57196 454684 57248
rect 454736 57236 454742 57248
rect 456610 57236 456616 57248
rect 454736 57208 456616 57236
rect 454736 57196 454742 57208
rect 456610 57196 456616 57208
rect 456668 57196 456674 57248
rect 456794 57196 456800 57248
rect 456852 57236 456858 57248
rect 480530 57236 480536 57248
rect 456852 57208 480536 57236
rect 456852 57196 456858 57208
rect 480530 57196 480536 57208
rect 480588 57196 480594 57248
rect 482112 57168 482140 57276
rect 486326 57264 486332 57276
rect 486384 57264 486390 57316
rect 490190 57264 490196 57316
rect 490248 57304 490254 57316
rect 500770 57304 500776 57316
rect 490248 57276 500776 57304
rect 490248 57264 490254 57276
rect 500770 57264 500776 57276
rect 500828 57264 500834 57316
rect 545758 57264 545764 57316
rect 545816 57304 545822 57316
rect 564434 57304 564440 57316
rect 545816 57276 564440 57304
rect 545816 57264 545822 57276
rect 564434 57264 564440 57276
rect 564492 57264 564498 57316
rect 484394 57196 484400 57248
rect 484452 57236 484458 57248
rect 496814 57236 496820 57248
rect 484452 57208 496820 57236
rect 484452 57196 484458 57208
rect 496814 57196 496820 57208
rect 496872 57196 496878 57248
rect 498194 57196 498200 57248
rect 498252 57236 498258 57248
rect 505186 57236 505192 57248
rect 498252 57208 505192 57236
rect 498252 57196 498258 57208
rect 505186 57196 505192 57208
rect 505244 57196 505250 57248
rect 556614 57196 556620 57248
rect 556672 57236 556678 57248
rect 582374 57236 582380 57248
rect 556672 57208 582380 57236
rect 556672 57196 556678 57208
rect 582374 57196 582380 57208
rect 582432 57196 582438 57248
rect 488626 57168 488632 57180
rect 482112 57140 488632 57168
rect 488626 57128 488632 57140
rect 488684 57128 488690 57180
rect 264238 57060 264244 57112
rect 264296 57100 264302 57112
rect 266170 57100 266176 57112
rect 264296 57072 266176 57100
rect 264296 57060 264302 57072
rect 266170 57060 266176 57072
rect 266228 57060 266234 57112
rect 518894 57060 518900 57112
rect 518952 57100 518958 57112
rect 520274 57100 520280 57112
rect 518952 57072 520280 57100
rect 518952 57060 518958 57072
rect 520274 57060 520280 57072
rect 520332 57060 520338 57112
rect 531958 57060 531964 57112
rect 532016 57100 532022 57112
rect 538858 57100 538864 57112
rect 532016 57072 538864 57100
rect 532016 57060 532022 57072
rect 538858 57060 538864 57072
rect 538916 57060 538922 57112
rect 231118 56924 231124 56976
rect 231176 56964 231182 56976
rect 232866 56964 232872 56976
rect 231176 56936 232872 56964
rect 231176 56924 231182 56936
rect 232866 56924 232872 56936
rect 232924 56924 232930 56976
rect 277394 56788 277400 56840
rect 277452 56828 277458 56840
rect 278222 56828 278228 56840
rect 277452 56800 278228 56828
rect 277452 56788 277458 56800
rect 278222 56788 278228 56800
rect 278280 56788 278286 56840
rect 523310 56788 523316 56840
rect 523368 56828 523374 56840
rect 527174 56828 527180 56840
rect 523368 56800 527180 56828
rect 523368 56788 523374 56800
rect 527174 56788 527180 56800
rect 527232 56788 527238 56840
rect 499758 56720 499764 56772
rect 499816 56760 499822 56772
rect 506566 56760 506572 56772
rect 499816 56732 506572 56760
rect 499816 56720 499822 56732
rect 506566 56720 506572 56732
rect 506624 56720 506630 56772
rect 506474 56652 506480 56704
rect 506532 56692 506538 56704
rect 510614 56692 510620 56704
rect 506532 56664 510620 56692
rect 506532 56652 506538 56664
rect 510614 56652 510620 56664
rect 510672 56652 510678 56704
rect 233878 56584 233884 56636
rect 233936 56624 233942 56636
rect 239398 56624 239404 56636
rect 233936 56596 239404 56624
rect 233936 56584 233942 56596
rect 239398 56584 239404 56596
rect 239456 56584 239462 56636
rect 410518 56584 410524 56636
rect 410576 56624 410582 56636
rect 413186 56624 413192 56636
rect 410576 56596 413192 56624
rect 410576 56584 410582 56596
rect 413186 56584 413192 56596
rect 413244 56584 413250 56636
rect 442994 56584 443000 56636
rect 443052 56624 443058 56636
rect 444006 56624 444012 56636
rect 443052 56596 444012 56624
rect 443052 56584 443058 56596
rect 444006 56584 444012 56596
rect 444064 56584 444070 56636
rect 447778 56584 447784 56636
rect 447836 56624 447842 56636
rect 452286 56624 452292 56636
rect 447836 56596 452292 56624
rect 447836 56584 447842 56596
rect 452286 56584 452292 56596
rect 452344 56584 452350 56636
rect 476758 56584 476764 56636
rect 476816 56624 476822 56636
rect 482738 56624 482744 56636
rect 476816 56596 482744 56624
rect 476816 56584 476822 56596
rect 482738 56584 482744 56596
rect 482796 56584 482802 56636
rect 508498 56584 508504 56636
rect 508556 56624 508562 56636
rect 510246 56624 510252 56636
rect 508556 56596 510252 56624
rect 508556 56584 508562 56596
rect 510246 56584 510252 56596
rect 510304 56584 510310 56636
rect 527266 56244 527272 56296
rect 527324 56284 527330 56296
rect 528094 56284 528100 56296
rect 527324 56256 528100 56284
rect 527324 56244 527330 56256
rect 528094 56244 528100 56256
rect 528152 56244 528158 56296
rect 269758 55972 269764 56024
rect 269816 56012 269822 56024
rect 362494 56012 362500 56024
rect 269816 55984 362500 56012
rect 269816 55972 269822 55984
rect 362494 55972 362500 55984
rect 362552 55972 362558 56024
rect 258718 55904 258724 55956
rect 258776 55944 258782 55956
rect 355226 55944 355232 55956
rect 258776 55916 355232 55944
rect 258776 55904 258782 55916
rect 355226 55904 355232 55916
rect 355284 55904 355290 55956
rect 364334 55904 364340 55956
rect 364392 55944 364398 55956
rect 423306 55944 423312 55956
rect 364392 55916 423312 55944
rect 364392 55904 364398 55916
rect 423306 55904 423312 55916
rect 423364 55904 423370 55956
rect 426434 55904 426440 55956
rect 426492 55944 426498 55956
rect 461670 55944 461676 55956
rect 426492 55916 461676 55944
rect 426492 55904 426498 55916
rect 461670 55904 461676 55916
rect 461728 55904 461734 55956
rect 171226 55836 171232 55888
rect 171284 55876 171290 55888
rect 305270 55876 305276 55888
rect 171284 55848 305276 55876
rect 171284 55836 171290 55848
rect 305270 55836 305276 55848
rect 305328 55836 305334 55888
rect 308398 55836 308404 55888
rect 308456 55876 308462 55888
rect 382734 55876 382740 55888
rect 308456 55848 382740 55876
rect 308456 55836 308462 55848
rect 382734 55836 382740 55848
rect 382792 55836 382798 55888
rect 383654 55836 383660 55888
rect 383712 55876 383718 55888
rect 435634 55876 435640 55888
rect 383712 55848 435640 55876
rect 383712 55836 383718 55848
rect 435634 55836 435640 55848
rect 435692 55836 435698 55888
rect 448698 55836 448704 55888
rect 448756 55876 448762 55888
rect 474734 55876 474740 55888
rect 448756 55848 474740 55876
rect 448756 55836 448762 55848
rect 474734 55836 474740 55848
rect 474792 55836 474798 55888
rect 483014 55836 483020 55888
rect 483072 55876 483078 55888
rect 496446 55876 496452 55888
rect 483072 55848 496452 55876
rect 483072 55836 483078 55848
rect 496446 55836 496452 55848
rect 496504 55836 496510 55888
rect 533430 55836 533436 55888
rect 533488 55876 533494 55888
rect 543826 55876 543832 55888
rect 533488 55848 543832 55876
rect 533488 55836 533494 55848
rect 543826 55836 543832 55848
rect 543884 55836 543890 55888
rect 546402 55836 546408 55888
rect 546460 55876 546466 55888
rect 564526 55876 564532 55888
rect 546460 55848 564532 55876
rect 546460 55836 546466 55848
rect 564526 55836 564532 55848
rect 564584 55836 564590 55888
rect 471974 55564 471980 55616
rect 472032 55604 472038 55616
rect 472894 55604 472900 55616
rect 472032 55576 472900 55604
rect 472032 55564 472038 55576
rect 472894 55564 472900 55576
rect 472952 55564 472958 55616
rect 456886 55428 456892 55480
rect 456944 55468 456950 55480
rect 457806 55468 457812 55480
rect 456944 55440 457812 55468
rect 456944 55428 456950 55440
rect 457806 55428 457812 55440
rect 457864 55428 457870 55480
rect 454034 55360 454040 55412
rect 454092 55400 454098 55412
rect 454862 55400 454868 55412
rect 454092 55372 454868 55400
rect 454092 55360 454098 55372
rect 454862 55360 454868 55372
rect 454920 55360 454926 55412
rect 346394 54680 346400 54732
rect 346452 54720 346458 54732
rect 411898 54720 411904 54732
rect 346452 54692 411904 54720
rect 346452 54680 346458 54692
rect 411898 54680 411904 54692
rect 411956 54680 411962 54732
rect 276658 54612 276664 54664
rect 276716 54652 276722 54664
rect 358998 54652 359004 54664
rect 276716 54624 359004 54652
rect 276716 54612 276722 54624
rect 358998 54612 359004 54624
rect 359056 54612 359062 54664
rect 244918 54544 244924 54596
rect 244976 54584 244982 54596
rect 349246 54584 349252 54596
rect 244976 54556 349252 54584
rect 244976 54544 244982 54556
rect 349246 54544 349252 54556
rect 349304 54544 349310 54596
rect 440234 54544 440240 54596
rect 440292 54584 440298 54596
rect 469950 54584 469956 54596
rect 440292 54556 469956 54584
rect 440292 54544 440298 54556
rect 469950 54544 469956 54556
rect 470008 54544 470014 54596
rect 487246 54544 487252 54596
rect 487304 54584 487310 54596
rect 498378 54584 498384 54596
rect 487304 54556 498384 54584
rect 487304 54544 487310 54556
rect 498378 54544 498384 54556
rect 498436 54544 498442 54596
rect 178034 54476 178040 54528
rect 178092 54516 178098 54528
rect 309134 54516 309140 54528
rect 178092 54488 309140 54516
rect 178092 54476 178098 54488
rect 309134 54476 309140 54488
rect 309192 54476 309198 54528
rect 311158 54476 311164 54528
rect 311216 54516 311222 54528
rect 389266 54516 389272 54528
rect 311216 54488 389272 54516
rect 311216 54476 311222 54488
rect 389266 54476 389272 54488
rect 389324 54476 389330 54528
rect 405734 54476 405740 54528
rect 405792 54516 405798 54528
rect 448514 54516 448520 54528
rect 405792 54488 448520 54516
rect 405792 54476 405798 54488
rect 448514 54476 448520 54488
rect 448572 54476 448578 54528
rect 476206 54476 476212 54528
rect 476264 54516 476270 54528
rect 491478 54516 491484 54528
rect 476264 54488 491484 54516
rect 476264 54476 476270 54488
rect 491478 54476 491484 54488
rect 491536 54476 491542 54528
rect 552474 54476 552480 54528
rect 552532 54516 552538 54528
rect 574738 54516 574744 54528
rect 552532 54488 574744 54516
rect 552532 54476 552538 54488
rect 574738 54476 574744 54488
rect 574796 54476 574802 54528
rect 298738 53252 298744 53304
rect 298796 53292 298802 53304
rect 381538 53292 381544 53304
rect 298796 53264 381544 53292
rect 298796 53252 298802 53264
rect 381538 53252 381544 53264
rect 381596 53252 381602 53304
rect 268378 53184 268384 53236
rect 268436 53224 268442 53236
rect 361574 53224 361580 53236
rect 268436 53196 361580 53224
rect 268436 53184 268442 53196
rect 361574 53184 361580 53196
rect 361632 53184 361638 53236
rect 226426 53116 226432 53168
rect 226484 53156 226490 53168
rect 338666 53156 338672 53168
rect 226484 53128 338672 53156
rect 226484 53116 226490 53128
rect 338666 53116 338672 53128
rect 338724 53116 338730 53168
rect 412634 53116 412640 53168
rect 412692 53156 412698 53168
rect 452746 53156 452752 53168
rect 412692 53128 452752 53156
rect 412692 53116 412698 53128
rect 452746 53116 452752 53128
rect 452804 53116 452810 53168
rect 200298 53048 200304 53100
rect 200356 53088 200362 53100
rect 322014 53088 322020 53100
rect 200356 53060 322020 53088
rect 200356 53048 200362 53060
rect 322014 53048 322020 53060
rect 322072 53048 322078 53100
rect 367186 53048 367192 53100
rect 367244 53088 367250 53100
rect 425146 53088 425152 53100
rect 367244 53060 425152 53088
rect 367244 53048 367250 53060
rect 425146 53048 425152 53060
rect 425204 53048 425210 53100
rect 444374 53048 444380 53100
rect 444432 53088 444438 53100
rect 472066 53088 472072 53100
rect 444432 53060 472072 53088
rect 444432 53048 444438 53060
rect 472066 53048 472072 53060
rect 472124 53048 472130 53100
rect 473354 53048 473360 53100
rect 473412 53088 473418 53100
rect 489914 53088 489920 53100
rect 473412 53060 489920 53088
rect 473412 53048 473418 53060
rect 489914 53048 489920 53060
rect 489972 53048 489978 53100
rect 554866 53048 554872 53100
rect 554924 53088 554930 53100
rect 578878 53088 578884 53100
rect 554924 53060 578884 53088
rect 554924 53048 554930 53060
rect 578878 53048 578884 53060
rect 578936 53048 578942 53100
rect 285030 51892 285036 51944
rect 285088 51932 285094 51944
rect 372706 51932 372712 51944
rect 285088 51904 372712 51932
rect 285088 51892 285094 51904
rect 372706 51892 372712 51904
rect 372764 51892 372770 51944
rect 266354 51824 266360 51876
rect 266412 51864 266418 51876
rect 363046 51864 363052 51876
rect 266412 51836 363052 51864
rect 266412 51824 266418 51836
rect 363046 51824 363052 51836
rect 363104 51824 363110 51876
rect 209774 51756 209780 51808
rect 209832 51796 209838 51808
rect 328546 51796 328552 51808
rect 209832 51768 328552 51796
rect 209832 51756 209838 51768
rect 328546 51756 328552 51768
rect 328604 51756 328610 51808
rect 379606 51756 379612 51808
rect 379664 51796 379670 51808
rect 432138 51796 432144 51808
rect 379664 51768 432144 51796
rect 379664 51756 379670 51768
rect 432138 51756 432144 51768
rect 432196 51756 432202 51808
rect 184934 51688 184940 51740
rect 184992 51728 184998 51740
rect 313274 51728 313280 51740
rect 184992 51700 313280 51728
rect 184992 51688 184998 51700
rect 313274 51688 313280 51700
rect 313332 51688 313338 51740
rect 360194 51688 360200 51740
rect 360252 51728 360258 51740
rect 421006 51728 421012 51740
rect 360252 51700 421012 51728
rect 360252 51688 360258 51700
rect 421006 51688 421012 51700
rect 421064 51688 421070 51740
rect 430666 51688 430672 51740
rect 430724 51728 430730 51740
rect 463786 51728 463792 51740
rect 430724 51700 463792 51728
rect 430724 51688 430730 51700
rect 463786 51688 463792 51700
rect 463844 51688 463850 51740
rect 554774 51688 554780 51740
rect 554832 51728 554838 51740
rect 580258 51728 580264 51740
rect 554832 51700 580264 51728
rect 554832 51688 554838 51700
rect 580258 51688 580264 51700
rect 580316 51688 580322 51740
rect 309134 50464 309140 50516
rect 309192 50504 309198 50516
rect 389174 50504 389180 50516
rect 309192 50476 389180 50504
rect 309192 50464 309198 50476
rect 389174 50464 389180 50476
rect 389232 50464 389238 50516
rect 238018 50396 238024 50448
rect 238076 50436 238082 50448
rect 345106 50436 345112 50448
rect 238076 50408 345112 50436
rect 238076 50396 238082 50408
rect 345106 50396 345112 50408
rect 345164 50396 345170 50448
rect 218698 50328 218704 50380
rect 218756 50368 218762 50380
rect 331306 50368 331312 50380
rect 218756 50340 331312 50368
rect 218756 50328 218762 50340
rect 331306 50328 331312 50340
rect 331364 50328 331370 50380
rect 374086 50328 374092 50380
rect 374144 50368 374150 50380
rect 429194 50368 429200 50380
rect 374144 50340 429200 50368
rect 374144 50328 374150 50340
rect 429194 50328 429200 50340
rect 429252 50328 429258 50380
rect 433426 50328 433432 50380
rect 433484 50368 433490 50380
rect 465534 50368 465540 50380
rect 433484 50340 465540 50368
rect 433484 50328 433490 50340
rect 465534 50328 465540 50340
rect 465592 50328 465598 50380
rect 330478 49172 330484 49224
rect 330536 49212 330542 49224
rect 394694 49212 394700 49224
rect 330536 49184 394700 49212
rect 330536 49172 330542 49184
rect 394694 49172 394700 49184
rect 394752 49172 394758 49224
rect 313274 49104 313280 49156
rect 313332 49144 313338 49156
rect 392026 49144 392032 49156
rect 313332 49116 392032 49144
rect 313332 49104 313338 49116
rect 392026 49104 392032 49116
rect 392084 49104 392090 49156
rect 226978 49036 226984 49088
rect 227036 49076 227042 49088
rect 333146 49076 333152 49088
rect 227036 49048 333152 49076
rect 227036 49036 227042 49048
rect 333146 49036 333152 49048
rect 333204 49036 333210 49088
rect 173526 48968 173532 49020
rect 173584 49008 173590 49020
rect 226518 49008 226524 49020
rect 173584 48980 226524 49008
rect 173584 48968 173590 48980
rect 226518 48968 226524 48980
rect 226576 48968 226582 49020
rect 233326 48968 233332 49020
rect 233384 49008 233390 49020
rect 342254 49008 342260 49020
rect 233384 48980 342260 49008
rect 233384 48968 233390 48980
rect 342254 48968 342260 48980
rect 342312 48968 342318 49020
rect 394694 48968 394700 49020
rect 394752 49008 394758 49020
rect 441706 49008 441712 49020
rect 394752 48980 441712 49008
rect 394752 48968 394758 48980
rect 441706 48968 441712 48980
rect 441764 48968 441770 49020
rect 455414 48968 455420 49020
rect 455472 49008 455478 49020
rect 478966 49008 478972 49020
rect 455472 48980 478972 49008
rect 455472 48968 455478 48980
rect 478966 48968 478972 48980
rect 479024 48968 479030 49020
rect 334618 47744 334624 47796
rect 334676 47784 334682 47796
rect 399478 47784 399484 47796
rect 334676 47756 399484 47784
rect 334676 47744 334682 47756
rect 399478 47744 399484 47756
rect 399536 47744 399542 47796
rect 257338 47676 257344 47728
rect 257396 47716 257402 47728
rect 351914 47716 351920 47728
rect 257396 47688 351920 47716
rect 257396 47676 257402 47688
rect 351914 47676 351920 47688
rect 351972 47676 351978 47728
rect 407390 47676 407396 47728
rect 407448 47716 407454 47728
rect 448606 47716 448612 47728
rect 407448 47688 448612 47716
rect 407448 47676 407454 47688
rect 448606 47676 448612 47688
rect 448664 47676 448670 47728
rect 220814 47608 220820 47660
rect 220872 47648 220878 47660
rect 335354 47648 335360 47660
rect 220872 47620 335360 47648
rect 220872 47608 220878 47620
rect 335354 47608 335360 47620
rect 335412 47608 335418 47660
rect 218238 47540 218244 47592
rect 218296 47580 218302 47592
rect 334066 47580 334072 47592
rect 218296 47552 334072 47580
rect 218296 47540 218302 47552
rect 334066 47540 334072 47552
rect 334124 47540 334130 47592
rect 339678 47540 339684 47592
rect 339736 47580 339742 47592
rect 407206 47580 407212 47592
rect 339736 47552 407212 47580
rect 339736 47540 339742 47552
rect 407206 47540 407212 47552
rect 407264 47540 407270 47592
rect 447870 47540 447876 47592
rect 447928 47580 447934 47592
rect 471974 47580 471980 47592
rect 447928 47552 471980 47580
rect 447928 47540 447934 47552
rect 471974 47540 471980 47552
rect 472032 47540 472038 47592
rect 574830 46860 574836 46912
rect 574888 46900 574894 46912
rect 580166 46900 580172 46912
rect 574888 46872 580172 46900
rect 574888 46860 574894 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 276750 46316 276756 46368
rect 276808 46356 276814 46368
rect 366174 46356 366180 46368
rect 276808 46328 366180 46356
rect 276808 46316 276814 46328
rect 366174 46316 366180 46328
rect 366232 46316 366238 46368
rect 416958 46316 416964 46368
rect 417016 46356 417022 46368
rect 455506 46356 455512 46368
rect 417016 46328 455512 46356
rect 417016 46316 417022 46328
rect 455506 46316 455512 46328
rect 455564 46316 455570 46368
rect 240778 46248 240784 46300
rect 240836 46288 240842 46300
rect 339494 46288 339500 46300
rect 240836 46260 339500 46288
rect 240836 46248 240842 46260
rect 339494 46248 339500 46260
rect 339552 46248 339558 46300
rect 179414 46180 179420 46232
rect 179472 46220 179478 46232
rect 309870 46220 309876 46232
rect 179472 46192 309876 46220
rect 179472 46180 179478 46192
rect 309870 46180 309876 46192
rect 309928 46180 309934 46232
rect 353386 46180 353392 46232
rect 353444 46220 353450 46232
rect 416866 46220 416872 46232
rect 353444 46192 416872 46220
rect 353444 46180 353450 46192
rect 416866 46180 416872 46192
rect 416924 46180 416930 46232
rect 250438 45024 250444 45076
rect 250496 45064 250502 45076
rect 340966 45064 340972 45076
rect 250496 45036 340972 45064
rect 250496 45024 250502 45036
rect 340966 45024 340972 45036
rect 341024 45024 341030 45076
rect 280154 44956 280160 45008
rect 280212 44996 280218 45008
rect 371234 44996 371240 45008
rect 280212 44968 371240 44996
rect 280212 44956 280218 44968
rect 371234 44956 371240 44968
rect 371292 44956 371298 45008
rect 191834 44888 191840 44940
rect 191892 44928 191898 44940
rect 317414 44928 317420 44940
rect 191892 44900 317420 44928
rect 191892 44888 191898 44900
rect 317414 44888 317420 44900
rect 317472 44888 317478 44940
rect 450538 44888 450544 44940
rect 450596 44928 450602 44940
rect 473446 44928 473452 44940
rect 450596 44900 473452 44928
rect 450596 44888 450602 44900
rect 473446 44888 473452 44900
rect 473504 44888 473510 44940
rect 172514 44820 172520 44872
rect 172572 44860 172578 44872
rect 304994 44860 305000 44872
rect 172572 44832 305000 44860
rect 172572 44820 172578 44832
rect 304994 44820 305000 44832
rect 305052 44820 305058 44872
rect 340966 44820 340972 44872
rect 341024 44860 341030 44872
rect 408586 44860 408592 44872
rect 341024 44832 408592 44860
rect 341024 44820 341030 44832
rect 408586 44820 408592 44832
rect 408644 44820 408650 44872
rect 409874 44820 409880 44872
rect 409932 44860 409938 44872
rect 451366 44860 451372 44872
rect 409932 44832 451372 44860
rect 409932 44820 409938 44832
rect 451366 44820 451372 44832
rect 451424 44820 451430 44872
rect 317414 43596 317420 43648
rect 317472 43636 317478 43648
rect 394786 43636 394792 43648
rect 317472 43608 394792 43636
rect 317472 43596 317478 43608
rect 394786 43596 394792 43608
rect 394844 43596 394850 43648
rect 236638 43528 236644 43580
rect 236696 43568 236702 43580
rect 343818 43568 343824 43580
rect 236696 43540 343824 43568
rect 236696 43528 236702 43540
rect 343818 43528 343824 43540
rect 343876 43528 343882 43580
rect 216766 43460 216772 43512
rect 216824 43500 216830 43512
rect 332594 43500 332600 43512
rect 216824 43472 332600 43500
rect 216824 43460 216830 43472
rect 332594 43460 332600 43472
rect 332652 43460 332658 43512
rect 193214 43392 193220 43444
rect 193272 43432 193278 43444
rect 318886 43432 318892 43444
rect 193272 43404 318892 43432
rect 193272 43392 193278 43404
rect 318886 43392 318892 43404
rect 318944 43392 318950 43444
rect 348418 43392 348424 43444
rect 348476 43432 348482 43444
rect 401686 43432 401692 43444
rect 348476 43404 401692 43432
rect 348476 43392 348482 43404
rect 401686 43392 401692 43404
rect 401744 43392 401750 43444
rect 414106 43392 414112 43444
rect 414164 43432 414170 43444
rect 452654 43432 452660 43444
rect 414164 43404 452660 43432
rect 414164 43392 414170 43404
rect 452654 43392 452660 43404
rect 452712 43392 452718 43444
rect 287146 42236 287152 42288
rect 287204 42276 287210 42288
rect 375466 42276 375472 42288
rect 287204 42248 375472 42276
rect 287204 42236 287210 42248
rect 375466 42236 375472 42248
rect 375524 42236 375530 42288
rect 247770 42168 247776 42220
rect 247828 42208 247834 42220
rect 347866 42208 347872 42220
rect 247828 42180 347872 42208
rect 247828 42168 247834 42180
rect 347866 42168 347872 42180
rect 347924 42168 347930 42220
rect 194594 42100 194600 42152
rect 194652 42140 194658 42152
rect 318794 42140 318800 42152
rect 194652 42112 318800 42140
rect 194652 42100 194658 42112
rect 318794 42100 318800 42112
rect 318852 42100 318858 42152
rect 176654 42032 176660 42084
rect 176712 42072 176718 42084
rect 307846 42072 307852 42084
rect 176712 42044 307852 42072
rect 176712 42032 176718 42044
rect 307846 42032 307852 42044
rect 307904 42032 307910 42084
rect 351914 42032 351920 42084
rect 351972 42072 351978 42084
rect 415486 42072 415492 42084
rect 351972 42044 415492 42072
rect 351972 42032 351978 42044
rect 415486 42032 415492 42044
rect 415544 42032 415550 42084
rect 427998 42032 428004 42084
rect 428056 42072 428062 42084
rect 462406 42072 462412 42084
rect 428056 42044 462412 42072
rect 428056 42032 428062 42044
rect 462406 42032 462412 42044
rect 462464 42032 462470 42084
rect 304258 40876 304264 40928
rect 304316 40916 304322 40928
rect 378226 40916 378232 40928
rect 304316 40888 378232 40916
rect 304316 40876 304322 40888
rect 378226 40876 378232 40888
rect 378284 40876 378290 40928
rect 245746 40808 245752 40860
rect 245804 40848 245810 40860
rect 350718 40848 350724 40860
rect 245804 40820 350724 40848
rect 245804 40808 245810 40820
rect 350718 40808 350724 40820
rect 350776 40808 350782 40860
rect 198734 40740 198740 40792
rect 198792 40780 198798 40792
rect 321554 40780 321560 40792
rect 198792 40752 321560 40780
rect 198792 40740 198798 40752
rect 321554 40740 321560 40752
rect 321612 40740 321618 40792
rect 183554 40672 183560 40724
rect 183612 40712 183618 40724
rect 311894 40712 311900 40724
rect 183612 40684 311900 40712
rect 183612 40672 183618 40684
rect 311894 40672 311900 40684
rect 311952 40672 311958 40724
rect 342254 40672 342260 40724
rect 342312 40712 342318 40724
rect 409966 40712 409972 40724
rect 342312 40684 409972 40712
rect 342312 40672 342318 40684
rect 409966 40672 409972 40684
rect 410024 40672 410030 40724
rect 240870 39448 240876 39500
rect 240928 39488 240934 39500
rect 346578 39488 346584 39500
rect 240928 39460 346584 39488
rect 240928 39448 240934 39460
rect 346578 39448 346584 39460
rect 346636 39448 346642 39500
rect 205726 39380 205732 39432
rect 205784 39420 205790 39432
rect 325786 39420 325792 39432
rect 205784 39392 325792 39420
rect 205784 39380 205790 39392
rect 325786 39380 325792 39392
rect 325844 39380 325850 39432
rect 327718 39380 327724 39432
rect 327776 39420 327782 39432
rect 393498 39420 393504 39432
rect 327776 39392 393504 39420
rect 327776 39380 327782 39392
rect 393498 39380 393504 39392
rect 393556 39380 393562 39432
rect 397638 39380 397644 39432
rect 397696 39420 397702 39432
rect 443086 39420 443092 39432
rect 397696 39392 443092 39420
rect 397696 39380 397702 39392
rect 443086 39380 443092 39392
rect 443144 39380 443150 39432
rect 186314 39312 186320 39364
rect 186372 39352 186378 39364
rect 314746 39352 314752 39364
rect 186372 39324 314752 39352
rect 186372 39312 186378 39324
rect 314746 39312 314752 39324
rect 314804 39312 314810 39364
rect 335354 39312 335360 39364
rect 335412 39352 335418 39364
rect 405826 39352 405832 39364
rect 335412 39324 405832 39352
rect 335412 39312 335418 39324
rect 405826 39312 405832 39324
rect 405884 39312 405890 39364
rect 297358 38020 297364 38072
rect 297416 38060 297422 38072
rect 380894 38060 380900 38072
rect 297416 38032 380900 38060
rect 297416 38020 297422 38032
rect 380894 38020 380900 38032
rect 380952 38020 380958 38072
rect 259638 37952 259644 38004
rect 259696 37992 259702 38004
rect 358814 37992 358820 38004
rect 259696 37964 358820 37992
rect 259696 37952 259702 37964
rect 358814 37952 358820 37964
rect 358872 37952 358878 38004
rect 231210 37884 231216 37936
rect 231268 37924 231274 37936
rect 339586 37924 339592 37936
rect 231268 37896 339592 37924
rect 231268 37884 231274 37896
rect 339586 37884 339592 37896
rect 339644 37884 339650 37936
rect 356698 37884 356704 37936
rect 356756 37924 356762 37936
rect 408494 37924 408500 37936
rect 356756 37896 408500 37924
rect 356756 37884 356762 37896
rect 408494 37884 408500 37896
rect 408552 37884 408558 37936
rect 289906 36660 289912 36712
rect 289964 36700 289970 36712
rect 376846 36700 376852 36712
rect 289964 36672 376852 36700
rect 289964 36660 289970 36672
rect 376846 36660 376852 36672
rect 376904 36660 376910 36712
rect 254762 36592 254768 36644
rect 254820 36632 254826 36644
rect 352006 36632 352012 36644
rect 254820 36604 352012 36632
rect 254820 36592 254826 36604
rect 352006 36592 352012 36604
rect 352064 36592 352070 36644
rect 209958 36524 209964 36576
rect 210016 36564 210022 36576
rect 328454 36564 328460 36576
rect 210016 36536 328460 36564
rect 210016 36524 210022 36536
rect 328454 36524 328460 36536
rect 328512 36524 328518 36576
rect 378226 36524 378232 36576
rect 378284 36564 378290 36576
rect 431954 36564 431960 36576
rect 378284 36536 431960 36564
rect 378284 36524 378290 36536
rect 431954 36524 431960 36536
rect 432012 36524 432018 36576
rect 316678 35368 316684 35420
rect 316736 35408 316742 35420
rect 383838 35408 383844 35420
rect 316736 35380 383844 35408
rect 316736 35368 316742 35380
rect 383838 35368 383844 35380
rect 383896 35368 383902 35420
rect 236730 35300 236736 35352
rect 236788 35340 236794 35352
rect 336826 35340 336832 35352
rect 236788 35312 336832 35340
rect 236788 35300 236794 35312
rect 336826 35300 336832 35312
rect 336884 35300 336890 35352
rect 201678 35232 201684 35284
rect 201736 35272 201742 35284
rect 323026 35272 323032 35284
rect 201736 35244 323032 35272
rect 201736 35232 201742 35244
rect 323026 35232 323032 35244
rect 323084 35232 323090 35284
rect 384298 35232 384304 35284
rect 384356 35272 384362 35284
rect 434714 35272 434720 35284
rect 384356 35244 434720 35272
rect 384356 35232 384362 35244
rect 434714 35232 434720 35244
rect 434772 35232 434778 35284
rect 190454 35164 190460 35216
rect 190512 35204 190518 35216
rect 316218 35204 316224 35216
rect 190512 35176 316224 35204
rect 190512 35164 190518 35176
rect 316218 35164 316224 35176
rect 316276 35164 316282 35216
rect 332594 35164 332600 35216
rect 332652 35204 332658 35216
rect 403158 35204 403164 35216
rect 332652 35176 403164 35204
rect 332652 35164 332658 35176
rect 403158 35164 403164 35176
rect 403216 35164 403222 35216
rect 250622 33872 250628 33924
rect 250680 33912 250686 33924
rect 347774 33912 347780 33924
rect 250680 33884 347780 33912
rect 250680 33872 250686 33884
rect 347774 33872 347780 33884
rect 347832 33872 347838 33924
rect 172146 33804 172152 33856
rect 172204 33844 172210 33856
rect 212626 33844 212632 33856
rect 172204 33816 212632 33844
rect 172204 33804 172210 33816
rect 212626 33804 212632 33816
rect 212684 33804 212690 33856
rect 217318 33804 217324 33856
rect 217376 33844 217382 33856
rect 331214 33844 331220 33856
rect 217376 33816 331220 33844
rect 217376 33804 217382 33816
rect 331214 33804 331220 33816
rect 331272 33804 331278 33856
rect 365806 33804 365812 33856
rect 365864 33844 365870 33856
rect 423766 33844 423772 33856
rect 365864 33816 423772 33844
rect 365864 33804 365870 33816
rect 423766 33804 423772 33816
rect 423824 33804 423830 33856
rect 207198 33736 207204 33788
rect 207256 33776 207262 33788
rect 325694 33776 325700 33788
rect 207256 33748 325700 33776
rect 207256 33736 207262 33748
rect 325694 33736 325700 33748
rect 325752 33736 325758 33788
rect 328454 33736 328460 33788
rect 328512 33776 328518 33788
rect 401594 33776 401600 33788
rect 328512 33748 401600 33776
rect 328512 33736 328518 33748
rect 401594 33736 401600 33748
rect 401652 33736 401658 33788
rect 320358 32580 320364 32632
rect 320416 32620 320422 32632
rect 396166 32620 396172 32632
rect 320416 32592 396172 32620
rect 320416 32580 320422 32592
rect 396166 32580 396172 32592
rect 396224 32580 396230 32632
rect 264330 32512 264336 32564
rect 264388 32552 264394 32564
rect 356054 32552 356060 32564
rect 264388 32524 356060 32552
rect 264388 32512 264394 32524
rect 356054 32512 356060 32524
rect 356112 32512 356118 32564
rect 228358 32444 228364 32496
rect 228416 32484 228422 32496
rect 338114 32484 338120 32496
rect 228416 32456 338120 32484
rect 228416 32444 228422 32456
rect 338114 32444 338120 32456
rect 338172 32444 338178 32496
rect 195974 32376 195980 32428
rect 196032 32416 196038 32428
rect 320266 32416 320272 32428
rect 196032 32388 320272 32416
rect 196032 32376 196038 32388
rect 320266 32376 320272 32388
rect 320324 32376 320330 32428
rect 396166 32376 396172 32428
rect 396224 32416 396230 32428
rect 441614 32416 441620 32428
rect 396224 32388 441620 32416
rect 396224 32376 396230 32388
rect 441614 32376 441620 32388
rect 441672 32376 441678 32428
rect 169386 31220 169392 31272
rect 169444 31260 169450 31272
rect 276106 31260 276112 31272
rect 169444 31232 276112 31260
rect 169444 31220 169450 31232
rect 276106 31220 276112 31232
rect 276164 31220 276170 31272
rect 283006 31220 283012 31272
rect 283064 31260 283070 31272
rect 372798 31260 372804 31272
rect 283064 31232 372804 31260
rect 283064 31220 283070 31232
rect 372798 31220 372804 31232
rect 372856 31220 372862 31272
rect 208578 31152 208584 31204
rect 208636 31192 208642 31204
rect 327074 31192 327080 31204
rect 208636 31164 327080 31192
rect 208636 31152 208642 31164
rect 327074 31152 327080 31164
rect 327132 31152 327138 31204
rect 189074 31084 189080 31136
rect 189132 31124 189138 31136
rect 316034 31124 316040 31136
rect 189132 31096 316040 31124
rect 189132 31084 189138 31096
rect 316034 31084 316040 31096
rect 316092 31084 316098 31136
rect 382366 31084 382372 31136
rect 382424 31124 382430 31136
rect 433518 31124 433524 31136
rect 382424 31096 433524 31124
rect 382424 31084 382430 31096
rect 433518 31084 433524 31096
rect 433576 31084 433582 31136
rect 168374 31016 168380 31068
rect 168432 31056 168438 31068
rect 303706 31056 303712 31068
rect 168432 31028 303712 31056
rect 168432 31016 168438 31028
rect 303706 31016 303712 31028
rect 303764 31016 303770 31068
rect 318058 31016 318064 31068
rect 318116 31056 318122 31068
rect 386598 31056 386604 31068
rect 318116 31028 386604 31056
rect 318116 31016 318122 31028
rect 386598 31016 386604 31028
rect 386656 31016 386662 31068
rect 433978 31016 433984 31068
rect 434036 31056 434042 31068
rect 465074 31056 465080 31068
rect 434036 31028 465080 31056
rect 434036 31016 434042 31028
rect 465074 31016 465080 31028
rect 465132 31016 465138 31068
rect 143166 29860 143172 29912
rect 143224 29900 143230 29912
rect 198182 29900 198188 29912
rect 143224 29872 198188 29900
rect 143224 29860 143230 29872
rect 198182 29860 198188 29872
rect 198240 29860 198246 29912
rect 135806 29792 135812 29844
rect 135864 29832 135870 29844
rect 198090 29832 198096 29844
rect 135864 29804 198096 29832
rect 135864 29792 135870 29804
rect 198090 29792 198096 29804
rect 198148 29792 198154 29844
rect 128354 29724 128360 29776
rect 128412 29764 128418 29776
rect 198550 29764 198556 29776
rect 128412 29736 198556 29764
rect 128412 29724 128418 29736
rect 198550 29724 198556 29736
rect 198608 29724 198614 29776
rect 237558 29724 237564 29776
rect 237616 29764 237622 29776
rect 345014 29764 345020 29776
rect 237616 29736 345020 29764
rect 237616 29724 237622 29736
rect 345014 29724 345020 29736
rect 345072 29724 345078 29776
rect 127618 29656 127624 29708
rect 127676 29696 127682 29708
rect 198366 29696 198372 29708
rect 127676 29668 198372 29696
rect 127676 29656 127682 29668
rect 198366 29656 198372 29668
rect 198424 29656 198430 29708
rect 211246 29656 211252 29708
rect 211304 29696 211310 29708
rect 329926 29696 329932 29708
rect 211304 29668 329932 29696
rect 211304 29656 211310 29668
rect 329926 29656 329932 29668
rect 329984 29656 329990 29708
rect 370498 29656 370504 29708
rect 370556 29696 370562 29708
rect 425054 29696 425060 29708
rect 370556 29668 425060 29696
rect 370556 29656 370562 29668
rect 425054 29656 425060 29668
rect 425112 29656 425118 29708
rect 124030 29588 124036 29640
rect 124088 29628 124094 29640
rect 198274 29628 198280 29640
rect 124088 29600 198280 29628
rect 124088 29588 124094 29600
rect 198274 29588 198280 29600
rect 198332 29588 198338 29640
rect 204898 29588 204904 29640
rect 204956 29628 204962 29640
rect 324406 29628 324412 29640
rect 204956 29600 324412 29628
rect 204956 29588 204962 29600
rect 324406 29588 324412 29600
rect 324464 29588 324470 29640
rect 331214 29588 331220 29640
rect 331272 29628 331278 29640
rect 402974 29628 402980 29640
rect 331272 29600 402980 29628
rect 331272 29588 331278 29600
rect 402974 29588 402980 29600
rect 403032 29588 403038 29640
rect 429194 29588 429200 29640
rect 429252 29628 429258 29640
rect 462314 29628 462320 29640
rect 429252 29600 462320 29628
rect 429252 29588 429258 29600
rect 462314 29588 462320 29600
rect 462372 29588 462378 29640
rect 166166 29520 166172 29572
rect 166224 29560 166230 29572
rect 198642 29560 198648 29572
rect 166224 29532 198648 29560
rect 166224 29520 166230 29532
rect 198642 29520 198648 29532
rect 198700 29520 198706 29572
rect 166258 29452 166264 29504
rect 166316 29492 166322 29504
rect 198458 29492 198464 29504
rect 166316 29464 198464 29492
rect 166316 29452 166322 29464
rect 198458 29452 198464 29464
rect 198516 29452 198522 29504
rect 166350 29384 166356 29436
rect 166408 29424 166414 29436
rect 197998 29424 198004 29436
rect 166408 29396 198004 29424
rect 166408 29384 166414 29396
rect 197998 29384 198004 29396
rect 198056 29384 198062 29436
rect 130562 29044 130568 29096
rect 130620 29084 130626 29096
rect 170950 29084 170956 29096
rect 130620 29056 170956 29084
rect 130620 29044 130626 29056
rect 170950 29044 170956 29056
rect 171008 29044 171014 29096
rect 138934 28976 138940 29028
rect 138992 29016 138998 29028
rect 188430 29016 188436 29028
rect 138992 28988 188436 29016
rect 138992 28976 138998 28988
rect 188430 28976 188436 28988
rect 188488 28976 188494 29028
rect 134242 28908 134248 28960
rect 134300 28948 134306 28960
rect 186958 28948 186964 28960
rect 134300 28920 186964 28948
rect 134300 28908 134306 28920
rect 186958 28908 186964 28920
rect 187016 28908 187022 28960
rect 143258 28840 143264 28892
rect 143316 28880 143322 28892
rect 197906 28880 197912 28892
rect 143316 28852 197912 28880
rect 143316 28840 143322 28852
rect 197906 28840 197912 28852
rect 197964 28840 197970 28892
rect 103146 28772 103152 28824
rect 103204 28812 103210 28824
rect 168190 28812 168196 28824
rect 103204 28784 168196 28812
rect 103204 28772 103210 28784
rect 168190 28772 168196 28784
rect 168248 28772 168254 28824
rect 90726 28704 90732 28756
rect 90784 28744 90790 28756
rect 168006 28744 168012 28756
rect 90784 28716 168012 28744
rect 90784 28704 90790 28716
rect 168006 28704 168012 28716
rect 168064 28704 168070 28756
rect 88058 28636 88064 28688
rect 88116 28676 88122 28688
rect 169018 28676 169024 28688
rect 88116 28648 169024 28676
rect 88116 28636 88122 28648
rect 169018 28636 169024 28648
rect 169076 28636 169082 28688
rect 83090 28568 83096 28620
rect 83148 28608 83154 28620
rect 174814 28608 174820 28620
rect 83148 28580 174820 28608
rect 83148 28568 83154 28580
rect 174814 28568 174820 28580
rect 174872 28568 174878 28620
rect 80698 28500 80704 28552
rect 80756 28540 80762 28552
rect 176194 28540 176200 28552
rect 80756 28512 176200 28540
rect 80756 28500 80762 28512
rect 176194 28500 176200 28512
rect 176252 28500 176258 28552
rect 78122 28432 78128 28484
rect 78180 28472 78186 28484
rect 177758 28472 177764 28484
rect 78180 28444 177764 28472
rect 78180 28432 78186 28444
rect 177758 28432 177764 28444
rect 177816 28432 177822 28484
rect 75546 28364 75552 28416
rect 75604 28404 75610 28416
rect 176102 28404 176108 28416
rect 75604 28376 176108 28404
rect 75604 28364 75610 28376
rect 176102 28364 176108 28376
rect 176160 28364 176166 28416
rect 60642 28296 60648 28348
rect 60700 28336 60706 28348
rect 167822 28336 167828 28348
rect 60700 28308 167828 28336
rect 60700 28296 60706 28308
rect 167822 28296 167828 28308
rect 167880 28296 167886 28348
rect 244458 28296 244464 28348
rect 244516 28336 244522 28348
rect 349154 28336 349160 28348
rect 244516 28308 349160 28336
rect 244516 28296 244522 28308
rect 349154 28296 349160 28308
rect 349212 28296 349218 28348
rect 68186 28228 68192 28280
rect 68244 28268 68250 28280
rect 178954 28268 178960 28280
rect 68244 28240 178960 28268
rect 68244 28228 68250 28240
rect 178954 28228 178960 28240
rect 179012 28228 179018 28280
rect 224310 28228 224316 28280
rect 224368 28268 224374 28280
rect 335446 28268 335452 28280
rect 224368 28240 335452 28268
rect 224368 28228 224374 28240
rect 335446 28228 335452 28240
rect 335504 28228 335510 28280
rect 389174 28228 389180 28280
rect 389232 28268 389238 28280
rect 437566 28268 437572 28280
rect 389232 28240 437572 28268
rect 389232 28228 389238 28240
rect 437566 28228 437572 28240
rect 437624 28228 437630 28280
rect 128538 28160 128544 28212
rect 128596 28200 128602 28212
rect 174722 28200 174728 28212
rect 128596 28172 174728 28200
rect 128596 28160 128602 28172
rect 174722 28160 174728 28172
rect 174780 28160 174786 28212
rect 135898 28092 135904 28144
rect 135956 28132 135962 28144
rect 172054 28132 172060 28144
rect 135956 28104 172060 28132
rect 135956 28092 135962 28104
rect 172054 28092 172060 28104
rect 172112 28092 172118 28144
rect 138290 28024 138296 28076
rect 138348 28064 138354 28076
rect 169294 28064 169300 28076
rect 138348 28036 169300 28064
rect 138348 28024 138354 28036
rect 169294 28024 169300 28036
rect 169352 28024 169358 28076
rect 28626 27548 28632 27600
rect 28684 27588 28690 27600
rect 42794 27588 42800 27600
rect 28684 27560 42800 27588
rect 28684 27548 28690 27560
rect 42794 27548 42800 27560
rect 42852 27548 42858 27600
rect 120626 27548 120632 27600
rect 120684 27588 120690 27600
rect 127618 27588 127624 27600
rect 120684 27560 127624 27588
rect 120684 27548 120690 27560
rect 127618 27548 127624 27560
rect 127676 27548 127682 27600
rect 132770 27548 132776 27600
rect 132828 27588 132834 27600
rect 143258 27588 143264 27600
rect 132828 27560 143264 27588
rect 132828 27548 132834 27560
rect 143258 27548 143264 27560
rect 143316 27548 143322 27600
rect 150618 27548 150624 27600
rect 150676 27588 150682 27600
rect 167086 27588 167092 27600
rect 150676 27560 167092 27588
rect 150676 27548 150682 27560
rect 167086 27548 167092 27560
rect 167144 27548 167150 27600
rect 28810 27480 28816 27532
rect 28868 27520 28874 27532
rect 43622 27520 43628 27532
rect 28868 27492 43628 27520
rect 28868 27480 28874 27492
rect 43622 27480 43628 27492
rect 43680 27480 43686 27532
rect 143442 27480 143448 27532
rect 143500 27520 143506 27532
rect 176010 27520 176016 27532
rect 143500 27492 176016 27520
rect 143500 27480 143506 27492
rect 176010 27480 176016 27492
rect 176068 27480 176074 27532
rect 118418 27412 118424 27464
rect 118476 27452 118482 27464
rect 118476 27424 127664 27452
rect 118476 27412 118482 27424
rect 115658 27344 115664 27396
rect 115716 27384 115722 27396
rect 124030 27384 124036 27396
rect 115716 27356 124036 27384
rect 115716 27344 115722 27356
rect 124030 27344 124036 27356
rect 124088 27344 124094 27396
rect 127636 27384 127664 27424
rect 132034 27412 132040 27464
rect 132092 27452 132098 27464
rect 178862 27452 178868 27464
rect 132092 27424 178868 27452
rect 132092 27412 132098 27424
rect 178862 27412 178868 27424
rect 178920 27412 178926 27464
rect 176286 27384 176292 27396
rect 127636 27356 176292 27384
rect 176286 27344 176292 27356
rect 176344 27344 176350 27396
rect 124122 27276 124128 27328
rect 124180 27316 124186 27328
rect 180150 27316 180156 27328
rect 124180 27288 180156 27316
rect 124180 27276 124186 27288
rect 180150 27276 180156 27288
rect 180208 27276 180214 27328
rect 129642 27208 129648 27260
rect 129700 27248 129706 27260
rect 184290 27248 184296 27260
rect 129700 27220 184296 27248
rect 129700 27208 129706 27220
rect 184290 27208 184296 27220
rect 184348 27208 184354 27260
rect 126330 27140 126336 27192
rect 126388 27180 126394 27192
rect 177390 27180 177396 27192
rect 126388 27152 177396 27180
rect 126388 27140 126394 27152
rect 177390 27140 177396 27152
rect 177448 27140 177454 27192
rect 123754 27072 123760 27124
rect 123812 27112 123818 27124
rect 166258 27112 166264 27124
rect 123812 27084 166264 27112
rect 123812 27072 123818 27084
rect 166258 27072 166264 27084
rect 166316 27072 166322 27124
rect 128170 27004 128176 27056
rect 128228 27044 128234 27056
rect 166166 27044 166172 27056
rect 128228 27016 166172 27044
rect 128228 27004 128234 27016
rect 166166 27004 166172 27016
rect 166224 27004 166230 27056
rect 214742 27004 214748 27056
rect 214800 27044 214806 27056
rect 329834 27044 329840 27056
rect 214800 27016 329840 27044
rect 214800 27004 214806 27016
rect 329834 27004 329840 27016
rect 329892 27004 329898 27056
rect 112162 26936 112168 26988
rect 112220 26976 112226 26988
rect 149054 26976 149060 26988
rect 112220 26948 149060 26976
rect 112220 26936 112226 26948
rect 149054 26936 149060 26948
rect 149112 26936 149118 26988
rect 150066 26936 150072 26988
rect 150124 26976 150130 26988
rect 166994 26976 167000 26988
rect 150124 26948 167000 26976
rect 150124 26936 150130 26948
rect 166994 26936 167000 26948
rect 167052 26936 167058 26988
rect 204438 26936 204444 26988
rect 204496 26976 204502 26988
rect 324314 26976 324320 26988
rect 204496 26948 324320 26976
rect 204496 26936 204502 26948
rect 324314 26936 324320 26948
rect 324372 26936 324378 26988
rect 324958 26936 324964 26988
rect 325016 26976 325022 26988
rect 390646 26976 390652 26988
rect 325016 26948 390652 26976
rect 325016 26936 325022 26948
rect 390646 26936 390652 26948
rect 390704 26936 390710 26988
rect 110322 26868 110328 26920
rect 110380 26908 110386 26920
rect 143350 26908 143356 26920
rect 110380 26880 143356 26908
rect 110380 26868 110386 26880
rect 143350 26868 143356 26880
rect 143408 26868 143414 26920
rect 143442 26868 143448 26920
rect 143500 26908 143506 26920
rect 175918 26908 175924 26920
rect 143500 26880 175924 26908
rect 143500 26868 143506 26880
rect 175918 26868 175924 26880
rect 175976 26868 175982 26920
rect 193306 26868 193312 26920
rect 193364 26908 193370 26920
rect 317506 26908 317512 26920
rect 193364 26880 317512 26908
rect 193364 26868 193370 26880
rect 317506 26868 317512 26880
rect 317564 26868 317570 26920
rect 327074 26868 327080 26920
rect 327132 26908 327138 26920
rect 400306 26908 400312 26920
rect 327132 26880 400312 26908
rect 327132 26868 327138 26880
rect 400306 26868 400312 26880
rect 400364 26868 400370 26920
rect 418338 26868 418344 26920
rect 418396 26908 418402 26920
rect 454678 26908 454684 26920
rect 418396 26880 454684 26908
rect 418396 26868 418402 26880
rect 454678 26868 454684 26880
rect 454736 26868 454742 26920
rect 64874 26800 64880 26852
rect 64932 26840 64938 26852
rect 135806 26840 135812 26852
rect 64932 26812 135812 26840
rect 64932 26800 64938 26812
rect 135806 26800 135812 26812
rect 135864 26800 135870 26852
rect 140130 26800 140136 26852
rect 140188 26840 140194 26852
rect 167638 26840 167644 26852
rect 140188 26812 167644 26840
rect 140188 26800 140194 26812
rect 167638 26800 167644 26812
rect 167696 26800 167702 26852
rect 141234 26732 141240 26784
rect 141292 26772 141298 26784
rect 167730 26772 167736 26784
rect 141292 26744 167736 26772
rect 141292 26732 141298 26744
rect 167730 26732 167736 26744
rect 167788 26732 167794 26784
rect 63218 26664 63224 26716
rect 63276 26704 63282 26716
rect 166350 26704 166356 26716
rect 63276 26676 166356 26704
rect 63276 26664 63282 26676
rect 166350 26664 166356 26676
rect 166408 26664 166414 26716
rect 71590 26596 71596 26648
rect 71648 26636 71654 26648
rect 143166 26636 143172 26648
rect 71648 26608 143172 26636
rect 71648 26596 71654 26608
rect 143166 26596 143172 26608
rect 143224 26596 143230 26648
rect 98270 26188 98276 26240
rect 98328 26228 98334 26240
rect 174998 26228 175004 26240
rect 98328 26200 175004 26228
rect 98328 26188 98334 26200
rect 174998 26188 175004 26200
rect 175056 26188 175062 26240
rect 100202 26120 100208 26172
rect 100260 26160 100266 26172
rect 169110 26160 169116 26172
rect 100260 26132 169116 26160
rect 100260 26120 100266 26132
rect 169110 26120 169116 26132
rect 169168 26120 169174 26172
rect 105538 26052 105544 26104
rect 105596 26092 105602 26104
rect 171778 26092 171784 26104
rect 105596 26064 171784 26092
rect 105596 26052 105602 26064
rect 171778 26052 171784 26064
rect 171836 26052 171842 26104
rect 142154 25984 142160 26036
rect 142212 26024 142218 26036
rect 271138 26024 271144 26036
rect 142212 25996 271144 26024
rect 142212 25984 142218 25996
rect 271138 25984 271144 25996
rect 271196 25984 271202 26036
rect 157334 25916 157340 25968
rect 157392 25956 157398 25968
rect 295426 25956 295432 25968
rect 157392 25928 295432 25956
rect 157392 25916 157398 25928
rect 295426 25916 295432 25928
rect 295484 25916 295490 25968
rect 154574 25848 154580 25900
rect 154632 25888 154638 25900
rect 294046 25888 294052 25900
rect 154632 25860 294052 25888
rect 154632 25848 154638 25860
rect 294046 25848 294052 25860
rect 294104 25848 294110 25900
rect 128354 25780 128360 25832
rect 128412 25820 128418 25832
rect 278038 25820 278044 25832
rect 128412 25792 278044 25820
rect 128412 25780 128418 25792
rect 278038 25780 278044 25792
rect 278096 25780 278102 25832
rect 114554 25712 114560 25764
rect 114612 25752 114618 25764
rect 270586 25752 270592 25764
rect 114612 25724 270592 25752
rect 114612 25712 114618 25724
rect 270586 25712 270592 25724
rect 270644 25712 270650 25764
rect 104894 25644 104900 25696
rect 104952 25684 104958 25696
rect 263686 25684 263692 25696
rect 104952 25656 263692 25684
rect 104952 25644 104958 25656
rect 263686 25644 263692 25656
rect 263744 25644 263750 25696
rect 60734 25576 60740 25628
rect 60792 25616 60798 25628
rect 236086 25616 236092 25628
rect 60792 25588 236092 25616
rect 60792 25576 60798 25588
rect 236086 25576 236092 25588
rect 236144 25576 236150 25628
rect 294598 25576 294604 25628
rect 294656 25616 294662 25628
rect 364518 25616 364524 25628
rect 294656 25588 364524 25616
rect 294656 25576 294662 25588
rect 364518 25576 364524 25588
rect 364576 25576 364582 25628
rect 60826 25508 60832 25560
rect 60884 25548 60890 25560
rect 237466 25548 237472 25560
rect 60884 25520 237472 25548
rect 60884 25508 60890 25520
rect 237466 25508 237472 25520
rect 237524 25508 237530 25560
rect 271230 25508 271236 25560
rect 271288 25548 271294 25560
rect 362954 25548 362960 25560
rect 271288 25520 362960 25548
rect 271288 25508 271294 25520
rect 362954 25508 362960 25520
rect 363012 25508 363018 25560
rect 363046 25508 363052 25560
rect 363104 25548 363110 25560
rect 422294 25548 422300 25560
rect 363104 25520 422300 25548
rect 363104 25508 363110 25520
rect 422294 25508 422300 25520
rect 422352 25508 422358 25560
rect 431954 25508 431960 25560
rect 432012 25548 432018 25560
rect 463694 25548 463700 25560
rect 432012 25520 463700 25548
rect 432012 25508 432018 25520
rect 463694 25508 463700 25520
rect 463752 25508 463758 25560
rect 111518 25440 111524 25492
rect 111576 25480 111582 25492
rect 169202 25480 169208 25492
rect 111576 25452 169208 25480
rect 111576 25440 111582 25452
rect 169202 25440 169208 25452
rect 169260 25440 169266 25492
rect 112898 25372 112904 25424
rect 112956 25412 112962 25424
rect 173434 25412 173440 25424
rect 112956 25384 173440 25412
rect 112956 25372 112962 25384
rect 173434 25372 173440 25384
rect 173492 25372 173498 25424
rect 108022 25304 108028 25356
rect 108080 25344 108086 25356
rect 168098 25344 168104 25356
rect 108080 25316 168104 25344
rect 108080 25304 108086 25316
rect 168098 25304 168104 25316
rect 168156 25304 168162 25356
rect 147674 24760 147680 24812
rect 147732 24800 147738 24812
rect 171134 24800 171140 24812
rect 147732 24772 171140 24800
rect 147732 24760 147738 24772
rect 171134 24760 171140 24772
rect 171192 24760 171198 24812
rect 86586 24692 86592 24744
rect 86644 24732 86650 24744
rect 173158 24732 173164 24744
rect 86644 24704 173164 24732
rect 86644 24692 86650 24704
rect 173158 24692 173164 24704
rect 173216 24692 173222 24744
rect 92750 24624 92756 24676
rect 92808 24664 92814 24676
rect 174906 24664 174912 24676
rect 92808 24636 174912 24664
rect 92808 24624 92814 24636
rect 174906 24624 174912 24636
rect 174964 24624 174970 24676
rect 162854 24556 162860 24608
rect 162912 24596 162918 24608
rect 299566 24596 299572 24608
rect 162912 24568 299572 24596
rect 162912 24556 162918 24568
rect 299566 24556 299572 24568
rect 299624 24556 299630 24608
rect 146294 24488 146300 24540
rect 146352 24528 146358 24540
rect 289998 24528 290004 24540
rect 146352 24500 290004 24528
rect 146352 24488 146358 24500
rect 289998 24488 290004 24500
rect 290056 24488 290062 24540
rect 140774 24420 140780 24472
rect 140832 24460 140838 24472
rect 285766 24460 285772 24472
rect 140832 24432 285772 24460
rect 140832 24420 140838 24432
rect 285766 24420 285772 24432
rect 285824 24420 285830 24472
rect 111794 24352 111800 24404
rect 111852 24392 111858 24404
rect 267826 24392 267832 24404
rect 111852 24364 267832 24392
rect 111852 24352 111858 24364
rect 267826 24352 267832 24364
rect 267884 24352 267890 24404
rect 89714 24284 89720 24336
rect 89772 24324 89778 24336
rect 254854 24324 254860 24336
rect 89772 24296 254860 24324
rect 89772 24284 89778 24296
rect 254854 24284 254860 24296
rect 254912 24284 254918 24336
rect 85574 24216 85580 24268
rect 85632 24256 85638 24268
rect 251266 24256 251272 24268
rect 85632 24228 251272 24256
rect 85632 24216 85638 24228
rect 251266 24216 251272 24228
rect 251324 24216 251330 24268
rect 46934 24148 46940 24200
rect 46992 24188 46998 24200
rect 229186 24188 229192 24200
rect 46992 24160 229192 24188
rect 46992 24148 46998 24160
rect 229186 24148 229192 24160
rect 229244 24148 229250 24200
rect 10318 24080 10324 24132
rect 10376 24120 10382 24132
rect 204346 24120 204352 24132
rect 10376 24092 204352 24120
rect 10376 24080 10382 24092
rect 204346 24080 204352 24092
rect 204404 24080 204410 24132
rect 290458 24080 290464 24132
rect 290516 24120 290522 24132
rect 360378 24120 360384 24132
rect 290516 24092 360384 24120
rect 290516 24080 290522 24092
rect 360378 24080 360384 24092
rect 360436 24080 360442 24132
rect 392026 24080 392032 24132
rect 392084 24120 392090 24132
rect 440326 24120 440332 24132
rect 392084 24092 440332 24120
rect 392084 24080 392090 24092
rect 440326 24080 440332 24092
rect 440384 24080 440390 24132
rect 454218 24080 454224 24132
rect 454276 24120 454282 24132
rect 477586 24120 477592 24132
rect 454276 24092 477592 24120
rect 454276 24080 454282 24092
rect 477586 24080 477592 24092
rect 477644 24080 477650 24132
rect 135346 24012 135352 24064
rect 135404 24052 135410 24064
rect 177574 24052 177580 24064
rect 135404 24024 177580 24052
rect 135404 24012 135410 24024
rect 177574 24012 177580 24024
rect 177632 24012 177638 24064
rect 73982 23944 73988 23996
rect 74040 23984 74046 23996
rect 167914 23984 167920 23996
rect 74040 23956 167920 23984
rect 74040 23944 74046 23956
rect 167914 23944 167920 23956
rect 167972 23944 167978 23996
rect 95234 23876 95240 23928
rect 95292 23916 95298 23928
rect 173250 23916 173256 23928
rect 95292 23888 173256 23916
rect 95292 23876 95298 23888
rect 173250 23876 173256 23888
rect 173308 23876 173314 23928
rect 106274 23400 106280 23452
rect 106332 23440 106338 23452
rect 185578 23440 185584 23452
rect 106332 23412 185584 23440
rect 106332 23400 106338 23412
rect 185578 23400 185584 23412
rect 185636 23400 185642 23452
rect 88334 23332 88340 23384
rect 88392 23372 88398 23384
rect 170858 23372 170864 23384
rect 88392 23344 170864 23372
rect 88392 23332 88398 23344
rect 170858 23332 170864 23344
rect 170916 23332 170922 23384
rect 165614 23264 165620 23316
rect 165672 23304 165678 23316
rect 301038 23304 301044 23316
rect 165672 23276 301044 23304
rect 165672 23264 165678 23276
rect 301038 23264 301044 23276
rect 301096 23264 301102 23316
rect 166994 23196 167000 23248
rect 167052 23236 167058 23248
rect 302326 23236 302332 23248
rect 167052 23208 302332 23236
rect 167052 23196 167058 23208
rect 302326 23196 302332 23208
rect 302384 23196 302390 23248
rect 164234 23128 164240 23180
rect 164292 23168 164298 23180
rect 300854 23168 300860 23180
rect 164292 23140 300860 23168
rect 164292 23128 164298 23140
rect 300854 23128 300860 23140
rect 300912 23128 300918 23180
rect 139394 23060 139400 23112
rect 139452 23100 139458 23112
rect 285674 23100 285680 23112
rect 139452 23072 285680 23100
rect 139452 23060 139458 23072
rect 285674 23060 285680 23072
rect 285732 23060 285738 23112
rect 107654 22992 107660 23044
rect 107712 23032 107718 23044
rect 264238 23032 264244 23044
rect 107712 23004 264244 23032
rect 107712 22992 107718 23004
rect 264238 22992 264244 23004
rect 264296 22992 264302 23044
rect 69014 22924 69020 22976
rect 69072 22964 69078 22976
rect 242986 22964 242992 22976
rect 69072 22936 242992 22964
rect 69072 22924 69078 22936
rect 242986 22924 242992 22936
rect 243044 22924 243050 22976
rect 53834 22856 53840 22908
rect 53892 22896 53898 22908
rect 233418 22896 233424 22908
rect 53892 22868 233424 22896
rect 53892 22856 53898 22868
rect 233418 22856 233424 22868
rect 233476 22856 233482 22908
rect 37274 22788 37280 22840
rect 37332 22828 37338 22840
rect 222286 22828 222292 22840
rect 37332 22800 222292 22828
rect 37332 22788 37338 22800
rect 222286 22788 222292 22800
rect 222344 22788 222350 22840
rect 306558 22788 306564 22840
rect 306616 22828 306622 22840
rect 387886 22828 387892 22840
rect 306616 22800 387892 22828
rect 306616 22788 306622 22800
rect 387886 22788 387892 22800
rect 387944 22788 387950 22840
rect 2774 22720 2780 22772
rect 2832 22760 2838 22772
rect 201586 22760 201592 22772
rect 2832 22732 201592 22760
rect 2832 22720 2838 22732
rect 201586 22720 201592 22732
rect 201644 22720 201650 22772
rect 286318 22720 286324 22772
rect 286376 22760 286382 22772
rect 368566 22760 368572 22772
rect 286376 22732 368572 22760
rect 286376 22720 286382 22732
rect 368566 22720 368572 22732
rect 368624 22720 368630 22772
rect 385126 22720 385132 22772
rect 385184 22760 385190 22772
rect 436186 22760 436192 22772
rect 385184 22732 436192 22760
rect 385184 22720 385190 22732
rect 436186 22720 436192 22732
rect 436244 22720 436250 22772
rect 440326 22720 440332 22772
rect 440384 22760 440390 22772
rect 469214 22760 469220 22772
rect 440384 22732 469220 22760
rect 440384 22720 440390 22732
rect 469214 22720 469220 22732
rect 469272 22720 469278 22772
rect 118234 22652 118240 22704
rect 118292 22692 118298 22704
rect 195238 22692 195244 22704
rect 118292 22664 195244 22692
rect 118292 22652 118298 22664
rect 195238 22652 195244 22664
rect 195296 22652 195302 22704
rect 110966 22584 110972 22636
rect 111024 22624 111030 22636
rect 180058 22624 180064 22636
rect 111024 22596 180064 22624
rect 111024 22584 111030 22596
rect 180058 22584 180064 22596
rect 180116 22584 180122 22636
rect 120810 22516 120816 22568
rect 120868 22556 120874 22568
rect 173342 22556 173348 22568
rect 120868 22528 173348 22556
rect 120868 22516 120874 22528
rect 173342 22516 173348 22528
rect 173400 22516 173406 22568
rect 108758 22040 108764 22092
rect 108816 22080 108822 22092
rect 182818 22080 182824 22092
rect 108816 22052 182824 22080
rect 108816 22040 108822 22052
rect 182818 22040 182824 22052
rect 182876 22040 182882 22092
rect 120074 21972 120080 22024
rect 120132 22012 120138 22024
rect 191098 22012 191104 22024
rect 120132 21984 191104 22012
rect 120132 21972 120138 21984
rect 191098 21972 191104 21984
rect 191156 21972 191162 22024
rect 149054 21904 149060 21956
rect 149112 21944 149118 21956
rect 258810 21944 258816 21956
rect 149112 21916 258816 21944
rect 149112 21904 149118 21916
rect 258810 21904 258816 21916
rect 258868 21904 258874 21956
rect 158714 21836 158720 21888
rect 158772 21876 158778 21888
rect 296806 21876 296812 21888
rect 158772 21848 296812 21876
rect 158772 21836 158778 21848
rect 296806 21836 296812 21848
rect 296864 21836 296870 21888
rect 132494 21768 132500 21820
rect 132552 21808 132558 21820
rect 280338 21808 280344 21820
rect 132552 21780 280344 21808
rect 132552 21768 132558 21780
rect 280338 21768 280344 21780
rect 280396 21768 280402 21820
rect 126974 21700 126980 21752
rect 127032 21740 127038 21752
rect 277486 21740 277492 21752
rect 127032 21712 277492 21740
rect 127032 21700 127038 21712
rect 277486 21700 277492 21712
rect 277544 21700 277550 21752
rect 4154 21632 4160 21684
rect 4212 21672 4218 21684
rect 171962 21672 171968 21684
rect 4212 21644 171968 21672
rect 4212 21632 4218 21644
rect 171962 21632 171968 21644
rect 172020 21632 172026 21684
rect 185026 21632 185032 21684
rect 185084 21672 185090 21684
rect 313366 21672 313372 21684
rect 185084 21644 313372 21672
rect 185084 21632 185090 21644
rect 313366 21632 313372 21644
rect 313424 21632 313430 21684
rect 62114 21564 62120 21616
rect 62172 21604 62178 21616
rect 237374 21604 237380 21616
rect 62172 21576 237380 21604
rect 62172 21564 62178 21576
rect 237374 21564 237380 21576
rect 237432 21564 237438 21616
rect 57974 21496 57980 21548
rect 58032 21536 58038 21548
rect 234706 21536 234712 21548
rect 58032 21508 234712 21536
rect 58032 21496 58038 21508
rect 234706 21496 234712 21508
rect 234764 21496 234770 21548
rect 360838 21496 360844 21548
rect 360896 21536 360902 21548
rect 419626 21536 419632 21548
rect 360896 21508 419632 21536
rect 360896 21496 360902 21508
rect 419626 21496 419632 21508
rect 419684 21496 419690 21548
rect 34514 21428 34520 21480
rect 34572 21468 34578 21480
rect 220906 21468 220912 21480
rect 34572 21440 220912 21468
rect 34572 21428 34578 21440
rect 220906 21428 220912 21440
rect 220964 21428 220970 21480
rect 316034 21428 316040 21480
rect 316092 21468 316098 21480
rect 393406 21468 393412 21480
rect 316092 21440 393412 21468
rect 316092 21428 316098 21440
rect 393406 21428 393412 21440
rect 393464 21428 393470 21480
rect 16574 21360 16580 21412
rect 16632 21400 16638 21412
rect 209866 21400 209872 21412
rect 16632 21372 209872 21400
rect 16632 21360 16638 21372
rect 209866 21360 209872 21372
rect 209924 21360 209930 21412
rect 278038 21360 278044 21412
rect 278096 21400 278102 21412
rect 368474 21400 368480 21412
rect 278096 21372 368480 21400
rect 278096 21360 278102 21372
rect 368474 21360 368480 21372
rect 368532 21360 368538 21412
rect 415394 21360 415400 21412
rect 415452 21400 415458 21412
rect 454126 21400 454132 21412
rect 415452 21372 454132 21400
rect 415452 21360 415458 21372
rect 454126 21360 454132 21372
rect 454184 21360 454190 21412
rect 117130 21292 117136 21344
rect 117188 21332 117194 21344
rect 174538 21332 174544 21344
rect 117188 21304 174544 21332
rect 117188 21292 117194 21304
rect 174538 21292 174544 21304
rect 174596 21292 174602 21344
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 184198 20652 184204 20664
rect 3476 20624 184204 20652
rect 3476 20612 3482 20624
rect 184198 20612 184204 20624
rect 184256 20612 184262 20664
rect 577498 20612 577504 20664
rect 577556 20652 577562 20664
rect 579614 20652 579620 20664
rect 577556 20624 579620 20652
rect 577556 20612 577562 20624
rect 579614 20612 579620 20624
rect 579672 20612 579678 20664
rect 138014 20476 138020 20528
rect 138072 20516 138078 20528
rect 254670 20516 254676 20528
rect 138072 20488 254676 20516
rect 138072 20476 138078 20488
rect 254670 20476 254676 20488
rect 254728 20476 254734 20528
rect 182174 20408 182180 20460
rect 182232 20448 182238 20460
rect 310606 20448 310612 20460
rect 182232 20420 310612 20448
rect 182232 20408 182238 20420
rect 310606 20408 310612 20420
rect 310664 20408 310670 20460
rect 150434 20340 150440 20392
rect 150492 20380 150498 20392
rect 291286 20380 291292 20392
rect 150492 20352 291292 20380
rect 150492 20340 150498 20352
rect 291286 20340 291292 20352
rect 291344 20340 291350 20392
rect 147674 20272 147680 20324
rect 147732 20312 147738 20324
rect 289814 20312 289820 20324
rect 147732 20284 289820 20312
rect 147732 20272 147738 20284
rect 289814 20272 289820 20284
rect 289872 20272 289878 20324
rect 96614 20204 96620 20256
rect 96672 20244 96678 20256
rect 259546 20244 259552 20256
rect 96672 20216 259552 20244
rect 96672 20204 96678 20216
rect 259546 20204 259552 20216
rect 259604 20204 259610 20256
rect 38654 20136 38660 20188
rect 38712 20176 38718 20188
rect 214650 20176 214656 20188
rect 38712 20148 214656 20176
rect 38712 20136 38718 20148
rect 214650 20136 214656 20148
rect 214708 20136 214714 20188
rect 51074 20068 51080 20120
rect 51132 20108 51138 20120
rect 230566 20108 230572 20120
rect 51132 20080 230572 20108
rect 51132 20068 51138 20080
rect 230566 20068 230572 20080
rect 230624 20068 230630 20120
rect 48314 20000 48320 20052
rect 48372 20040 48378 20052
rect 229094 20040 229100 20052
rect 48372 20012 229100 20040
rect 48372 20000 48378 20012
rect 229094 20000 229100 20012
rect 229152 20000 229158 20052
rect 324314 20000 324320 20052
rect 324372 20040 324378 20052
rect 397546 20040 397552 20052
rect 324372 20012 397552 20040
rect 324372 20000 324378 20012
rect 397546 20000 397552 20012
rect 397604 20000 397610 20052
rect 22094 19932 22100 19984
rect 22152 19972 22158 19984
rect 214006 19972 214012 19984
rect 22152 19944 214012 19972
rect 22152 19932 22158 19944
rect 214006 19932 214012 19944
rect 214064 19932 214070 19984
rect 253934 19932 253940 19984
rect 253992 19972 253998 19984
rect 354674 19972 354680 19984
rect 253992 19944 354680 19972
rect 253992 19932 253998 19944
rect 354674 19932 354680 19944
rect 354732 19932 354738 19984
rect 402974 19932 402980 19984
rect 403032 19972 403038 19984
rect 447226 19972 447232 19984
rect 403032 19944 447232 19972
rect 403032 19932 403038 19944
rect 447226 19932 447232 19944
rect 447284 19932 447290 19984
rect 151814 19116 151820 19168
rect 151872 19156 151878 19168
rect 273898 19156 273904 19168
rect 151872 19128 273904 19156
rect 151872 19116 151878 19128
rect 273898 19116 273904 19128
rect 273956 19116 273962 19168
rect 161474 19048 161480 19100
rect 161532 19088 161538 19100
rect 299474 19088 299480 19100
rect 161532 19060 299480 19088
rect 161532 19048 161538 19060
rect 299474 19048 299480 19060
rect 299532 19048 299538 19100
rect 135254 18980 135260 19032
rect 135312 19020 135318 19032
rect 282914 19020 282920 19032
rect 135312 18992 282920 19020
rect 135312 18980 135318 18992
rect 282914 18980 282920 18992
rect 282972 18980 282978 19032
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 171870 18952 171876 18964
rect 23532 18924 171876 18952
rect 23532 18912 23538 18924
rect 171870 18912 171876 18924
rect 171928 18912 171934 18964
rect 175274 18912 175280 18964
rect 175332 18952 175338 18964
rect 306466 18952 306472 18964
rect 175332 18924 306472 18952
rect 175332 18912 175338 18924
rect 306466 18912 306472 18924
rect 306524 18912 306530 18964
rect 127066 18844 127072 18896
rect 127124 18884 127130 18896
rect 277394 18884 277400 18896
rect 127124 18856 277400 18884
rect 127124 18844 127130 18856
rect 277394 18844 277400 18856
rect 277452 18844 277458 18896
rect 84194 18776 84200 18828
rect 84252 18816 84258 18828
rect 246298 18816 246304 18828
rect 84252 18788 246304 18816
rect 84252 18776 84258 18788
rect 246298 18776 246304 18788
rect 246356 18776 246362 18828
rect 69106 18708 69112 18760
rect 69164 18748 69170 18760
rect 241606 18748 241612 18760
rect 69164 18720 241612 18748
rect 69164 18708 69170 18720
rect 241606 18708 241612 18720
rect 241664 18708 241670 18760
rect 357618 18708 357624 18760
rect 357676 18748 357682 18760
rect 418430 18748 418436 18760
rect 357676 18720 418436 18748
rect 357676 18708 357682 18720
rect 418430 18708 418436 18720
rect 418488 18708 418494 18760
rect 44174 18640 44180 18692
rect 44232 18680 44238 18692
rect 227806 18680 227812 18692
rect 44232 18652 227812 18680
rect 44232 18640 44238 18652
rect 227806 18640 227812 18652
rect 227864 18640 227870 18692
rect 302326 18640 302332 18692
rect 302384 18680 302390 18692
rect 385034 18680 385040 18692
rect 302384 18652 385040 18680
rect 302384 18640 302390 18652
rect 385034 18640 385040 18652
rect 385092 18640 385098 18692
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 215386 18612 215392 18624
rect 26292 18584 215392 18612
rect 26292 18572 26298 18584
rect 215386 18572 215392 18584
rect 215444 18572 215450 18624
rect 273346 18572 273352 18624
rect 273404 18612 273410 18624
rect 367278 18612 367284 18624
rect 273404 18584 367284 18612
rect 273404 18572 273410 18584
rect 367278 18572 367284 18584
rect 367336 18572 367342 18624
rect 423766 18572 423772 18624
rect 423824 18612 423830 18624
rect 458910 18612 458916 18624
rect 423824 18584 458916 18612
rect 423824 18572 423830 18584
rect 458910 18572 458916 18584
rect 458968 18572 458974 18624
rect 530026 18572 530032 18624
rect 530084 18612 530090 18624
rect 539778 18612 539784 18624
rect 530084 18584 539784 18612
rect 530084 18572 530090 18584
rect 539778 18572 539784 18584
rect 539836 18572 539842 18624
rect 118694 17756 118700 17808
rect 118752 17796 118758 17808
rect 247678 17796 247684 17808
rect 118752 17768 247684 17796
rect 118752 17756 118758 17768
rect 247678 17756 247684 17768
rect 247736 17756 247742 17808
rect 160186 17688 160192 17740
rect 160244 17728 160250 17740
rect 296714 17728 296720 17740
rect 160244 17700 296720 17728
rect 160244 17688 160250 17700
rect 296714 17688 296720 17700
rect 296772 17688 296778 17740
rect 160094 17620 160100 17672
rect 160152 17660 160158 17672
rect 298094 17660 298100 17672
rect 160152 17632 298100 17660
rect 160152 17620 160158 17632
rect 298094 17620 298100 17632
rect 298152 17620 298158 17672
rect 143534 17552 143540 17604
rect 143592 17592 143598 17604
rect 287238 17592 287244 17604
rect 143592 17564 287244 17592
rect 143592 17552 143598 17564
rect 287238 17552 287244 17564
rect 287296 17552 287302 17604
rect 136634 17484 136640 17536
rect 136692 17524 136698 17536
rect 284294 17524 284300 17536
rect 136692 17496 284300 17524
rect 136692 17484 136698 17496
rect 284294 17484 284300 17496
rect 284352 17484 284358 17536
rect 131114 17416 131120 17468
rect 131172 17456 131178 17468
rect 280246 17456 280252 17468
rect 131172 17428 280252 17456
rect 131172 17416 131178 17428
rect 280246 17416 280252 17428
rect 280304 17416 280310 17468
rect 67634 17348 67640 17400
rect 67692 17388 67698 17400
rect 224218 17388 224224 17400
rect 67692 17360 224224 17388
rect 67692 17348 67698 17360
rect 224218 17348 224224 17360
rect 224276 17348 224282 17400
rect 93854 17280 93860 17332
rect 93912 17320 93918 17332
rect 256878 17320 256884 17332
rect 93912 17292 256884 17320
rect 93912 17280 93918 17292
rect 256878 17280 256884 17292
rect 256936 17280 256942 17332
rect 299474 17280 299480 17332
rect 299532 17320 299538 17332
rect 382274 17320 382280 17332
rect 299532 17292 382280 17320
rect 299532 17280 299538 17292
rect 382274 17280 382280 17292
rect 382332 17280 382338 17332
rect 422294 17280 422300 17332
rect 422352 17320 422358 17332
rect 458174 17320 458180 17332
rect 422352 17292 458180 17320
rect 422352 17280 422358 17292
rect 458174 17280 458180 17292
rect 458232 17280 458238 17332
rect 33134 17212 33140 17264
rect 33192 17252 33198 17264
rect 219526 17252 219532 17264
rect 33192 17224 219532 17252
rect 33192 17212 33198 17224
rect 219526 17212 219532 17224
rect 219584 17212 219590 17264
rect 280798 17212 280804 17264
rect 280856 17252 280862 17264
rect 369946 17252 369952 17264
rect 280856 17224 369952 17252
rect 280856 17212 280862 17224
rect 369946 17212 369952 17224
rect 370004 17212 370010 17264
rect 371234 17212 371240 17264
rect 371292 17252 371298 17264
rect 426618 17252 426624 17264
rect 371292 17224 426624 17252
rect 371292 17212 371298 17224
rect 426618 17212 426624 17224
rect 426676 17212 426682 17264
rect 153746 16396 153752 16448
rect 153804 16436 153810 16448
rect 293954 16436 293960 16448
rect 153804 16408 293960 16436
rect 153804 16396 153810 16408
rect 293954 16396 293960 16408
rect 294012 16396 294018 16448
rect 144730 16328 144736 16380
rect 144788 16368 144794 16380
rect 288526 16368 288532 16380
rect 144788 16340 288532 16368
rect 144788 16328 144794 16340
rect 288526 16328 288532 16340
rect 288584 16328 288590 16380
rect 135346 16260 135352 16312
rect 135404 16300 135410 16312
rect 281626 16300 281632 16312
rect 135404 16272 281632 16300
rect 135404 16260 135410 16272
rect 281626 16260 281632 16272
rect 281684 16260 281690 16312
rect 125594 16192 125600 16244
rect 125652 16232 125658 16244
rect 276014 16232 276020 16244
rect 125652 16204 276020 16232
rect 125652 16192 125658 16204
rect 276014 16192 276020 16204
rect 276072 16192 276078 16244
rect 102134 16124 102140 16176
rect 102192 16164 102198 16176
rect 254578 16164 254584 16176
rect 102192 16136 254584 16164
rect 102192 16124 102198 16136
rect 254578 16124 254584 16136
rect 254636 16124 254642 16176
rect 116394 16056 116400 16108
rect 116452 16096 116458 16108
rect 270678 16096 270684 16108
rect 116452 16068 270684 16096
rect 116452 16056 116458 16068
rect 270678 16056 270684 16068
rect 270736 16056 270742 16108
rect 86402 15988 86408 16040
rect 86460 16028 86466 16040
rect 250530 16028 250536 16040
rect 86460 16000 250536 16028
rect 86460 15988 86466 16000
rect 250530 15988 250536 16000
rect 250588 15988 250594 16040
rect 334618 15988 334624 16040
rect 334676 16028 334682 16040
rect 404538 16028 404544 16040
rect 334676 16000 404544 16028
rect 334676 15988 334682 16000
rect 404538 15988 404544 16000
rect 404596 15988 404602 16040
rect 40218 15920 40224 15972
rect 40276 15960 40282 15972
rect 223666 15960 223672 15972
rect 40276 15932 223672 15960
rect 40276 15920 40282 15932
rect 223666 15920 223672 15932
rect 223724 15920 223730 15972
rect 294506 15920 294512 15972
rect 294564 15960 294570 15972
rect 379698 15960 379704 15972
rect 294564 15932 379704 15960
rect 294564 15920 294570 15932
rect 379698 15920 379704 15932
rect 379756 15920 379762 15972
rect 7650 15852 7656 15904
rect 7708 15892 7714 15904
rect 204254 15892 204260 15904
rect 7708 15864 204260 15892
rect 7708 15852 7714 15864
rect 204254 15852 204260 15864
rect 204312 15852 204318 15904
rect 270770 15852 270776 15904
rect 270828 15892 270834 15904
rect 365714 15892 365720 15904
rect 270828 15864 365720 15892
rect 270828 15852 270834 15864
rect 365714 15852 365720 15864
rect 365772 15852 365778 15904
rect 398926 15852 398932 15904
rect 398984 15892 398990 15904
rect 444466 15892 444472 15904
rect 398984 15864 444472 15892
rect 398984 15852 398990 15864
rect 444466 15852 444472 15864
rect 444524 15852 444530 15904
rect 120626 14900 120632 14952
rect 120684 14940 120690 14952
rect 273530 14940 273536 14952
rect 120684 14912 273536 14940
rect 120684 14900 120690 14912
rect 273530 14900 273536 14912
rect 273588 14900 273594 14952
rect 117314 14832 117320 14884
rect 117372 14872 117378 14884
rect 271966 14872 271972 14884
rect 117372 14844 271972 14872
rect 117372 14832 117378 14844
rect 271966 14832 271972 14844
rect 272024 14832 272030 14884
rect 110506 14764 110512 14816
rect 110564 14804 110570 14816
rect 266538 14804 266544 14816
rect 110564 14776 266544 14804
rect 110564 14764 110570 14776
rect 266538 14764 266544 14776
rect 266596 14764 266602 14816
rect 106458 14696 106464 14748
rect 106516 14736 106522 14748
rect 265066 14736 265072 14748
rect 106516 14708 265072 14736
rect 106516 14696 106522 14708
rect 265066 14696 265072 14708
rect 265124 14696 265130 14748
rect 99834 14628 99840 14680
rect 99892 14668 99898 14680
rect 260926 14668 260932 14680
rect 99892 14640 260932 14668
rect 99892 14628 99898 14640
rect 260926 14628 260932 14640
rect 260984 14628 260990 14680
rect 92474 14560 92480 14612
rect 92532 14600 92538 14612
rect 256694 14600 256700 14612
rect 92532 14572 256700 14600
rect 92532 14560 92538 14572
rect 256694 14560 256700 14572
rect 256752 14560 256758 14612
rect 338666 14560 338672 14612
rect 338724 14600 338730 14612
rect 407298 14600 407304 14612
rect 338724 14572 407304 14600
rect 338724 14560 338730 14572
rect 407298 14560 407304 14572
rect 407356 14560 407362 14612
rect 46658 14492 46664 14544
rect 46716 14532 46722 14544
rect 227714 14532 227720 14544
rect 46716 14504 227720 14532
rect 46716 14492 46722 14504
rect 227714 14492 227720 14504
rect 227772 14492 227778 14544
rect 273898 14492 273904 14544
rect 273956 14532 273962 14544
rect 353478 14532 353484 14544
rect 273956 14504 353484 14532
rect 273956 14492 273962 14504
rect 353478 14492 353484 14504
rect 353536 14492 353542 14544
rect 25314 14424 25320 14476
rect 25372 14464 25378 14476
rect 215294 14464 215300 14476
rect 25372 14436 215300 14464
rect 25372 14424 25378 14436
rect 215294 14424 215300 14436
rect 215352 14424 215358 14476
rect 277946 14424 277952 14476
rect 278004 14464 278010 14476
rect 369854 14464 369860 14476
rect 278004 14436 369860 14464
rect 278004 14424 278010 14436
rect 369854 14424 369860 14436
rect 369912 14424 369918 14476
rect 420178 14424 420184 14476
rect 420236 14464 420242 14476
rect 456978 14464 456984 14476
rect 420236 14436 456984 14464
rect 420236 14424 420242 14436
rect 456978 14424 456984 14436
rect 457036 14424 457042 14476
rect 475746 14424 475752 14476
rect 475804 14464 475810 14476
rect 491294 14464 491300 14476
rect 475804 14436 491300 14464
rect 475804 14424 475810 14436
rect 491294 14424 491300 14436
rect 491352 14424 491358 14476
rect 543918 14424 543924 14476
rect 543976 14464 543982 14476
rect 562042 14464 562048 14476
rect 543976 14436 562048 14464
rect 543976 14424 543982 14436
rect 562042 14424 562048 14436
rect 562100 14424 562106 14476
rect 81618 13540 81624 13592
rect 81676 13580 81682 13592
rect 214558 13580 214564 13592
rect 81676 13552 214564 13580
rect 81676 13540 81682 13552
rect 214558 13540 214564 13552
rect 214616 13540 214622 13592
rect 109034 13472 109040 13524
rect 109092 13512 109098 13524
rect 266446 13512 266452 13524
rect 109092 13484 266452 13512
rect 109092 13472 109098 13484
rect 266446 13472 266452 13484
rect 266504 13472 266510 13524
rect 102226 13404 102232 13456
rect 102284 13444 102290 13456
rect 262306 13444 262312 13456
rect 102284 13416 262312 13444
rect 102284 13404 102290 13416
rect 262306 13404 262312 13416
rect 262364 13404 262370 13456
rect 94682 13336 94688 13388
rect 94740 13376 94746 13388
rect 258166 13376 258172 13388
rect 94740 13348 258172 13376
rect 94740 13336 94746 13348
rect 258166 13336 258172 13348
rect 258224 13336 258230 13388
rect 91554 13268 91560 13320
rect 91612 13308 91618 13320
rect 255406 13308 255412 13320
rect 91612 13280 255412 13308
rect 91612 13268 91618 13280
rect 255406 13268 255412 13280
rect 255464 13268 255470 13320
rect 87506 13200 87512 13252
rect 87564 13240 87570 13252
rect 252646 13240 252652 13252
rect 87564 13212 252652 13240
rect 87564 13200 87570 13212
rect 252646 13200 252652 13212
rect 252704 13200 252710 13252
rect 349154 13200 349160 13252
rect 349212 13240 349218 13252
rect 412726 13240 412732 13252
rect 349212 13212 412732 13240
rect 349212 13200 349218 13212
rect 412726 13200 412732 13212
rect 412784 13200 412790 13252
rect 80882 13132 80888 13184
rect 80940 13172 80946 13184
rect 248506 13172 248512 13184
rect 80940 13144 248512 13172
rect 80940 13132 80946 13144
rect 248506 13132 248512 13144
rect 248564 13132 248570 13184
rect 297450 13132 297456 13184
rect 297508 13172 297514 13184
rect 374178 13172 374184 13184
rect 297508 13144 374184 13172
rect 297508 13132 297514 13144
rect 374178 13132 374184 13144
rect 374236 13132 374242 13184
rect 77386 13064 77392 13116
rect 77444 13104 77450 13116
rect 247126 13104 247132 13116
rect 77444 13076 247132 13104
rect 77444 13064 77450 13076
rect 247126 13064 247132 13076
rect 247184 13064 247190 13116
rect 294690 13064 294696 13116
rect 294748 13104 294754 13116
rect 378134 13104 378140 13116
rect 294748 13076 378140 13104
rect 294748 13064 294754 13076
rect 378134 13064 378140 13076
rect 378192 13064 378198 13116
rect 421006 13064 421012 13116
rect 421064 13104 421070 13116
rect 456886 13104 456892 13116
rect 421064 13076 456892 13104
rect 421064 13064 421070 13076
rect 456886 13064 456892 13076
rect 456944 13064 456950 13116
rect 56778 12180 56784 12232
rect 56836 12220 56842 12232
rect 234614 12220 234620 12232
rect 56836 12192 234620 12220
rect 56836 12180 56842 12192
rect 234614 12180 234620 12192
rect 234672 12180 234678 12232
rect 50154 12112 50160 12164
rect 50212 12152 50218 12164
rect 230474 12152 230480 12164
rect 50212 12124 230480 12152
rect 50212 12112 50218 12124
rect 230474 12112 230480 12124
rect 230532 12112 230538 12164
rect 41874 12044 41880 12096
rect 41932 12084 41938 12096
rect 224954 12084 224960 12096
rect 41932 12056 224960 12084
rect 41932 12044 41938 12056
rect 224954 12044 224960 12056
rect 225012 12044 225018 12096
rect 31938 11976 31944 12028
rect 31996 12016 32002 12028
rect 219434 12016 219440 12028
rect 31996 11988 219440 12016
rect 31996 11976 32002 11988
rect 219434 11976 219440 11988
rect 219492 11976 219498 12028
rect 18598 11908 18604 11960
rect 18656 11948 18662 11960
rect 208486 11948 208492 11960
rect 18656 11920 208492 11948
rect 18656 11908 18662 11920
rect 208486 11908 208492 11920
rect 208544 11908 208550 11960
rect 234614 11908 234620 11960
rect 234672 11948 234678 11960
rect 343726 11948 343732 11960
rect 234672 11920 343732 11948
rect 234672 11908 234678 11920
rect 343726 11908 343732 11920
rect 343784 11908 343790 11960
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 205818 11880 205824 11892
rect 9732 11852 205824 11880
rect 9732 11840 9738 11852
rect 205818 11840 205824 11852
rect 205876 11840 205882 11892
rect 231026 11840 231032 11892
rect 231084 11880 231090 11892
rect 340874 11880 340880 11892
rect 231084 11852 340880 11880
rect 231084 11840 231090 11852
rect 340874 11840 340880 11852
rect 340932 11840 340938 11892
rect 5994 11772 6000 11824
rect 6052 11812 6058 11824
rect 202966 11812 202972 11824
rect 6052 11784 202972 11812
rect 6052 11772 6058 11784
rect 202966 11772 202972 11784
rect 203024 11772 203030 11824
rect 223574 11772 223580 11824
rect 223632 11812 223638 11824
rect 336734 11812 336740 11824
rect 223632 11784 336740 11812
rect 223632 11772 223638 11784
rect 336734 11772 336740 11784
rect 336792 11772 336798 11824
rect 337378 11772 337384 11824
rect 337436 11812 337442 11824
rect 397454 11812 397460 11824
rect 337436 11784 397460 11812
rect 337436 11772 337442 11784
rect 397454 11772 397460 11784
rect 397512 11772 397518 11824
rect 113818 11704 113824 11756
rect 113876 11744 113882 11756
rect 200114 11744 200120 11756
rect 113876 11716 200120 11744
rect 113876 11704 113882 11716
rect 200114 11704 200120 11716
rect 200172 11704 200178 11756
rect 219986 11704 219992 11756
rect 220044 11744 220050 11756
rect 333974 11744 333980 11756
rect 220044 11716 333980 11744
rect 220044 11704 220050 11716
rect 333974 11704 333980 11716
rect 334032 11704 334038 11756
rect 345290 11704 345296 11756
rect 345348 11744 345354 11756
rect 411254 11744 411260 11756
rect 345348 11716 411260 11744
rect 345348 11704 345354 11716
rect 411254 11704 411260 11716
rect 411312 11704 411318 11756
rect 423858 11704 423864 11756
rect 423916 11744 423922 11756
rect 459646 11744 459652 11756
rect 423916 11716 459652 11744
rect 423916 11704 423922 11716
rect 459646 11704 459652 11716
rect 459704 11704 459710 11756
rect 160094 11636 160100 11688
rect 160152 11676 160158 11688
rect 161290 11676 161296 11688
rect 160152 11648 161296 11676
rect 160152 11636 160158 11648
rect 161290 11636 161296 11648
rect 161348 11636 161354 11688
rect 188522 10888 188528 10940
rect 188580 10928 188586 10940
rect 314838 10928 314844 10940
rect 188580 10900 314844 10928
rect 188580 10888 188586 10900
rect 314838 10888 314844 10900
rect 314896 10888 314902 10940
rect 180978 10820 180984 10872
rect 181036 10860 181042 10872
rect 310514 10860 310520 10872
rect 181036 10832 310520 10860
rect 181036 10820 181042 10832
rect 310514 10820 310520 10832
rect 310572 10820 310578 10872
rect 95786 10752 95792 10804
rect 95844 10792 95850 10804
rect 175182 10792 175188 10804
rect 95844 10764 175188 10792
rect 95844 10752 95850 10764
rect 175182 10752 175188 10764
rect 175240 10752 175246 10804
rect 177574 10752 177580 10804
rect 177632 10792 177638 10804
rect 307754 10792 307760 10804
rect 177632 10764 307760 10792
rect 177632 10752 177638 10764
rect 307754 10752 307760 10764
rect 307812 10752 307818 10804
rect 74994 10684 75000 10736
rect 75052 10724 75058 10736
rect 170766 10724 170772 10736
rect 75052 10696 170772 10724
rect 75052 10684 75058 10696
rect 170766 10684 170772 10696
rect 170824 10684 170830 10736
rect 173894 10684 173900 10736
rect 173952 10724 173958 10736
rect 306374 10724 306380 10736
rect 173952 10696 306380 10724
rect 173952 10684 173958 10696
rect 306374 10684 306380 10696
rect 306432 10684 306438 10736
rect 170306 10616 170312 10668
rect 170364 10656 170370 10668
rect 303614 10656 303620 10668
rect 170364 10628 303620 10656
rect 170364 10616 170370 10628
rect 303614 10616 303620 10628
rect 303672 10616 303678 10668
rect 111610 10548 111616 10600
rect 111668 10588 111674 10600
rect 267734 10588 267740 10600
rect 111668 10560 267740 10588
rect 111668 10548 111674 10560
rect 267734 10548 267740 10560
rect 267792 10548 267798 10600
rect 104066 10480 104072 10532
rect 104124 10520 104130 10532
rect 263594 10520 263600 10532
rect 104124 10492 263600 10520
rect 104124 10480 104130 10492
rect 263594 10480 263600 10492
rect 263652 10480 263658 10532
rect 64322 10412 64328 10464
rect 64380 10452 64386 10464
rect 233878 10452 233884 10464
rect 64380 10424 233884 10452
rect 64380 10412 64386 10424
rect 233878 10412 233884 10424
rect 233936 10412 233942 10464
rect 36722 10344 36728 10396
rect 36780 10384 36786 10396
rect 222194 10384 222200 10396
rect 36780 10356 222200 10384
rect 36780 10344 36786 10356
rect 222194 10344 222200 10356
rect 222252 10344 222258 10396
rect 349246 10344 349252 10396
rect 349304 10384 349310 10396
rect 414014 10384 414020 10396
rect 349304 10356 414020 10384
rect 349304 10344 349310 10356
rect 414014 10344 414020 10356
rect 414072 10344 414078 10396
rect 442626 10344 442632 10396
rect 442684 10384 442690 10396
rect 470686 10384 470692 10396
rect 442684 10356 470692 10384
rect 442684 10344 442690 10356
rect 470686 10344 470692 10356
rect 470744 10344 470750 10396
rect 17954 10276 17960 10328
rect 18012 10316 18018 10328
rect 211154 10316 211160 10328
rect 18012 10288 211160 10316
rect 18012 10276 18018 10288
rect 211154 10276 211160 10288
rect 211212 10276 211218 10328
rect 314746 10276 314752 10328
rect 314804 10316 314810 10328
rect 391934 10316 391940 10328
rect 314804 10288 391940 10316
rect 314804 10276 314810 10288
rect 391934 10276 391940 10288
rect 391992 10276 391998 10328
rect 409138 10276 409144 10328
rect 409196 10316 409202 10328
rect 449986 10316 449992 10328
rect 409196 10288 449992 10316
rect 409196 10276 409202 10288
rect 449986 10276 449992 10288
rect 450044 10276 450050 10328
rect 473906 10276 473912 10328
rect 473964 10316 473970 10328
rect 490006 10316 490012 10328
rect 473964 10288 490012 10316
rect 473964 10276 473970 10288
rect 490006 10276 490012 10288
rect 490064 10276 490070 10328
rect 490098 10276 490104 10328
rect 490156 10316 490162 10328
rect 499666 10316 499672 10328
rect 490156 10288 499672 10316
rect 490156 10276 490162 10288
rect 499666 10276 499672 10288
rect 499724 10276 499730 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 78582 9392 78588 9444
rect 78640 9432 78646 9444
rect 247034 9432 247040 9444
rect 78640 9404 247040 9432
rect 78640 9392 78646 9404
rect 247034 9392 247040 9404
rect 247092 9392 247098 9444
rect 66714 9324 66720 9376
rect 66772 9364 66778 9376
rect 240134 9364 240140 9376
rect 66772 9336 240140 9364
rect 66772 9324 66778 9336
rect 240134 9324 240140 9336
rect 240192 9324 240198 9376
rect 59630 9256 59636 9308
rect 59688 9296 59694 9308
rect 235994 9296 236000 9308
rect 59688 9268 236000 9296
rect 59688 9256 59694 9268
rect 235994 9256 236000 9268
rect 236052 9256 236058 9308
rect 286594 9256 286600 9308
rect 286652 9296 286658 9308
rect 375374 9296 375380 9308
rect 286652 9268 375380 9296
rect 286652 9256 286658 9268
rect 375374 9256 375380 9268
rect 375432 9256 375438 9308
rect 56042 9188 56048 9240
rect 56100 9228 56106 9240
rect 233234 9228 233240 9240
rect 56100 9200 233240 9228
rect 56100 9188 56106 9200
rect 233234 9188 233240 9200
rect 233292 9188 233298 9240
rect 261754 9188 261760 9240
rect 261812 9228 261818 9240
rect 360286 9228 360292 9240
rect 261812 9200 360292 9228
rect 261812 9188 261818 9200
rect 360286 9188 360292 9200
rect 360344 9188 360350 9240
rect 52546 9120 52552 9172
rect 52604 9160 52610 9172
rect 231946 9160 231952 9172
rect 52604 9132 231952 9160
rect 52604 9120 52610 9132
rect 231946 9120 231952 9132
rect 232004 9120 232010 9172
rect 258258 9120 258264 9172
rect 258316 9160 258322 9172
rect 357526 9160 357532 9172
rect 258316 9132 357532 9160
rect 258316 9120 258322 9132
rect 357526 9120 357532 9132
rect 357584 9120 357590 9172
rect 31294 9052 31300 9104
rect 31352 9092 31358 9104
rect 218146 9092 218152 9104
rect 31352 9064 218152 9092
rect 31352 9052 31358 9064
rect 218146 9052 218152 9064
rect 218204 9052 218210 9104
rect 251174 9052 251180 9104
rect 251232 9092 251238 9104
rect 353294 9092 353300 9104
rect 251232 9064 353300 9092
rect 251232 9052 251238 9064
rect 353294 9052 353300 9064
rect 353352 9052 353358 9104
rect 27706 8984 27712 9036
rect 27764 9024 27770 9036
rect 216858 9024 216864 9036
rect 27764 8996 216864 9024
rect 27764 8984 27770 8996
rect 216858 8984 216864 8996
rect 216916 8984 216922 9036
rect 247586 8984 247592 9036
rect 247644 9024 247650 9036
rect 350626 9024 350632 9036
rect 247644 8996 350632 9024
rect 247644 8984 247650 8996
rect 350626 8984 350632 8996
rect 350684 8984 350690 9036
rect 416682 8984 416688 9036
rect 416740 9024 416746 9036
rect 454034 9024 454040 9036
rect 416740 8996 454040 9024
rect 416740 8984 416746 8996
rect 454034 8984 454040 8996
rect 454092 8984 454098 9036
rect 480530 8984 480536 9036
rect 480588 9024 480594 9036
rect 494146 9024 494152 9036
rect 480588 8996 494152 9024
rect 480588 8984 480594 8996
rect 494146 8984 494152 8996
rect 494204 8984 494210 9036
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 207106 8956 207112 8968
rect 13596 8928 207112 8956
rect 13596 8916 13602 8928
rect 207106 8916 207112 8928
rect 207164 8916 207170 8968
rect 240502 8916 240508 8968
rect 240560 8956 240566 8968
rect 346486 8956 346492 8968
rect 240560 8928 346492 8956
rect 240560 8916 240566 8928
rect 346486 8916 346492 8928
rect 346544 8916 346550 8968
rect 359918 8916 359924 8968
rect 359976 8956 359982 8968
rect 419534 8956 419540 8968
rect 359976 8928 419540 8956
rect 359976 8916 359982 8928
rect 419534 8916 419540 8928
rect 419592 8916 419598 8968
rect 459186 8916 459192 8968
rect 459244 8956 459250 8968
rect 480438 8956 480444 8968
rect 459244 8928 480444 8956
rect 459244 8916 459250 8928
rect 480438 8916 480444 8928
rect 480496 8916 480502 8968
rect 532694 8916 532700 8968
rect 532752 8956 532758 8968
rect 543182 8956 543188 8968
rect 532752 8928 543188 8956
rect 532752 8916 532758 8928
rect 543182 8916 543188 8928
rect 543240 8916 543246 8968
rect 550726 8916 550732 8968
rect 550784 8956 550790 8968
rect 572714 8956 572720 8968
rect 550784 8928 572720 8956
rect 550784 8916 550790 8928
rect 572714 8916 572720 8928
rect 572772 8916 572778 8968
rect 151906 8100 151912 8152
rect 151964 8140 151970 8152
rect 292666 8140 292672 8152
rect 151964 8112 292672 8140
rect 151964 8100 151970 8112
rect 292666 8100 292672 8112
rect 292724 8100 292730 8152
rect 145926 8032 145932 8084
rect 145984 8072 145990 8084
rect 287698 8072 287704 8084
rect 145984 8044 287704 8072
rect 145984 8032 145990 8044
rect 287698 8032 287704 8044
rect 287756 8032 287762 8084
rect 134150 7964 134156 8016
rect 134208 8004 134214 8016
rect 281534 8004 281540 8016
rect 134208 7976 281540 8004
rect 134208 7964 134214 7976
rect 281534 7964 281540 7976
rect 281592 7964 281598 8016
rect 325602 7964 325608 8016
rect 325660 8004 325666 8016
rect 398834 8004 398840 8016
rect 325660 7976 398840 8004
rect 325660 7964 325666 7976
rect 398834 7964 398840 7976
rect 398892 7964 398898 8016
rect 130562 7896 130568 7948
rect 130620 7936 130626 7948
rect 278866 7936 278872 7948
rect 130620 7908 278872 7936
rect 130620 7896 130626 7908
rect 278866 7896 278872 7908
rect 278924 7896 278930 7948
rect 322106 7896 322112 7948
rect 322164 7936 322170 7948
rect 396074 7936 396080 7948
rect 322164 7908 396080 7936
rect 322164 7896 322170 7908
rect 396074 7896 396080 7908
rect 396132 7896 396138 7948
rect 123478 7828 123484 7880
rect 123536 7868 123542 7880
rect 274726 7868 274732 7880
rect 123536 7840 274732 7868
rect 123536 7828 123542 7840
rect 274726 7828 274732 7840
rect 274784 7828 274790 7880
rect 307938 7828 307944 7880
rect 307996 7868 308002 7880
rect 387978 7868 387984 7880
rect 307996 7840 387984 7868
rect 307996 7828 308002 7840
rect 387978 7828 387984 7840
rect 388036 7828 388042 7880
rect 122282 7760 122288 7812
rect 122340 7800 122346 7812
rect 274634 7800 274640 7812
rect 122340 7772 274640 7800
rect 122340 7760 122346 7772
rect 274634 7760 274640 7772
rect 274692 7760 274698 7812
rect 311434 7760 311440 7812
rect 311492 7800 311498 7812
rect 390554 7800 390560 7812
rect 311492 7772 390560 7800
rect 311492 7760 311498 7772
rect 390554 7760 390560 7772
rect 390612 7760 390618 7812
rect 72602 7692 72608 7744
rect 72660 7732 72666 7744
rect 244366 7732 244372 7744
rect 72660 7704 244372 7732
rect 72660 7692 72666 7704
rect 244366 7692 244372 7704
rect 244424 7692 244430 7744
rect 304350 7692 304356 7744
rect 304408 7732 304414 7744
rect 386506 7732 386512 7744
rect 304408 7704 386512 7732
rect 304408 7692 304414 7704
rect 386506 7692 386512 7704
rect 386564 7692 386570 7744
rect 14734 7624 14740 7676
rect 14792 7664 14798 7676
rect 208394 7664 208400 7676
rect 14792 7636 208400 7664
rect 14792 7624 14798 7636
rect 208394 7624 208400 7636
rect 208452 7624 208458 7676
rect 300762 7624 300768 7676
rect 300820 7664 300826 7676
rect 383746 7664 383752 7676
rect 300820 7636 383752 7664
rect 300820 7624 300826 7636
rect 383746 7624 383752 7636
rect 383804 7624 383810 7676
rect 435542 7624 435548 7676
rect 435600 7664 435606 7676
rect 466546 7664 466552 7676
rect 435600 7636 466552 7664
rect 435600 7624 435606 7636
rect 466546 7624 466552 7636
rect 466604 7624 466610 7676
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 201494 7596 201500 7608
rect 4120 7568 201500 7596
rect 4120 7556 4126 7568
rect 201494 7556 201500 7568
rect 201552 7556 201558 7608
rect 293678 7556 293684 7608
rect 293736 7596 293742 7608
rect 379514 7596 379520 7608
rect 293736 7568 379520 7596
rect 293736 7556 293742 7568
rect 379514 7556 379520 7568
rect 379572 7556 379578 7608
rect 402514 7556 402520 7608
rect 402572 7596 402578 7608
rect 445846 7596 445852 7608
rect 402572 7568 445852 7596
rect 402572 7556 402578 7568
rect 445846 7556 445852 7568
rect 445904 7556 445910 7608
rect 462774 7556 462780 7608
rect 462832 7596 462838 7608
rect 483106 7596 483112 7608
rect 462832 7568 483112 7596
rect 462832 7556 462838 7568
rect 483106 7556 483112 7568
rect 483164 7556 483170 7608
rect 540974 7556 540980 7608
rect 541032 7596 541038 7608
rect 558546 7596 558552 7608
rect 541032 7568 558552 7596
rect 541032 7556 541038 7568
rect 558546 7556 558552 7568
rect 558604 7556 558610 7608
rect 374086 7488 374092 7540
rect 374144 7528 374150 7540
rect 375282 7528 375288 7540
rect 374144 7500 375288 7528
rect 374144 7488 374150 7500
rect 375282 7488 375288 7500
rect 375340 7488 375346 7540
rect 570598 6808 570604 6860
rect 570656 6848 570662 6860
rect 580166 6848 580172 6860
rect 570656 6820 580172 6848
rect 570656 6808 570662 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 98638 6604 98644 6656
rect 98696 6644 98702 6656
rect 259546 6644 259552 6656
rect 98696 6616 259552 6644
rect 98696 6604 98702 6616
rect 259546 6604 259552 6616
rect 259604 6604 259610 6656
rect 83274 6536 83280 6588
rect 83332 6576 83338 6588
rect 249886 6576 249892 6588
rect 83332 6548 249892 6576
rect 83332 6536 83338 6548
rect 249886 6536 249892 6548
rect 249944 6536 249950 6588
rect 76190 6468 76196 6520
rect 76248 6508 76254 6520
rect 246022 6508 246028 6520
rect 76248 6480 246028 6508
rect 76248 6468 76254 6480
rect 246022 6468 246028 6480
rect 246080 6468 246086 6520
rect 79686 6400 79692 6452
rect 79744 6440 79750 6452
rect 248414 6440 248420 6452
rect 79744 6412 248420 6440
rect 79744 6400 79750 6412
rect 248414 6400 248420 6412
rect 248472 6400 248478 6452
rect 71498 6332 71504 6384
rect 71556 6372 71562 6384
rect 242894 6372 242900 6384
rect 71556 6344 242900 6372
rect 71556 6332 71562 6344
rect 242894 6332 242900 6344
rect 242952 6332 242958 6384
rect 288986 6332 288992 6384
rect 289044 6372 289050 6384
rect 376754 6372 376760 6384
rect 289044 6344 376760 6372
rect 289044 6332 289050 6344
rect 376754 6332 376760 6344
rect 376812 6332 376818 6384
rect 44266 6264 44272 6316
rect 44324 6304 44330 6316
rect 226610 6304 226616 6316
rect 44324 6276 226616 6304
rect 44324 6264 44330 6276
rect 226610 6264 226616 6276
rect 226668 6264 226674 6316
rect 285398 6264 285404 6316
rect 285456 6304 285462 6316
rect 373994 6304 374000 6316
rect 285456 6276 374000 6304
rect 285456 6264 285462 6276
rect 373994 6264 374000 6276
rect 374052 6264 374058 6316
rect 381170 6264 381176 6316
rect 381228 6304 381234 6316
rect 433334 6304 433340 6316
rect 381228 6276 433340 6304
rect 381228 6264 381234 6276
rect 433334 6264 433340 6276
rect 433392 6264 433398 6316
rect 30098 6196 30104 6248
rect 30156 6236 30162 6248
rect 218054 6236 218060 6248
rect 30156 6208 218060 6236
rect 30156 6196 30162 6208
rect 218054 6196 218060 6208
rect 218112 6196 218118 6248
rect 274818 6196 274824 6248
rect 274876 6236 274882 6248
rect 367094 6236 367100 6248
rect 274876 6208 367100 6236
rect 274876 6196 274882 6208
rect 367094 6196 367100 6208
rect 367152 6196 367158 6248
rect 377674 6196 377680 6248
rect 377732 6236 377738 6248
rect 430758 6236 430764 6248
rect 377732 6208 430764 6236
rect 377732 6196 377738 6208
rect 430758 6196 430764 6208
rect 430816 6196 430822 6248
rect 466270 6196 466276 6248
rect 466328 6236 466334 6248
rect 484486 6236 484492 6248
rect 466328 6208 484492 6236
rect 466328 6196 466334 6208
rect 484486 6196 484492 6208
rect 484544 6196 484550 6248
rect 536926 6196 536932 6248
rect 536984 6236 536990 6248
rect 551462 6236 551468 6248
rect 536984 6208 551468 6236
rect 536984 6196 536990 6208
rect 551462 6196 551468 6208
rect 551520 6196 551526 6248
rect 21818 6128 21824 6180
rect 21876 6168 21882 6180
rect 212718 6168 212724 6180
rect 21876 6140 212724 6168
rect 21876 6128 21882 6140
rect 212718 6128 212724 6140
rect 212776 6128 212782 6180
rect 257062 6128 257068 6180
rect 257120 6168 257126 6180
rect 357526 6168 357532 6180
rect 257120 6140 357532 6168
rect 257120 6128 257126 6140
rect 357526 6128 357532 6140
rect 357584 6128 357590 6180
rect 367002 6128 367008 6180
rect 367060 6168 367066 6180
rect 423674 6168 423680 6180
rect 367060 6140 423680 6168
rect 367060 6128 367066 6140
rect 423674 6128 423680 6140
rect 423732 6128 423738 6180
rect 437934 6128 437940 6180
rect 437992 6168 437998 6180
rect 467926 6168 467932 6180
rect 437992 6140 467932 6168
rect 437992 6128 437998 6140
rect 467926 6128 467932 6140
rect 467984 6128 467990 6180
rect 495894 6128 495900 6180
rect 495952 6168 495958 6180
rect 503806 6168 503812 6180
rect 495952 6140 503812 6168
rect 495952 6128 495958 6140
rect 503806 6128 503812 6140
rect 503864 6128 503870 6180
rect 547966 6128 547972 6180
rect 548024 6168 548030 6180
rect 569126 6168 569132 6180
rect 548024 6140 569132 6168
rect 548024 6128 548030 6140
rect 569126 6128 569132 6140
rect 569184 6128 569190 6180
rect 197906 5312 197912 5364
rect 197964 5352 197970 5364
rect 320174 5352 320180 5364
rect 197964 5324 320180 5352
rect 197964 5312 197970 5324
rect 320174 5312 320180 5324
rect 320232 5312 320238 5364
rect 156598 5244 156604 5296
rect 156656 5284 156662 5296
rect 284938 5284 284944 5296
rect 156656 5256 284944 5284
rect 156656 5244 156662 5256
rect 284938 5244 284944 5256
rect 284996 5244 285002 5296
rect 118786 5176 118792 5228
rect 118844 5216 118850 5228
rect 266998 5216 267004 5228
rect 118844 5188 267004 5216
rect 118844 5176 118850 5188
rect 266998 5176 267004 5188
rect 267056 5176 267062 5228
rect 101030 5108 101036 5160
rect 101088 5148 101094 5160
rect 260834 5148 260840 5160
rect 101088 5120 260840 5148
rect 101088 5108 101094 5120
rect 260834 5108 260840 5120
rect 260892 5108 260898 5160
rect 399018 5108 399024 5160
rect 399076 5148 399082 5160
rect 442994 5148 443000 5160
rect 399076 5120 443000 5148
rect 399076 5108 399082 5120
rect 442994 5108 443000 5120
rect 443052 5108 443058 5160
rect 73798 5040 73804 5092
rect 73856 5080 73862 5092
rect 244274 5080 244280 5092
rect 73856 5052 244280 5080
rect 73856 5040 73862 5052
rect 244274 5040 244280 5052
rect 244332 5040 244338 5092
rect 391842 5040 391848 5092
rect 391900 5080 391906 5092
rect 438946 5080 438952 5092
rect 391900 5052 438952 5080
rect 391900 5040 391906 5052
rect 438946 5040 438952 5052
rect 439004 5040 439010 5092
rect 65518 4972 65524 5024
rect 65576 5012 65582 5024
rect 238846 5012 238852 5024
rect 65576 4984 238852 5012
rect 65576 4972 65582 4984
rect 238846 4972 238852 4984
rect 238904 4972 238910 5024
rect 388254 4972 388260 5024
rect 388312 5012 388318 5024
rect 437474 5012 437480 5024
rect 388312 4984 437480 5012
rect 388312 4972 388318 4984
rect 437474 4972 437480 4984
rect 437532 4972 437538 5024
rect 53742 4904 53748 4956
rect 53800 4944 53806 4956
rect 231118 4944 231124 4956
rect 53800 4916 231124 4944
rect 53800 4904 53806 4916
rect 231118 4904 231124 4916
rect 231176 4904 231182 4956
rect 374178 4904 374184 4956
rect 374236 4944 374242 4956
rect 427906 4944 427912 4956
rect 374236 4916 427912 4944
rect 374236 4904 374242 4916
rect 427906 4904 427912 4916
rect 427964 4904 427970 4956
rect 12342 4836 12348 4888
rect 12400 4876 12406 4888
rect 207014 4876 207020 4888
rect 12400 4848 207020 4876
rect 12400 4836 12406 4848
rect 207014 4836 207020 4848
rect 207072 4836 207078 4888
rect 268838 4836 268844 4888
rect 268896 4876 268902 4888
rect 364426 4876 364432 4888
rect 268896 4848 364432 4876
rect 268896 4836 268902 4848
rect 364426 4836 364432 4848
rect 364484 4836 364490 4888
rect 370590 4836 370596 4888
rect 370648 4876 370654 4888
rect 426526 4876 426532 4888
rect 370648 4848 426532 4876
rect 370648 4836 370654 4848
rect 426526 4836 426532 4848
rect 426584 4836 426590 4888
rect 469858 4836 469864 4888
rect 469916 4876 469922 4888
rect 487154 4876 487160 4888
rect 469916 4848 487160 4876
rect 469916 4836 469922 4848
rect 487154 4836 487160 4848
rect 487212 4836 487218 4888
rect 547138 4836 547144 4888
rect 547196 4876 547202 4888
rect 547874 4876 547880 4888
rect 547196 4848 547880 4876
rect 547196 4836 547202 4848
rect 547874 4836 547880 4848
rect 547932 4836 547938 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 200206 4808 200212 4820
rect 1728 4780 200212 4808
rect 1728 4768 1734 4780
rect 200206 4768 200212 4780
rect 200264 4768 200270 4820
rect 201494 4768 201500 4820
rect 201552 4808 201558 4820
rect 322934 4808 322940 4820
rect 201552 4780 322940 4808
rect 201552 4768 201558 4780
rect 322934 4768 322940 4780
rect 322992 4768 322998 4820
rect 356330 4768 356336 4820
rect 356388 4808 356394 4820
rect 418154 4808 418160 4820
rect 356388 4780 418160 4808
rect 356388 4768 356394 4780
rect 418154 4768 418160 4780
rect 418212 4768 418218 4820
rect 452102 4768 452108 4820
rect 452160 4808 452166 4820
rect 476298 4808 476304 4820
rect 452160 4780 476304 4808
rect 452160 4768 452166 4780
rect 476298 4768 476304 4780
rect 476356 4768 476362 4820
rect 492306 4768 492312 4820
rect 492364 4808 492370 4820
rect 501046 4808 501052 4820
rect 492364 4780 501052 4808
rect 492364 4768 492370 4780
rect 501046 4768 501052 4780
rect 501104 4768 501110 4820
rect 539686 4768 539692 4820
rect 539744 4808 539750 4820
rect 554958 4808 554964 4820
rect 539744 4780 554964 4808
rect 539744 4768 539750 4780
rect 554958 4768 554964 4780
rect 555016 4768 555022 4820
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 18598 4128 18604 4140
rect 15988 4100 18604 4128
rect 15988 4088 15994 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 265342 4088 265348 4140
rect 265400 4128 265406 4140
rect 269758 4128 269764 4140
rect 265400 4100 269764 4128
rect 265400 4088 265406 4100
rect 269758 4088 269764 4100
rect 269816 4088 269822 4140
rect 296070 4088 296076 4140
rect 296128 4128 296134 4140
rect 297358 4128 297364 4140
rect 296128 4100 297364 4128
rect 296128 4088 296134 4100
rect 297358 4088 297364 4100
rect 297416 4088 297422 4140
rect 376478 4088 376484 4140
rect 376536 4128 376542 4140
rect 377398 4128 377404 4140
rect 376536 4100 377404 4128
rect 376536 4088 376542 4100
rect 377398 4088 377404 4100
rect 377456 4088 377462 4140
rect 383562 4088 383568 4140
rect 383620 4128 383626 4140
rect 384298 4128 384304 4140
rect 383620 4100 384304 4128
rect 383620 4088 383626 4100
rect 384298 4088 384304 4100
rect 384356 4088 384362 4140
rect 479334 4088 479340 4140
rect 479392 4128 479398 4140
rect 482278 4128 482284 4140
rect 479392 4100 482284 4128
rect 479392 4088 479398 4100
rect 482278 4088 482284 4100
rect 482336 4088 482342 4140
rect 527266 4088 527272 4140
rect 527324 4128 527330 4140
rect 527910 4128 527916 4140
rect 527324 4100 527916 4128
rect 527324 4088 527330 4100
rect 527910 4088 527916 4100
rect 527968 4088 527974 4140
rect 537478 4088 537484 4140
rect 537536 4128 537542 4140
rect 549070 4128 549076 4140
rect 537536 4100 549076 4128
rect 537536 4088 537542 4100
rect 549070 4088 549076 4100
rect 549128 4088 549134 4140
rect 135254 4020 135260 4072
rect 135312 4060 135318 4072
rect 136450 4060 136456 4072
rect 135312 4032 136456 4060
rect 135312 4020 135318 4032
rect 136450 4020 136456 4032
rect 136508 4020 136514 4072
rect 151814 4020 151820 4072
rect 151872 4060 151878 4072
rect 153010 4060 153016 4072
rect 151872 4032 153016 4060
rect 151872 4020 151878 4032
rect 153010 4020 153016 4032
rect 153068 4020 153074 4072
rect 241698 4020 241704 4072
rect 241756 4060 241762 4072
rect 250622 4060 250628 4072
rect 241756 4032 250628 4060
rect 241756 4020 241762 4032
rect 250622 4020 250628 4032
rect 250680 4020 250686 4072
rect 523034 4020 523040 4072
rect 523092 4060 523098 4072
rect 529014 4060 529020 4072
rect 523092 4032 529020 4060
rect 523092 4020 523098 4032
rect 529014 4020 529020 4032
rect 529072 4020 529078 4072
rect 536834 4020 536840 4072
rect 536892 4060 536898 4072
rect 550266 4060 550272 4072
rect 536892 4032 550272 4060
rect 536892 4020 536898 4032
rect 550266 4020 550272 4032
rect 550324 4020 550330 4072
rect 124674 3952 124680 4004
rect 124732 3992 124738 4004
rect 169386 3992 169392 4004
rect 124732 3964 169392 3992
rect 124732 3952 124738 3964
rect 169386 3952 169392 3964
rect 169444 3952 169450 4004
rect 538214 3952 538220 4004
rect 538272 3992 538278 4004
rect 553762 3992 553768 4004
rect 538272 3964 553768 3992
rect 538272 3952 538278 3964
rect 553762 3952 553768 3964
rect 553820 3952 553826 4004
rect 114002 3884 114008 3936
rect 114060 3924 114066 3936
rect 188614 3924 188620 3936
rect 114060 3896 188620 3924
rect 114060 3884 114066 3896
rect 188614 3884 188620 3896
rect 188672 3884 188678 3936
rect 534718 3884 534724 3936
rect 534776 3924 534782 3936
rect 538398 3924 538404 3936
rect 534776 3896 538404 3924
rect 534776 3884 534782 3896
rect 538398 3884 538404 3896
rect 538456 3884 538462 3936
rect 539594 3884 539600 3936
rect 539652 3924 539658 3936
rect 556154 3924 556160 3936
rect 539652 3896 556160 3924
rect 539652 3884 539658 3896
rect 556154 3884 556160 3896
rect 556212 3884 556218 3936
rect 43070 3816 43076 3868
rect 43128 3856 43134 3868
rect 173526 3856 173532 3868
rect 43128 3828 173532 3856
rect 43128 3816 43134 3828
rect 173526 3816 173532 3828
rect 173584 3816 173590 3868
rect 276014 3816 276020 3868
rect 276072 3856 276078 3868
rect 278038 3856 278044 3868
rect 276072 3828 278044 3856
rect 276072 3816 276078 3828
rect 278038 3816 278044 3828
rect 278096 3816 278102 3868
rect 409874 3816 409880 3868
rect 409932 3856 409938 3868
rect 410518 3856 410524 3868
rect 409932 3828 410524 3856
rect 409932 3816 409938 3828
rect 410518 3816 410524 3828
rect 410576 3816 410582 3868
rect 525794 3816 525800 3868
rect 525852 3856 525858 3868
rect 532510 3856 532516 3868
rect 525852 3828 532516 3856
rect 525852 3816 525858 3828
rect 532510 3816 532516 3828
rect 532568 3816 532574 3868
rect 546494 3816 546500 3868
rect 546552 3856 546558 3868
rect 566826 3856 566832 3868
rect 546552 3828 566832 3856
rect 546552 3816 546558 3828
rect 566826 3816 566832 3828
rect 566884 3816 566890 3868
rect 35986 3748 35992 3800
rect 36044 3788 36050 3800
rect 177666 3788 177672 3800
rect 36044 3760 177672 3788
rect 36044 3748 36050 3760
rect 177666 3748 177672 3760
rect 177724 3748 177730 3800
rect 284294 3748 284300 3800
rect 284352 3788 284358 3800
rect 297450 3788 297456 3800
rect 284352 3760 297456 3788
rect 284352 3748 284358 3760
rect 297450 3748 297456 3760
rect 297508 3748 297514 3800
rect 390646 3748 390652 3800
rect 390704 3788 390710 3800
rect 438118 3788 438124 3800
rect 390704 3760 438124 3788
rect 390704 3748 390710 3760
rect 438118 3748 438124 3760
rect 438176 3748 438182 3800
rect 456886 3748 456892 3800
rect 456944 3788 456950 3800
rect 464338 3788 464344 3800
rect 456944 3760 464344 3788
rect 456944 3748 456950 3760
rect 464338 3748 464344 3760
rect 464396 3748 464402 3800
rect 529934 3748 529940 3800
rect 529992 3788 529998 3800
rect 529992 3760 538214 3788
rect 529992 3748 529998 3760
rect 28902 3680 28908 3732
rect 28960 3720 28966 3732
rect 175090 3720 175096 3732
rect 28960 3692 175096 3720
rect 28960 3680 28966 3692
rect 175090 3680 175096 3692
rect 175148 3680 175154 3732
rect 260650 3680 260656 3732
rect 260708 3720 260714 3732
rect 276658 3720 276664 3732
rect 260708 3692 276664 3720
rect 260708 3680 260714 3692
rect 276658 3680 276664 3692
rect 276716 3680 276722 3732
rect 298462 3680 298468 3732
rect 298520 3720 298526 3732
rect 308398 3720 308404 3732
rect 298520 3692 308404 3720
rect 298520 3680 298526 3692
rect 308398 3680 308404 3692
rect 308456 3680 308462 3732
rect 316218 3680 316224 3732
rect 316276 3720 316282 3732
rect 327718 3720 327724 3732
rect 316276 3692 327724 3720
rect 316276 3680 316282 3692
rect 327718 3680 327724 3692
rect 327776 3680 327782 3732
rect 372890 3680 372896 3732
rect 372948 3720 372954 3732
rect 427814 3720 427820 3732
rect 372948 3692 427820 3720
rect 372948 3680 372954 3692
rect 427814 3680 427820 3692
rect 427872 3680 427878 3732
rect 443822 3680 443828 3732
rect 443880 3720 443886 3732
rect 458818 3720 458824 3732
rect 443880 3692 458824 3720
rect 443880 3680 443886 3692
rect 458818 3680 458824 3692
rect 458876 3680 458882 3732
rect 465166 3680 465172 3732
rect 465224 3720 465230 3732
rect 478230 3720 478236 3732
rect 465224 3692 478236 3720
rect 465224 3680 465230 3692
rect 478230 3680 478236 3692
rect 478288 3680 478294 3732
rect 527358 3680 527364 3732
rect 527416 3720 527422 3732
rect 534902 3720 534908 3732
rect 527416 3692 534908 3720
rect 527416 3680 527422 3692
rect 534902 3680 534908 3692
rect 534960 3680 534966 3732
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 172146 3652 172152 3664
rect 20680 3624 172152 3652
rect 20680 3612 20686 3624
rect 172146 3612 172152 3624
rect 172204 3612 172210 3664
rect 225138 3612 225144 3664
rect 225196 3652 225202 3664
rect 236730 3652 236736 3664
rect 225196 3624 236736 3652
rect 225196 3612 225202 3624
rect 236730 3612 236736 3624
rect 236788 3612 236794 3664
rect 252370 3612 252376 3664
rect 252428 3652 252434 3664
rect 273898 3652 273904 3664
rect 252428 3624 273904 3652
rect 252428 3612 252434 3624
rect 273898 3612 273904 3624
rect 273956 3612 273962 3664
rect 277118 3612 277124 3664
rect 277176 3652 277182 3664
rect 286318 3652 286324 3664
rect 277176 3624 286324 3652
rect 277176 3612 277182 3624
rect 286318 3612 286324 3624
rect 286376 3612 286382 3664
rect 294598 3652 294604 3664
rect 287026 3624 294604 3652
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 181438 3584 181444 3596
rect 19484 3556 181444 3584
rect 19484 3544 19490 3556
rect 181438 3544 181444 3556
rect 181496 3544 181502 3596
rect 193214 3544 193220 3596
rect 193272 3584 193278 3596
rect 194410 3584 194416 3596
rect 193272 3556 194416 3584
rect 193272 3544 193278 3556
rect 194410 3544 194416 3556
rect 194468 3544 194474 3596
rect 196618 3544 196624 3596
rect 196676 3544 196682 3596
rect 203886 3544 203892 3596
rect 203944 3584 203950 3596
rect 204898 3584 204904 3596
rect 203944 3556 204904 3584
rect 203944 3544 203950 3556
rect 204898 3544 204904 3556
rect 204956 3544 204962 3596
rect 214466 3544 214472 3596
rect 214524 3584 214530 3596
rect 218698 3584 218704 3596
rect 214524 3556 218704 3584
rect 214524 3544 214530 3556
rect 218698 3544 218704 3556
rect 218756 3544 218762 3596
rect 226978 3584 226984 3596
rect 219406 3556 226984 3584
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 10318 3516 10324 3528
rect 8812 3488 10324 3516
rect 8812 3476 8818 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 196636 3516 196664 3544
rect 11204 3488 196664 3516
rect 11204 3476 11210 3488
rect 213362 3476 213368 3528
rect 213420 3516 213426 3528
rect 214742 3516 214748 3528
rect 213420 3488 214748 3516
rect 213420 3476 213426 3488
rect 214742 3476 214748 3488
rect 214800 3476 214806 3528
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 217318 3516 217324 3528
rect 215720 3488 217324 3516
rect 215720 3476 215726 3488
rect 217318 3476 217324 3488
rect 217376 3476 217382 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 219406 3516 219434 3556
rect 226978 3544 226984 3556
rect 227036 3544 227042 3596
rect 228726 3544 228732 3596
rect 228784 3584 228790 3596
rect 240778 3584 240784 3596
rect 228784 3556 240784 3584
rect 228784 3544 228790 3556
rect 240778 3544 240784 3556
rect 240836 3544 240842 3596
rect 244090 3544 244096 3596
rect 244148 3584 244154 3596
rect 244918 3584 244924 3596
rect 244148 3556 244924 3584
rect 244148 3544 244154 3556
rect 244918 3544 244924 3556
rect 244976 3544 244982 3596
rect 250438 3584 250444 3596
rect 248386 3556 250444 3584
rect 218112 3488 219434 3516
rect 218112 3476 218118 3488
rect 222746 3476 222752 3528
rect 222804 3516 222810 3528
rect 224310 3516 224316 3528
rect 222804 3488 224316 3516
rect 222804 3476 222810 3488
rect 224310 3476 224316 3488
rect 224368 3476 224374 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 228358 3516 228364 3528
rect 226392 3488 228364 3516
rect 226392 3476 226398 3488
rect 228358 3476 228364 3488
rect 228416 3476 228422 3528
rect 235810 3476 235816 3528
rect 235868 3516 235874 3528
rect 236638 3516 236644 3528
rect 235868 3488 236644 3516
rect 235868 3476 235874 3488
rect 236638 3476 236644 3488
rect 236696 3476 236702 3528
rect 248386 3516 248414 3556
rect 250438 3544 250444 3556
rect 250496 3544 250502 3596
rect 255866 3544 255872 3596
rect 255924 3584 255930 3596
rect 264330 3584 264336 3596
rect 255924 3556 264336 3584
rect 255924 3544 255930 3556
rect 264330 3544 264336 3556
rect 264388 3544 264394 3596
rect 270034 3544 270040 3596
rect 270092 3584 270098 3596
rect 287026 3584 287054 3624
rect 294598 3612 294604 3624
rect 294656 3612 294662 3664
rect 319714 3612 319720 3664
rect 319772 3652 319778 3664
rect 330478 3652 330484 3664
rect 319772 3624 330484 3652
rect 319772 3612 319778 3624
rect 330478 3612 330484 3624
rect 330536 3612 330542 3664
rect 341058 3612 341064 3664
rect 341116 3652 341122 3664
rect 356698 3652 356704 3664
rect 341116 3624 356704 3652
rect 341116 3612 341122 3624
rect 356698 3612 356704 3624
rect 356756 3612 356762 3664
rect 356808 3624 360976 3652
rect 270092 3556 287054 3584
rect 270092 3544 270098 3556
rect 292574 3544 292580 3596
rect 292632 3584 292638 3596
rect 294690 3584 294696 3596
rect 292632 3556 294696 3584
rect 292632 3544 292638 3556
rect 294690 3544 294696 3556
rect 294748 3544 294754 3596
rect 304258 3584 304264 3596
rect 296686 3556 304264 3584
rect 236748 3488 248414 3516
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 113818 3448 113824 3460
rect 624 3420 113824 3448
rect 624 3408 630 3420
rect 113818 3408 113824 3420
rect 113876 3408 113882 3460
rect 118694 3408 118700 3460
rect 118752 3448 118758 3460
rect 119890 3448 119896 3460
rect 118752 3420 119896 3448
rect 118752 3408 118758 3420
rect 119890 3408 119896 3420
rect 119948 3408 119954 3460
rect 168374 3408 168380 3460
rect 168432 3448 168438 3460
rect 169570 3448 169576 3460
rect 168432 3420 169576 3448
rect 168432 3408 168438 3420
rect 169570 3408 169576 3420
rect 169628 3408 169634 3460
rect 171106 3420 232176 3448
rect 69014 3340 69020 3392
rect 69072 3380 69078 3392
rect 69934 3380 69940 3392
rect 69072 3352 69940 3380
rect 69072 3340 69078 3352
rect 69934 3340 69940 3352
rect 69992 3340 69998 3392
rect 102134 3340 102140 3392
rect 102192 3380 102198 3392
rect 103330 3380 103336 3392
rect 102192 3352 103336 3380
rect 102192 3340 102198 3352
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 168374 3272 168380 3324
rect 168432 3312 168438 3324
rect 171106 3312 171134 3420
rect 168432 3284 171134 3312
rect 168432 3272 168438 3284
rect 229830 3272 229836 3324
rect 229888 3312 229894 3324
rect 231210 3312 231216 3324
rect 229888 3284 231216 3312
rect 229888 3272 229894 3284
rect 231210 3272 231216 3284
rect 231268 3272 231274 3324
rect 232148 3312 232176 3420
rect 232222 3340 232228 3392
rect 232280 3380 232286 3392
rect 236748 3380 236776 3488
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 254762 3516 254768 3528
rect 250036 3488 254768 3516
rect 250036 3476 250042 3488
rect 254762 3476 254768 3488
rect 254820 3476 254826 3528
rect 262950 3476 262956 3528
rect 263008 3516 263014 3528
rect 290458 3516 290464 3528
rect 263008 3488 290464 3516
rect 263008 3476 263014 3488
rect 290458 3476 290464 3488
rect 290516 3476 290522 3528
rect 291378 3476 291384 3528
rect 291436 3516 291442 3528
rect 296686 3516 296714 3556
rect 304258 3544 304264 3556
rect 304316 3544 304322 3596
rect 305546 3544 305552 3596
rect 305604 3584 305610 3596
rect 318150 3584 318156 3596
rect 305604 3556 318156 3584
rect 305604 3544 305610 3556
rect 318150 3544 318156 3556
rect 318208 3544 318214 3596
rect 330386 3544 330392 3596
rect 330444 3584 330450 3596
rect 330444 3556 345014 3584
rect 330444 3544 330450 3556
rect 291436 3488 296714 3516
rect 291436 3476 291442 3488
rect 297266 3476 297272 3528
rect 297324 3516 297330 3528
rect 298738 3516 298744 3528
rect 297324 3488 298744 3516
rect 297324 3476 297330 3488
rect 298738 3476 298744 3488
rect 298796 3476 298802 3528
rect 301958 3476 301964 3528
rect 302016 3516 302022 3528
rect 316678 3516 316684 3528
rect 302016 3488 316684 3516
rect 302016 3476 302022 3488
rect 316678 3476 316684 3488
rect 316736 3476 316742 3528
rect 323302 3476 323308 3528
rect 323360 3516 323366 3528
rect 337378 3516 337384 3528
rect 323360 3488 337384 3516
rect 323360 3476 323366 3488
rect 337378 3476 337384 3488
rect 337436 3476 337442 3528
rect 337470 3476 337476 3528
rect 337528 3516 337534 3528
rect 338758 3516 338764 3528
rect 337528 3488 338764 3516
rect 337528 3476 337534 3488
rect 338758 3476 338764 3488
rect 338816 3476 338822 3528
rect 340966 3476 340972 3528
rect 341024 3516 341030 3528
rect 342162 3516 342168 3528
rect 341024 3488 342168 3516
rect 341024 3476 341030 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 344986 3516 345014 3556
rect 348050 3544 348056 3596
rect 348108 3584 348114 3596
rect 348108 3556 354674 3584
rect 348108 3544 348114 3556
rect 348418 3516 348424 3528
rect 344986 3488 348424 3516
rect 348418 3476 348424 3488
rect 348476 3476 348482 3528
rect 349246 3476 349252 3528
rect 349304 3516 349310 3528
rect 350442 3516 350448 3528
rect 349304 3488 350448 3516
rect 349304 3476 349310 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 354646 3516 354674 3556
rect 355226 3544 355232 3596
rect 355284 3584 355290 3596
rect 356808 3584 356836 3624
rect 355284 3556 356836 3584
rect 355284 3544 355290 3556
rect 358722 3544 358728 3596
rect 358780 3584 358786 3596
rect 360838 3584 360844 3596
rect 358780 3556 360844 3584
rect 358780 3544 358786 3556
rect 360838 3544 360844 3556
rect 360896 3544 360902 3596
rect 360948 3584 360976 3624
rect 362310 3612 362316 3664
rect 362368 3652 362374 3664
rect 420914 3652 420920 3664
rect 362368 3624 420920 3652
rect 362368 3612 362374 3624
rect 420914 3612 420920 3624
rect 420972 3612 420978 3664
rect 439130 3612 439136 3664
rect 439188 3652 439194 3664
rect 440878 3652 440884 3664
rect 439188 3624 440884 3652
rect 439188 3612 439194 3624
rect 440878 3612 440884 3624
rect 440936 3612 440942 3664
rect 449802 3612 449808 3664
rect 449860 3652 449866 3664
rect 467098 3652 467104 3664
rect 449860 3624 467104 3652
rect 449860 3612 449866 3624
rect 467098 3612 467104 3624
rect 467156 3612 467162 3664
rect 467208 3624 468616 3652
rect 417050 3584 417056 3596
rect 360948 3556 417056 3584
rect 417050 3544 417056 3556
rect 417108 3544 417114 3596
rect 423766 3544 423772 3596
rect 423824 3584 423830 3596
rect 424962 3584 424968 3596
rect 423824 3556 424968 3584
rect 423824 3544 423830 3556
rect 424962 3544 424968 3556
rect 425020 3544 425026 3596
rect 426158 3544 426164 3596
rect 426216 3584 426222 3596
rect 441614 3584 441620 3596
rect 426216 3556 441620 3584
rect 426216 3544 426222 3556
rect 441614 3544 441620 3556
rect 441672 3544 441678 3596
rect 447778 3584 447784 3596
rect 444760 3556 447784 3584
rect 354646 3488 404768 3516
rect 302234 3448 302240 3460
rect 238726 3420 302240 3448
rect 232280 3352 236776 3380
rect 232280 3340 232286 3352
rect 237006 3340 237012 3392
rect 237064 3380 237070 3392
rect 238018 3380 238024 3392
rect 237064 3352 238024 3380
rect 237064 3340 237070 3352
rect 238018 3340 238024 3352
rect 238076 3340 238082 3392
rect 238726 3312 238754 3420
rect 302234 3408 302240 3420
rect 302292 3408 302298 3460
rect 309042 3408 309048 3460
rect 309100 3448 309106 3460
rect 311158 3448 311164 3460
rect 309100 3420 311164 3448
rect 309100 3408 309106 3420
rect 311158 3408 311164 3420
rect 311216 3408 311222 3460
rect 312630 3408 312636 3460
rect 312688 3448 312694 3460
rect 324958 3448 324964 3460
rect 312688 3420 324964 3448
rect 312688 3408 312694 3420
rect 324958 3408 324964 3420
rect 325016 3408 325022 3460
rect 333882 3408 333888 3460
rect 333940 3448 333946 3460
rect 404354 3448 404360 3460
rect 333940 3420 404360 3448
rect 333940 3408 333946 3420
rect 404354 3408 404360 3420
rect 404412 3408 404418 3460
rect 267734 3340 267740 3392
rect 267792 3380 267798 3392
rect 271230 3380 271236 3392
rect 267792 3352 271236 3380
rect 267792 3340 267798 3352
rect 271230 3340 271236 3352
rect 271288 3340 271294 3392
rect 281902 3340 281908 3392
rect 281960 3380 281966 3392
rect 285030 3380 285036 3392
rect 281960 3352 285036 3380
rect 281960 3340 281966 3352
rect 285030 3340 285036 3352
rect 285088 3340 285094 3392
rect 326798 3340 326804 3392
rect 326856 3380 326862 3392
rect 334710 3380 334716 3392
rect 326856 3352 334716 3380
rect 326856 3340 326862 3352
rect 334710 3340 334716 3352
rect 334768 3340 334774 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 404740 3380 404768 3488
rect 407114 3476 407120 3528
rect 407172 3516 407178 3528
rect 408402 3516 408408 3528
rect 407172 3488 408408 3516
rect 407172 3476 407178 3488
rect 408402 3476 408408 3488
rect 408460 3476 408466 3528
rect 411898 3476 411904 3528
rect 411956 3516 411962 3528
rect 444760 3516 444788 3556
rect 447778 3544 447784 3556
rect 447836 3544 447842 3596
rect 460934 3584 460940 3596
rect 447980 3556 460940 3584
rect 411956 3488 444788 3516
rect 411956 3476 411962 3488
rect 446214 3476 446220 3528
rect 446272 3516 446278 3528
rect 447870 3516 447876 3528
rect 446272 3488 447876 3516
rect 446272 3476 446278 3488
rect 447870 3476 447876 3488
rect 447928 3476 447934 3528
rect 404814 3408 404820 3460
rect 404872 3448 404878 3460
rect 446398 3448 446404 3460
rect 404872 3420 446404 3448
rect 404872 3408 404878 3420
rect 446398 3408 446404 3420
rect 446456 3408 446462 3460
rect 409874 3380 409880 3392
rect 404740 3352 409880 3380
rect 409874 3340 409880 3352
rect 409932 3340 409938 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 441614 3340 441620 3392
rect 441672 3380 441678 3392
rect 447980 3380 448008 3556
rect 460934 3544 460940 3556
rect 460992 3544 460998 3596
rect 461578 3544 461584 3596
rect 461636 3584 461642 3596
rect 467208 3584 467236 3624
rect 461636 3556 467236 3584
rect 461636 3544 461642 3556
rect 467466 3544 467472 3596
rect 467524 3584 467530 3596
rect 468478 3584 468484 3596
rect 467524 3556 468484 3584
rect 467524 3544 467530 3556
rect 468478 3544 468484 3556
rect 468536 3544 468542 3596
rect 468588 3584 468616 3624
rect 468662 3612 468668 3664
rect 468720 3652 468726 3664
rect 480898 3652 480904 3664
rect 468720 3624 480904 3652
rect 468720 3612 468726 3624
rect 480898 3612 480904 3624
rect 480956 3612 480962 3664
rect 525978 3612 525984 3664
rect 526036 3652 526042 3664
rect 533706 3652 533712 3664
rect 526036 3624 533712 3652
rect 526036 3612 526042 3624
rect 533706 3612 533712 3624
rect 533764 3612 533770 3664
rect 538186 3652 538214 3760
rect 543734 3748 543740 3800
rect 543792 3788 543798 3800
rect 563238 3788 563244 3800
rect 543792 3760 563244 3788
rect 543792 3748 543798 3760
rect 563238 3748 563244 3760
rect 563296 3748 563302 3800
rect 566458 3748 566464 3800
rect 566516 3788 566522 3800
rect 570322 3788 570328 3800
rect 566516 3760 570328 3788
rect 566516 3748 566522 3760
rect 570322 3748 570328 3760
rect 570380 3748 570386 3800
rect 547966 3680 547972 3732
rect 548024 3720 548030 3732
rect 568022 3720 568028 3732
rect 548024 3692 568028 3720
rect 548024 3680 548030 3692
rect 568022 3680 568028 3692
rect 568080 3680 568086 3732
rect 539594 3652 539600 3664
rect 538186 3624 539600 3652
rect 539594 3612 539600 3624
rect 539652 3612 539658 3664
rect 550634 3612 550640 3664
rect 550692 3652 550698 3664
rect 573910 3652 573916 3664
rect 550692 3624 573916 3652
rect 550692 3612 550698 3624
rect 573910 3612 573916 3624
rect 573968 3612 573974 3664
rect 468588 3556 472204 3584
rect 456794 3476 456800 3528
rect 456852 3516 456858 3528
rect 458082 3516 458088 3528
rect 456852 3488 458088 3516
rect 456852 3476 456858 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 471238 3516 471244 3528
rect 458284 3488 471244 3516
rect 450906 3408 450912 3460
rect 450964 3448 450970 3460
rect 450964 3420 451274 3448
rect 450964 3408 450970 3420
rect 441672 3352 448008 3380
rect 441672 3340 441678 3352
rect 232148 3284 238754 3312
rect 239306 3272 239312 3324
rect 239364 3312 239370 3324
rect 240870 3312 240876 3324
rect 239364 3284 240876 3312
rect 239364 3272 239370 3284
rect 240870 3272 240876 3284
rect 240928 3272 240934 3324
rect 253474 3272 253480 3324
rect 253532 3312 253538 3324
rect 258718 3312 258724 3324
rect 253532 3284 258724 3312
rect 253532 3272 253538 3284
rect 258718 3272 258724 3284
rect 258776 3272 258782 3324
rect 272426 3272 272432 3324
rect 272484 3312 272490 3324
rect 276750 3312 276756 3324
rect 272484 3284 276756 3312
rect 272484 3272 272490 3284
rect 276750 3272 276756 3284
rect 276808 3272 276814 3324
rect 451246 3312 451274 3420
rect 453298 3340 453304 3392
rect 453356 3380 453362 3392
rect 458284 3380 458312 3488
rect 471238 3476 471244 3488
rect 471296 3476 471302 3528
rect 472176 3516 472204 3556
rect 472250 3544 472256 3596
rect 472308 3584 472314 3596
rect 486418 3584 486424 3596
rect 472308 3556 486424 3584
rect 472308 3544 472314 3556
rect 486418 3544 486424 3556
rect 486476 3544 486482 3596
rect 493502 3544 493508 3596
rect 493560 3584 493566 3596
rect 500218 3584 500224 3596
rect 493560 3556 500224 3584
rect 493560 3544 493566 3556
rect 500218 3544 500224 3556
rect 500276 3544 500282 3596
rect 501782 3544 501788 3596
rect 501840 3584 501846 3596
rect 506750 3584 506756 3596
rect 501840 3556 506756 3584
rect 501840 3544 501846 3556
rect 506750 3544 506756 3556
rect 506808 3544 506814 3596
rect 508866 3544 508872 3596
rect 508924 3584 508930 3596
rect 510706 3584 510712 3596
rect 508924 3556 510712 3584
rect 508924 3544 508930 3556
rect 510706 3544 510712 3556
rect 510764 3544 510770 3596
rect 534166 3544 534172 3596
rect 534224 3584 534230 3596
rect 545482 3584 545488 3596
rect 534224 3556 545488 3584
rect 534224 3544 534230 3556
rect 545482 3544 545488 3556
rect 545540 3544 545546 3596
rect 549254 3544 549260 3596
rect 549312 3584 549318 3596
rect 571518 3584 571524 3596
rect 549312 3556 571524 3584
rect 549312 3544 549318 3556
rect 571518 3544 571524 3556
rect 571576 3544 571582 3596
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 576302 3584 576308 3596
rect 574796 3556 576308 3584
rect 574796 3544 574802 3556
rect 576302 3544 576308 3556
rect 576360 3544 576366 3596
rect 476758 3516 476764 3528
rect 472176 3488 476764 3516
rect 476758 3476 476764 3488
rect 476816 3476 476822 3528
rect 481726 3476 481732 3528
rect 481784 3516 481790 3528
rect 485038 3516 485044 3528
rect 481784 3488 485044 3516
rect 481784 3476 481790 3488
rect 485038 3476 485044 3488
rect 485096 3476 485102 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 508498 3516 508504 3528
rect 506532 3488 508504 3516
rect 506532 3476 506538 3488
rect 508498 3476 508504 3488
rect 508556 3476 508562 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 518986 3476 518992 3528
rect 519044 3516 519050 3528
rect 521838 3516 521844 3528
rect 519044 3488 521844 3516
rect 519044 3476 519050 3488
rect 521838 3476 521844 3488
rect 521896 3476 521902 3528
rect 524414 3476 524420 3528
rect 524472 3516 524478 3528
rect 531314 3516 531320 3528
rect 524472 3488 531320 3516
rect 524472 3476 524478 3488
rect 531314 3476 531320 3488
rect 531372 3476 531378 3528
rect 534074 3476 534080 3528
rect 534132 3516 534138 3528
rect 534132 3488 538214 3516
rect 534132 3476 534138 3488
rect 473998 3448 474004 3460
rect 453356 3352 458312 3380
rect 460906 3420 474004 3448
rect 453356 3340 453362 3352
rect 460906 3312 460934 3420
rect 473998 3408 474004 3420
rect 474056 3408 474062 3460
rect 486418 3408 486424 3460
rect 486476 3448 486482 3460
rect 496906 3448 496912 3460
rect 486476 3420 496912 3448
rect 486476 3408 486482 3420
rect 496906 3408 496912 3420
rect 496964 3408 496970 3460
rect 521654 3408 521660 3460
rect 521712 3448 521718 3460
rect 525426 3448 525432 3460
rect 521712 3420 525432 3448
rect 521712 3408 521718 3420
rect 525426 3408 525432 3420
rect 525484 3408 525490 3460
rect 527910 3408 527916 3460
rect 527968 3448 527974 3460
rect 536098 3448 536104 3460
rect 527968 3420 536104 3448
rect 527968 3408 527974 3420
rect 536098 3408 536104 3420
rect 536156 3408 536162 3460
rect 538186 3448 538214 3488
rect 538858 3476 538864 3528
rect 538916 3516 538922 3528
rect 541986 3516 541992 3528
rect 538916 3488 541992 3516
rect 538916 3476 538922 3488
rect 541986 3476 541992 3488
rect 542044 3476 542050 3528
rect 553394 3476 553400 3528
rect 553452 3516 553458 3528
rect 577406 3516 577412 3528
rect 553452 3488 577412 3516
rect 553452 3476 553458 3488
rect 577406 3476 577412 3488
rect 577464 3476 577470 3528
rect 578878 3476 578884 3528
rect 578936 3516 578942 3528
rect 580994 3516 581000 3528
rect 578936 3488 581000 3516
rect 578936 3476 578942 3488
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 546678 3448 546684 3460
rect 538186 3420 546684 3448
rect 546678 3408 546684 3420
rect 546736 3408 546742 3460
rect 553486 3408 553492 3460
rect 553544 3448 553550 3460
rect 578602 3448 578608 3460
rect 553544 3420 578608 3448
rect 553544 3408 553550 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 482830 3340 482836 3392
rect 482888 3380 482894 3392
rect 487798 3380 487804 3392
rect 482888 3352 487804 3380
rect 482888 3340 482894 3352
rect 487798 3340 487804 3352
rect 487856 3340 487862 3392
rect 538306 3340 538312 3392
rect 538364 3380 538370 3392
rect 552658 3380 552664 3392
rect 538364 3352 552664 3380
rect 538364 3340 538370 3352
rect 552658 3340 552664 3352
rect 552716 3340 552722 3392
rect 451246 3284 460934 3312
rect 558178 3272 558184 3324
rect 558236 3312 558242 3324
rect 559742 3312 559748 3324
rect 558236 3284 559748 3312
rect 558236 3272 558242 3284
rect 559742 3272 559748 3284
rect 559800 3272 559806 3324
rect 580258 3272 580264 3324
rect 580316 3312 580322 3324
rect 582190 3312 582196 3324
rect 580316 3284 582196 3312
rect 580316 3272 580322 3284
rect 582190 3272 582196 3284
rect 582248 3272 582254 3324
rect 242894 3204 242900 3256
rect 242952 3244 242958 3256
rect 247770 3244 247776 3256
rect 242952 3216 247776 3244
rect 242952 3204 242958 3216
rect 247770 3204 247776 3216
rect 247828 3204 247834 3256
rect 463970 3204 463976 3256
rect 464028 3244 464034 3256
rect 467190 3244 467196 3256
rect 464028 3216 467196 3244
rect 464028 3204 464034 3216
rect 467190 3204 467196 3216
rect 467248 3204 467254 3256
rect 517606 3204 517612 3256
rect 517664 3244 517670 3256
rect 519538 3244 519544 3256
rect 517664 3216 519544 3244
rect 517664 3204 517670 3216
rect 519538 3204 519544 3216
rect 519596 3204 519602 3256
rect 520458 3204 520464 3256
rect 520516 3244 520522 3256
rect 524230 3244 524236 3256
rect 520516 3216 524236 3244
rect 520516 3204 520522 3216
rect 524230 3204 524236 3216
rect 524288 3204 524294 3256
rect 369394 3136 369400 3188
rect 369452 3176 369458 3188
rect 370498 3176 370504 3188
rect 369452 3148 370504 3176
rect 369452 3136 369458 3148
rect 370498 3136 370504 3148
rect 370556 3136 370562 3188
rect 447410 3136 447416 3188
rect 447468 3176 447474 3188
rect 450538 3176 450544 3188
rect 447468 3148 450544 3176
rect 447468 3136 447474 3148
rect 450538 3136 450544 3148
rect 450596 3136 450602 3188
rect 512454 3136 512460 3188
rect 512512 3176 512518 3188
rect 513466 3176 513472 3188
rect 512512 3148 513472 3176
rect 512512 3136 512518 3148
rect 513466 3136 513472 3148
rect 513524 3136 513530 3188
rect 520366 3136 520372 3188
rect 520424 3176 520430 3188
rect 523034 3176 523040 3188
rect 520424 3148 523040 3176
rect 520424 3136 520430 3148
rect 523034 3136 523040 3148
rect 523092 3136 523098 3188
rect 524506 3136 524512 3188
rect 524564 3176 524570 3188
rect 530118 3176 530124 3188
rect 524564 3148 530124 3176
rect 524564 3136 524570 3148
rect 530118 3136 530124 3148
rect 530176 3136 530182 3188
rect 248782 3068 248788 3120
rect 248840 3108 248846 3120
rect 257338 3108 257344 3120
rect 248840 3080 257344 3108
rect 248840 3068 248846 3080
rect 257338 3068 257344 3080
rect 257396 3068 257402 3120
rect 279510 3000 279516 3052
rect 279568 3040 279574 3052
rect 280798 3040 280804 3052
rect 279568 3012 280804 3040
rect 279568 3000 279574 3012
rect 280798 3000 280804 3012
rect 280856 3000 280862 3052
rect 530578 3000 530584 3052
rect 530636 3040 530642 3052
rect 537202 3040 537208 3052
rect 530636 3012 537208 3040
rect 530636 3000 530642 3012
rect 537202 3000 537208 3012
rect 537260 3000 537266 3052
rect 433242 2932 433248 2984
rect 433300 2972 433306 2984
rect 434070 2972 434076 2984
rect 433300 2944 434076 2972
rect 433300 2932 433306 2944
rect 434070 2932 434076 2944
rect 434128 2932 434134 2984
rect 567838 2932 567844 2984
rect 567896 2972 567902 2984
rect 575106 2972 575112 2984
rect 567896 2944 575112 2972
rect 567896 2932 567902 2944
rect 575106 2932 575112 2944
rect 575164 2932 575170 2984
rect 264146 2864 264152 2916
rect 264204 2904 264210 2916
rect 268378 2904 268384 2916
rect 264204 2876 268384 2904
rect 264204 2864 264210 2876
rect 268378 2864 268384 2876
rect 268436 2864 268442 2916
rect 316034 960 316040 1012
rect 316092 1000 316098 1012
rect 317322 1000 317328 1012
rect 316092 972 317328 1000
rect 316092 960 316098 972
rect 317322 960 317328 972
rect 317380 960 317386 1012
<< via1 >>
rect 300124 700680 300176 700732
rect 356704 700680 356756 700732
rect 283840 700612 283892 700664
rect 344284 700612 344336 700664
rect 348792 700612 348844 700664
rect 396724 700612 396776 700664
rect 332508 700544 332560 700596
rect 405004 700544 405056 700596
rect 170312 700476 170364 700528
rect 177304 700476 177356 700528
rect 267648 700476 267700 700528
rect 351184 700476 351236 700528
rect 137836 700408 137888 700460
rect 184204 700408 184256 700460
rect 235172 700408 235224 700460
rect 358084 700408 358136 700460
rect 408408 700408 408460 700460
rect 429844 700408 429896 700460
rect 72976 700340 73028 700392
rect 186964 700340 187016 700392
rect 218980 700340 219032 700392
rect 348424 700340 348476 700392
rect 409788 700340 409840 700392
rect 462320 700340 462372 700392
rect 527180 700340 527232 700392
rect 546684 700340 546736 700392
rect 8116 700272 8168 700324
rect 188344 700272 188396 700324
rect 202788 700272 202840 700324
rect 353944 700272 353996 700324
rect 364984 700272 365036 700324
rect 393964 700272 394016 700324
rect 408316 700272 408368 700324
rect 478512 700272 478564 700324
rect 494796 700272 494848 700324
rect 546776 700272 546828 700324
rect 548524 700272 548576 700324
rect 559656 700272 559708 700324
rect 409696 699660 409748 699712
rect 413652 699660 413704 699712
rect 543464 699660 543516 699712
rect 547880 699660 547932 699712
rect 105452 698912 105504 698964
rect 407764 698912 407816 698964
rect 577504 696940 577556 696992
rect 580448 696940 580500 696992
rect 3424 683136 3476 683188
rect 178776 683136 178828 683188
rect 28724 674976 28776 675028
rect 28632 674908 28684 674960
rect 34520 674908 34572 674960
rect 46204 674908 46256 674960
rect 28816 674840 28868 674892
rect 46940 674840 46992 674892
rect 570604 670692 570656 670744
rect 580172 670692 580224 670744
rect 340144 660288 340196 660340
rect 488908 660288 488960 660340
rect 246304 659676 246356 659728
rect 337108 659676 337160 659728
rect 408224 659676 408276 659728
rect 499856 659676 499908 659728
rect 560944 643084 560996 643136
rect 580172 643084 580224 643136
rect 2964 618264 3016 618316
rect 21364 618264 21416 618316
rect 567844 616836 567896 616888
rect 580172 616836 580224 616888
rect 339408 612008 339460 612060
rect 407120 612008 407172 612060
rect 339408 610580 339460 610632
rect 407120 610580 407172 610632
rect 338304 608608 338356 608660
rect 407120 608608 407172 608660
rect 338120 607180 338172 607232
rect 407120 607180 407172 607232
rect 338396 605820 338448 605872
rect 407120 605820 407172 605872
rect 338212 604460 338264 604512
rect 339408 604460 339460 604512
rect 407120 604460 407172 604512
rect 339224 603712 339276 603764
rect 407120 603712 407172 603764
rect 574744 590656 574796 590708
rect 580172 590656 580224 590708
rect 99196 587392 99248 587444
rect 170864 587392 170916 587444
rect 149520 587324 149572 587376
rect 171600 587324 171652 587376
rect 143448 587256 143500 587308
rect 167000 587256 167052 587308
rect 142712 587188 142764 587240
rect 168104 587188 168156 587240
rect 140136 587120 140188 587172
rect 168012 587120 168064 587172
rect 137928 587052 137980 587104
rect 167828 587052 167880 587104
rect 139032 586984 139084 587036
rect 171416 586984 171468 587036
rect 136548 586916 136600 586968
rect 169760 586916 169812 586968
rect 133144 586848 133196 586900
rect 167920 586848 167972 586900
rect 129648 586780 129700 586832
rect 172796 586780 172848 586832
rect 126888 586712 126940 586764
rect 173532 586712 173584 586764
rect 100576 586644 100628 586696
rect 170772 586644 170824 586696
rect 28540 586576 28592 586628
rect 43076 586576 43128 586628
rect 103152 586576 103204 586628
rect 174636 586576 174688 586628
rect 28448 586508 28500 586560
rect 43536 586508 43588 586560
rect 150716 586508 150768 586560
rect 167092 586508 167144 586560
rect 139308 585828 139360 585880
rect 181536 585828 181588 585880
rect 105084 585760 105136 585812
rect 174728 585760 174780 585812
rect 339224 585760 339276 585812
rect 407120 585760 407172 585812
rect 130568 585080 130620 585132
rect 172888 585080 172940 585132
rect 120540 585012 120592 585064
rect 167184 585012 167236 585064
rect 125048 584944 125100 584996
rect 175372 584944 175424 584996
rect 129372 584876 129424 584928
rect 180800 584876 180852 584928
rect 122656 584808 122708 584860
rect 178040 584808 178092 584860
rect 117136 584740 117188 584792
rect 172520 584740 172572 584792
rect 114836 584672 114888 584724
rect 171232 584672 171284 584724
rect 113824 584604 113876 584656
rect 172612 584604 172664 584656
rect 109500 584536 109552 584588
rect 171324 584536 171376 584588
rect 110512 584468 110564 584520
rect 187148 584468 187200 584520
rect 62948 584400 63000 584452
rect 196900 584400 196952 584452
rect 131120 584332 131172 584384
rect 173256 584332 173308 584384
rect 136456 584264 136508 584316
rect 167644 584264 167696 584316
rect 147680 584196 147732 584248
rect 171508 584196 171560 584248
rect 132592 582972 132644 583024
rect 178960 582972 179012 583024
rect 339408 582972 339460 583024
rect 407120 582972 407172 583024
rect 122840 581680 122892 581732
rect 180064 581680 180116 581732
rect 95240 581612 95292 581664
rect 185676 581612 185728 581664
rect 64880 580252 64932 580304
rect 189816 580252 189868 580304
rect 3148 579640 3200 579692
rect 181444 579640 181496 579692
rect 120172 578960 120224 579012
rect 191196 578960 191248 579012
rect 83832 578892 83884 578944
rect 194048 578892 194100 578944
rect 114560 577532 114612 577584
rect 184296 577532 184348 577584
rect 86408 577464 86460 577516
rect 195428 577464 195480 577516
rect 565084 576852 565136 576904
rect 580172 576852 580224 576904
rect 113088 576172 113140 576224
rect 177488 576172 177540 576224
rect 93768 576104 93820 576156
rect 196808 576104 196860 576156
rect 338028 575492 338080 575544
rect 425060 575492 425112 575544
rect 330208 575424 330260 575476
rect 337108 575424 337160 575476
rect 408224 575424 408276 575476
rect 415400 575424 415452 575476
rect 199384 575152 199436 575204
rect 293960 575152 294012 575204
rect 195704 575084 195756 575136
rect 289820 575084 289872 575136
rect 198648 575016 198700 575068
rect 293960 575016 294012 575068
rect 301872 575016 301924 575068
rect 342352 575016 342404 575068
rect 199844 574948 199896 575000
rect 280160 574948 280212 575000
rect 320456 574948 320508 575000
rect 330484 574948 330536 575000
rect 340144 574948 340196 575000
rect 466460 574948 466512 575000
rect 195888 574880 195940 574932
rect 280252 574880 280304 574932
rect 307576 574880 307628 574932
rect 339592 574880 339644 574932
rect 409420 574880 409472 574932
rect 426440 574880 426492 574932
rect 118608 574812 118660 574864
rect 188436 574812 188488 574864
rect 197084 574812 197136 574864
rect 281540 574812 281592 574864
rect 304632 574812 304684 574864
rect 336832 574812 336884 574864
rect 409512 574812 409564 574864
rect 437480 574812 437532 574864
rect 81348 574744 81400 574796
rect 191288 574744 191340 574796
rect 197176 574744 197228 574796
rect 284300 574744 284352 574796
rect 305552 574744 305604 574796
rect 339684 574744 339736 574796
rect 406568 574744 406620 574796
rect 438860 574744 438912 574796
rect 195612 574676 195664 574728
rect 284392 574676 284444 574728
rect 306288 574676 306340 574728
rect 339776 574676 339828 574728
rect 406476 574676 406528 574728
rect 444380 574676 444432 574728
rect 285312 574608 285364 574660
rect 339960 574608 340012 574660
rect 409236 574608 409288 574660
rect 451280 574608 451332 574660
rect 195796 574540 195848 574592
rect 287520 574540 287572 574592
rect 302884 574540 302936 574592
rect 337476 574540 337528 574592
rect 405280 574540 405332 574592
rect 448520 574540 448572 574592
rect 287888 574472 287940 574524
rect 341432 574472 341484 574524
rect 405096 574472 405148 574524
rect 451280 574472 451332 574524
rect 490564 574472 490616 574524
rect 492680 574472 492732 574524
rect 198556 574404 198608 574456
rect 291200 574404 291252 574456
rect 300676 574404 300728 574456
rect 342444 574404 342496 574456
rect 406384 574404 406436 574456
rect 455420 574404 455472 574456
rect 199752 574336 199804 574388
rect 292580 574336 292632 574388
rect 297916 574336 297968 574388
rect 340972 574336 341024 574388
rect 400864 574336 400916 574388
rect 458180 574336 458232 574388
rect 284208 574268 284260 574320
rect 342260 574268 342312 574320
rect 398104 574268 398156 574320
rect 462872 574268 462924 574320
rect 480904 574268 480956 574320
rect 492680 574268 492732 574320
rect 196716 574200 196768 574252
rect 288440 574200 288492 574252
rect 292488 574200 292540 574252
rect 339500 574200 339552 574252
rect 396816 574200 396868 574252
rect 465080 574200 465132 574252
rect 487804 574200 487856 574252
rect 492772 574200 492824 574252
rect 196992 574132 197044 574184
rect 285680 574132 285732 574184
rect 286600 574132 286652 574184
rect 341524 574132 341576 574184
rect 391204 574132 391256 574184
rect 459560 574132 459612 574184
rect 485044 574132 485096 574184
rect 492956 574132 493008 574184
rect 195520 574064 195572 574116
rect 306472 574064 306524 574116
rect 68928 573384 68980 573436
rect 177580 573384 177632 573436
rect 191748 573384 191800 573436
rect 269120 573384 269172 573436
rect 360200 573384 360252 573436
rect 447140 573384 447192 573436
rect 3608 573316 3660 573368
rect 407856 573316 407908 573368
rect 199568 572636 199620 572688
rect 276020 572636 276072 572688
rect 291016 572636 291068 572688
rect 337108 572636 337160 572688
rect 402244 572636 402296 572688
rect 443092 572636 443144 572688
rect 198464 572568 198516 572620
rect 277676 572568 277728 572620
rect 291108 572568 291160 572620
rect 337200 572568 337252 572620
rect 402428 572568 402480 572620
rect 445852 572568 445904 572620
rect 196624 572500 196676 572552
rect 278780 572500 278832 572552
rect 289728 572500 289780 572552
rect 337292 572500 337344 572552
rect 402704 572500 402756 572552
rect 447232 572500 447284 572552
rect 193036 572432 193088 572484
rect 295340 572432 295392 572484
rect 296536 572432 296588 572484
rect 340880 572432 340932 572484
rect 402336 572432 402388 572484
rect 449992 572432 450044 572484
rect 194416 572364 194468 572416
rect 298100 572364 298152 572416
rect 299204 572364 299256 572416
rect 341340 572364 341392 572416
rect 402612 572364 402664 572416
rect 452660 572364 452712 572416
rect 194324 572296 194376 572348
rect 299480 572296 299532 572348
rect 399760 572296 399812 572348
rect 454132 572296 454184 572348
rect 192944 572228 192996 572280
rect 298192 572228 298244 572280
rect 298928 572228 298980 572280
rect 342536 572228 342588 572280
rect 399576 572228 399628 572280
rect 456892 572228 456944 572280
rect 194508 572160 194560 572212
rect 302240 572160 302292 572212
rect 399668 572160 399720 572212
rect 459284 572160 459336 572212
rect 193128 572092 193180 572144
rect 300860 572092 300912 572144
rect 399944 572092 399996 572144
rect 461308 572092 461360 572144
rect 192760 572024 192812 572076
rect 303620 572024 303672 572076
rect 399484 572024 399536 572076
rect 463792 572024 463844 572076
rect 71688 571956 71740 572008
rect 182916 571956 182968 572008
rect 194140 571956 194192 572008
rect 305000 571956 305052 572008
rect 399852 571956 399904 572008
rect 466460 571956 466512 572008
rect 199476 571888 199528 571940
rect 274640 571888 274692 571940
rect 293776 571888 293828 571940
rect 338580 571888 338632 571940
rect 402520 571888 402572 571940
rect 441804 571888 441856 571940
rect 199660 571820 199712 571872
rect 273260 571820 273312 571872
rect 294696 571820 294748 571872
rect 339868 571820 339920 571872
rect 405464 571820 405516 571872
rect 440332 571820 440384 571872
rect 405648 571752 405700 571804
rect 436192 571752 436244 571804
rect 125508 570664 125560 570716
rect 193956 570664 194008 570716
rect 88248 570596 88300 570648
rect 181628 570596 181680 570648
rect 237196 570596 237248 570648
rect 344376 570596 344428 570648
rect 365260 570596 365312 570648
rect 452752 570596 452804 570648
rect 128268 569440 128320 569492
rect 195336 569440 195388 569492
rect 194232 569372 194284 569424
rect 270500 569372 270552 569424
rect 191656 569304 191708 569356
rect 269212 569304 269264 569356
rect 192852 569236 192904 569288
rect 271880 569236 271932 569288
rect 91008 569168 91060 569220
rect 192484 569168 192536 569220
rect 253756 569168 253808 569220
rect 347044 569168 347096 569220
rect 367744 569168 367796 569220
rect 455512 569168 455564 569220
rect 131028 567876 131080 567928
rect 167736 567876 167788 567928
rect 108948 567808 109000 567860
rect 176200 567808 176252 567860
rect 253112 567808 253164 567860
rect 347136 567808 347188 567860
rect 374000 567808 374052 567860
rect 461124 567808 461176 567860
rect 74448 566448 74500 566500
rect 184480 566448 184532 566500
rect 356428 566448 356480 566500
rect 444472 566448 444524 566500
rect 3424 565836 3476 565888
rect 400956 565836 401008 565888
rect 75828 565156 75880 565208
rect 188528 565156 188580 565208
rect 3516 565088 3568 565140
rect 408040 565088 408092 565140
rect 142068 563796 142120 563848
rect 168196 563796 168248 563848
rect 78588 563728 78640 563780
rect 170956 563728 171008 563780
rect 357716 563728 357768 563780
rect 444564 563728 444616 563780
rect 3792 563660 3844 563712
rect 408132 563660 408184 563712
rect 29736 563116 29788 563168
rect 29644 563048 29696 563100
rect 35716 563048 35768 563100
rect 46756 563048 46808 563100
rect 566464 563048 566516 563100
rect 580172 563048 580224 563100
rect 28724 562572 28776 562624
rect 29736 562572 29788 562624
rect 28816 562300 28868 562352
rect 29828 562300 29880 562352
rect 48044 562300 48096 562352
rect 60648 562300 60700 562352
rect 179052 562300 179104 562352
rect 253848 562300 253900 562352
rect 348516 562300 348568 562352
rect 351368 562300 351420 562352
rect 438952 562300 439004 562352
rect 28632 561960 28684 562012
rect 29644 561960 29696 562012
rect 375288 560940 375340 560992
rect 462412 560940 462464 560992
rect 377772 559512 377824 559564
rect 464344 559512 464396 559564
rect 379060 558152 379112 558204
rect 466644 558152 466696 558204
rect 355140 556792 355192 556844
rect 443000 556792 443052 556844
rect 381544 555432 381596 555484
rect 468484 555432 468536 555484
rect 380348 554004 380400 554056
rect 467840 554004 467892 554056
rect 3424 553392 3476 553444
rect 28264 553392 28316 553444
rect 376576 552644 376628 552696
rect 463700 552644 463752 552696
rect 369032 551284 369084 551336
rect 455604 551284 455656 551336
rect 348516 550536 348568 550588
rect 485044 550536 485096 550588
rect 347136 549176 347188 549228
rect 347596 549176 347648 549228
rect 487804 549176 487856 549228
rect 347044 547816 347096 547868
rect 490564 547816 490616 547868
rect 346400 546456 346452 546508
rect 347044 546456 347096 546508
rect 254584 545708 254636 545760
rect 345112 545708 345164 545760
rect 480904 545708 480956 545760
rect 343824 545028 343876 545080
rect 344376 545028 344428 545080
rect 507952 545028 508004 545080
rect 238576 544348 238628 544400
rect 342628 544348 342680 544400
rect 342628 543668 342680 543720
rect 506480 543668 506532 543720
rect 238668 542988 238720 543040
rect 341616 542988 341668 543040
rect 358912 541696 358964 541748
rect 445760 541696 445812 541748
rect 361488 541628 361540 541680
rect 448612 541628 448664 541680
rect 384120 540812 384172 540864
rect 470692 540812 470744 540864
rect 385316 540744 385368 540796
rect 471980 540744 472032 540796
rect 386604 540676 386656 540728
rect 473360 540676 473412 540728
rect 387892 540608 387944 540660
rect 474740 540608 474792 540660
rect 389088 540540 389140 540592
rect 476120 540540 476172 540592
rect 352656 540472 352708 540524
rect 440240 540472 440292 540524
rect 280068 540404 280120 540456
rect 338764 540404 338816 540456
rect 382832 540404 382884 540456
rect 470600 540404 470652 540456
rect 278688 540336 278740 540388
rect 338672 540336 338724 540388
rect 353300 540336 353352 540388
rect 441620 540336 441672 540388
rect 218060 540268 218112 540320
rect 527180 540268 527232 540320
rect 217600 540200 217652 540252
rect 528836 540200 528888 540252
rect 187056 539928 187108 539980
rect 205732 539928 205784 539980
rect 190368 539860 190420 539912
rect 218060 539860 218112 539912
rect 169300 539792 169352 539844
rect 338856 539792 338908 539844
rect 169208 539724 169260 539776
rect 340052 539724 340104 539776
rect 169116 539656 169168 539708
rect 340328 539656 340380 539708
rect 169024 539588 169076 539640
rect 340236 539588 340288 539640
rect 370228 539316 370280 539368
rect 456800 539316 456852 539368
rect 371516 539248 371568 539300
rect 458364 539248 458416 539300
rect 372804 539180 372856 539232
rect 459652 539180 459704 539232
rect 362684 539112 362736 539164
rect 449900 539112 449952 539164
rect 318708 539044 318760 539096
rect 342720 539044 342772 539096
rect 363972 539044 364024 539096
rect 451280 539044 451332 539096
rect 284208 538976 284260 539028
rect 342812 538976 342864 539028
rect 350172 538976 350224 539028
rect 437572 538976 437624 539028
rect 282828 538908 282880 538960
rect 342904 538908 342956 538960
rect 366456 538908 366508 538960
rect 454040 538908 454092 538960
rect 281448 538840 281500 538892
rect 341708 538840 341760 538892
rect 407672 538840 407724 538892
rect 540796 538840 540848 538892
rect 570696 524424 570748 524476
rect 580172 524424 580224 524476
rect 3516 514768 3568 514820
rect 18604 514768 18656 514820
rect 565176 510620 565228 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 28724 500964 28776 501016
rect 339316 491240 339368 491292
rect 340328 491240 340380 491292
rect 407212 491240 407264 491292
rect 339408 491172 339460 491224
rect 340236 491172 340288 491224
rect 407120 491172 407172 491224
rect 340052 488452 340104 488504
rect 407120 488452 407172 488504
rect 169668 487092 169720 487144
rect 187056 487092 187108 487144
rect 338856 487092 338908 487144
rect 407120 487092 407172 487144
rect 168840 486412 168892 486464
rect 178684 486412 178736 486464
rect 339408 484372 339460 484424
rect 340236 484372 340288 484424
rect 407120 484372 407172 484424
rect 577596 484372 577648 484424
rect 580632 484372 580684 484424
rect 340052 483012 340104 483064
rect 407120 483012 407172 483064
rect 338856 481652 338908 481704
rect 407120 481652 407172 481704
rect 165528 476076 165580 476128
rect 167184 476076 167236 476128
rect 3516 475532 3568 475584
rect 166724 475532 166776 475584
rect 28540 475464 28592 475516
rect 42800 475464 42852 475516
rect 151360 475396 151412 475448
rect 151728 475396 151780 475448
rect 167092 475396 167144 475448
rect 29644 475328 29696 475380
rect 34520 475328 34572 475380
rect 28448 475260 28500 475312
rect 42800 475328 42852 475380
rect 141792 475328 141844 475380
rect 175924 475328 175976 475380
rect 129648 475260 129700 475312
rect 173900 475260 173952 475312
rect 174912 475260 174964 475312
rect 126888 475192 126940 475244
rect 176660 475192 176712 475244
rect 131028 475124 131080 475176
rect 181904 475124 181956 475176
rect 128268 475056 128320 475108
rect 187700 475056 187752 475108
rect 115480 474988 115532 475040
rect 175280 474988 175332 475040
rect 110328 474920 110380 474972
rect 171784 474920 171836 474972
rect 172428 474920 172480 474972
rect 121184 474852 121236 474904
rect 129004 474852 129056 474904
rect 129556 474852 129608 474904
rect 193864 474852 193916 474904
rect 60648 474784 60700 474836
rect 167552 474784 167604 474836
rect 175924 474784 175976 474836
rect 199200 474784 199252 474836
rect 121368 474716 121420 474768
rect 126244 474716 126296 474768
rect 174912 474716 174964 474768
rect 199292 474716 199344 474768
rect 28448 474648 28500 474700
rect 29644 474648 29696 474700
rect 136548 474172 136600 474224
rect 137284 474172 137336 474224
rect 139308 474104 139360 474156
rect 181720 474104 181772 474156
rect 136364 474036 136416 474088
rect 192576 474036 192628 474088
rect 96528 473968 96580 474020
rect 179144 473968 179196 474020
rect 143356 472744 143408 472796
rect 177396 472744 177448 472796
rect 133696 472676 133748 472728
rect 191380 472676 191432 472728
rect 93768 472608 93820 472660
rect 180156 472608 180208 472660
rect 177396 471996 177448 472048
rect 195244 471996 195296 472048
rect 131028 471384 131080 471436
rect 189908 471384 189960 471436
rect 112996 471316 113048 471368
rect 180248 471316 180300 471368
rect 86868 471248 86920 471300
rect 183100 471248 183152 471300
rect 566556 470568 566608 470620
rect 580172 470568 580224 470620
rect 124036 469956 124088 470008
rect 174820 469956 174872 470008
rect 111616 469888 111668 469940
rect 191472 469888 191524 469940
rect 84108 469820 84160 469872
rect 185860 469820 185912 469872
rect 121276 468596 121328 468648
rect 192668 468596 192720 468648
rect 108856 468528 108908 468580
rect 187240 468528 187292 468580
rect 75828 468460 75880 468512
rect 193772 468460 193824 468512
rect 115756 467236 115808 467288
rect 176292 467236 176344 467288
rect 106188 467168 106240 467220
rect 184664 467168 184716 467220
rect 78588 467100 78640 467152
rect 195152 467100 195204 467152
rect 74448 465672 74500 465724
rect 177764 465672 177816 465724
rect 136548 464448 136600 464500
rect 169852 464448 169904 464500
rect 100668 464380 100720 464432
rect 177672 464380 177724 464432
rect 68928 464312 68980 464364
rect 187424 464312 187476 464364
rect 169852 463700 169904 463752
rect 170404 463700 170456 463752
rect 176476 463700 176528 463752
rect 339408 463700 339460 463752
rect 340328 463700 340380 463752
rect 407120 463700 407172 463752
rect 339132 462952 339184 463004
rect 407120 462952 407172 463004
rect 407672 462952 407724 463004
rect 3516 462340 3568 462392
rect 191564 462340 191616 462392
rect 103428 461660 103480 461712
rect 188620 461660 188672 461712
rect 81348 461592 81400 461644
rect 190000 461592 190052 461644
rect 339040 461592 339092 461644
rect 407120 461592 407172 461644
rect 128268 460232 128320 460284
rect 183008 460232 183060 460284
rect 88248 460164 88300 460216
rect 174912 460164 174964 460216
rect 118516 458872 118568 458924
rect 185768 458872 185820 458924
rect 91008 458804 91060 458856
rect 176384 458804 176436 458856
rect 195060 457716 195112 457768
rect 195520 457716 195572 457768
rect 195244 457580 195296 457632
rect 195520 457580 195572 457632
rect 125508 457512 125560 457564
rect 168288 457512 168340 457564
rect 99288 457444 99340 457496
rect 181812 457444 181864 457496
rect 561036 456764 561088 456816
rect 580172 456764 580224 456816
rect 135168 456696 135220 456748
rect 168748 456696 168800 456748
rect 197084 456152 197136 456204
rect 137928 456084 137980 456136
rect 172428 456084 172480 456136
rect 63408 456016 63460 456068
rect 188712 456016 188764 456068
rect 197176 455948 197228 456000
rect 171876 455472 171928 455524
rect 172428 455472 172480 455524
rect 195244 455472 195296 455524
rect 168748 455404 168800 455456
rect 196072 455404 196124 455456
rect 169852 455336 169904 455388
rect 171048 455336 171100 455388
rect 171600 455336 171652 455388
rect 150348 454928 150400 454980
rect 169852 454928 169904 454980
rect 148324 454860 148376 454912
rect 183468 454860 183520 454912
rect 113088 454792 113140 454844
rect 172428 454792 172480 454844
rect 114376 454724 114428 454776
rect 176108 454724 176160 454776
rect 71688 454656 71740 454708
rect 184756 454656 184808 454708
rect 183192 454180 183244 454232
rect 183468 454180 183520 454232
rect 197360 454180 197412 454232
rect 176108 454112 176160 454164
rect 198740 454112 198792 454164
rect 172060 454044 172112 454096
rect 172428 454044 172480 454096
rect 195980 454044 196032 454096
rect 193588 453976 193640 454028
rect 193864 453976 193916 454028
rect 143448 453908 143500 453960
rect 176016 453908 176068 453960
rect 129004 453840 129056 453892
rect 172704 453840 172756 453892
rect 336280 453840 336332 453892
rect 336924 453840 336976 453892
rect 126244 453772 126296 453824
rect 173440 453772 173492 453824
rect 122748 453704 122800 453756
rect 169852 453704 169904 453756
rect 291016 453704 291068 453756
rect 338672 453704 338724 453756
rect 124128 453636 124180 453688
rect 179420 453636 179472 453688
rect 289820 453636 289872 453688
rect 338764 453636 338816 453688
rect 117228 453568 117280 453620
rect 174084 453568 174136 453620
rect 324964 453568 325016 453620
rect 399944 453568 399996 453620
rect 132408 453500 132460 453552
rect 191104 453500 191156 453552
rect 278044 453500 278096 453552
rect 311164 453500 311216 453552
rect 405280 453500 405332 453552
rect 114468 453432 114520 453484
rect 174544 453432 174596 453484
rect 118608 453364 118660 453416
rect 185952 453364 186004 453416
rect 281448 453432 281500 453484
rect 301228 453432 301280 453484
rect 406568 453432 406620 453484
rect 196164 453364 196216 453416
rect 294788 453364 294840 453416
rect 298560 453364 298612 453416
rect 405648 453364 405700 453416
rect 119988 453296 120040 453348
rect 189724 453296 189776 453348
rect 288900 453296 288952 453348
rect 299848 453296 299900 453348
rect 409512 453296 409564 453348
rect 409696 453296 409748 453348
rect 468300 453296 468352 453348
rect 199292 453228 199344 453280
rect 298468 453228 298520 453280
rect 193588 453160 193640 453212
rect 299572 453160 299624 453212
rect 174544 453092 174596 453144
rect 284300 453092 284352 453144
rect 199200 453024 199252 453076
rect 311072 453024 311124 453076
rect 174084 452956 174136 453008
rect 286784 452956 286836 453008
rect 179420 452888 179472 452940
rect 293684 452888 293736 452940
rect 172704 452820 172756 452872
rect 290188 452820 290240 452872
rect 173440 452752 173492 452804
rect 291200 452752 291252 452804
rect 169852 452684 169904 452736
rect 170680 452684 170732 452736
rect 292580 452684 292632 452736
rect 335084 452684 335136 452736
rect 337384 452684 337436 452736
rect 176016 452616 176068 452668
rect 312360 452616 312412 452668
rect 29552 452548 29604 452600
rect 29736 452548 29788 452600
rect 140688 452548 140740 452600
rect 167276 452548 167328 452600
rect 176476 452548 176528 452600
rect 305276 452548 305328 452600
rect 195520 452480 195572 452532
rect 313372 452480 313424 452532
rect 330024 452480 330076 452532
rect 399852 452480 399904 452532
rect 466184 452480 466236 452532
rect 467104 452480 467156 452532
rect 473544 452480 473596 452532
rect 476764 452480 476816 452532
rect 481088 452480 481140 452532
rect 485136 452480 485188 452532
rect 493600 452480 493652 452532
rect 497464 452480 497516 452532
rect 503536 452480 503588 452532
rect 504364 452480 504416 452532
rect 505928 452480 505980 452532
rect 507124 452480 507176 452532
rect 197360 452412 197412 452464
rect 314660 452412 314712 452464
rect 317420 452412 317472 452464
rect 399760 452412 399812 452464
rect 483480 452412 483532 452464
rect 487804 452412 487856 452464
rect 195244 452344 195296 452396
rect 307852 452344 307904 452396
rect 316224 452344 316276 452396
rect 402612 452344 402664 452396
rect 196072 452276 196124 452328
rect 304172 452276 304224 452328
rect 312452 452276 312504 452328
rect 402336 452276 402388 452328
rect 151728 452208 151780 452260
rect 169944 452208 169996 452260
rect 195980 452208 196032 452260
rect 282092 452208 282144 452260
rect 309968 452208 310020 452260
rect 402704 452208 402756 452260
rect 139216 452140 139268 452192
rect 171968 452140 172020 452192
rect 198740 452140 198792 452192
rect 283196 452140 283248 452192
rect 308680 452140 308732 452192
rect 402428 452140 402480 452192
rect 137284 452072 137336 452124
rect 170496 452072 170548 452124
rect 278044 452072 278096 452124
rect 301964 452072 302016 452124
rect 306104 452072 306156 452124
rect 402244 452072 402296 452124
rect 133788 452004 133840 452056
rect 187056 452004 187108 452056
rect 303620 452004 303672 452056
rect 402520 452004 402572 452056
rect 28540 451936 28592 451988
rect 34520 451936 34572 451988
rect 66168 451936 66220 451988
rect 175004 451936 175056 451988
rect 302332 451936 302384 451988
rect 405464 451936 405516 451988
rect 29552 451868 29604 451920
rect 45652 451868 45704 451920
rect 167276 451868 167328 451920
rect 309876 451868 309928 451920
rect 320180 451868 320232 451920
rect 425428 451868 425480 451920
rect 280988 451800 281040 451852
rect 341432 451800 341484 451852
rect 282276 451732 282328 451784
rect 341524 451732 341576 451784
rect 283472 451664 283524 451716
rect 339960 451664 340012 451716
rect 195060 451596 195112 451648
rect 201776 451596 201828 451648
rect 198372 451528 198424 451580
rect 200212 451528 200264 451580
rect 187056 451460 187108 451512
rect 303068 451460 303120 451512
rect 171968 451392 172020 451444
rect 308956 451392 309008 451444
rect 170496 451324 170548 451376
rect 306380 451324 306432 451376
rect 318800 451324 318852 451376
rect 319444 451324 319496 451376
rect 426900 451324 426952 451376
rect 495992 451324 496044 451376
rect 530584 451324 530636 451376
rect 169944 451256 169996 451308
rect 320180 451256 320232 451308
rect 468668 451256 468720 451308
rect 474004 451256 474056 451308
rect 476028 451256 476080 451308
rect 480904 451256 480956 451308
rect 29828 451188 29880 451240
rect 48044 451188 48096 451240
rect 170312 451188 170364 451240
rect 452844 451188 452896 451240
rect 173808 451120 173860 451172
rect 450268 451120 450320 451172
rect 169300 451052 169352 451104
rect 340236 451052 340288 451104
rect 194140 450916 194192 450968
rect 203064 450916 203116 450968
rect 168012 450848 168064 450900
rect 193680 450848 193732 450900
rect 436284 450848 436336 450900
rect 168196 450780 168248 450832
rect 187332 450780 187384 450832
rect 434720 450780 434772 450832
rect 168104 450712 168156 450764
rect 179236 450712 179288 450764
rect 433708 450712 433760 450764
rect 165528 450644 165580 450696
rect 184572 450644 184624 450696
rect 454132 450644 454184 450696
rect 516048 450644 516100 450696
rect 556344 450644 556396 450696
rect 28724 450576 28776 450628
rect 429384 450576 429436 450628
rect 443644 450576 443696 450628
rect 519912 450576 519964 450628
rect 18604 450508 18656 450560
rect 430580 450508 430632 450560
rect 438676 450508 438728 450560
rect 517336 450508 517388 450560
rect 169300 450168 169352 450220
rect 169484 450168 169536 450220
rect 28356 450100 28408 450152
rect 421840 450100 421892 450152
rect 28448 450032 28500 450084
rect 423036 450032 423088 450084
rect 3332 449964 3384 450016
rect 410524 449964 410576 450016
rect 3516 449896 3568 449948
rect 413284 449896 413336 449948
rect 169024 449828 169076 449880
rect 340052 449828 340104 449880
rect 171048 449760 171100 449812
rect 318800 449760 318852 449812
rect 182088 449692 182140 449744
rect 300124 449692 300176 449744
rect 247040 449420 247092 449472
rect 338304 449420 338356 449472
rect 175188 449352 175240 449404
rect 338856 449352 338908 449404
rect 396724 449352 396776 449404
rect 464528 449352 464580 449404
rect 280160 449284 280212 449336
rect 490932 449284 490984 449336
rect 166724 449216 166776 449268
rect 424324 449216 424376 449268
rect 478420 449216 478472 449268
rect 537484 449216 537536 449268
rect 169116 449148 169168 449200
rect 174176 449148 174228 449200
rect 175188 449148 175240 449200
rect 243176 449148 243228 449200
rect 509792 449148 509844 449200
rect 197912 448468 197964 448520
rect 549720 448468 549772 448520
rect 169392 448400 169444 448452
rect 340328 448400 340380 448452
rect 169300 448332 169352 448384
rect 169668 448332 169720 448384
rect 339040 448332 339092 448384
rect 199384 448264 199436 448316
rect 214380 448264 214432 448316
rect 199752 448196 199804 448248
rect 215576 448196 215628 448248
rect 198556 448128 198608 448180
rect 216864 448128 216916 448180
rect 264612 448128 264664 448180
rect 337476 448128 337528 448180
rect 196716 448060 196768 448112
rect 219348 448060 219400 448112
rect 322480 448060 322532 448112
rect 399668 448060 399720 448112
rect 195704 447992 195756 448044
rect 218152 447992 218204 448044
rect 319996 447992 320048 448044
rect 399576 447992 399628 448044
rect 195796 447924 195848 447976
rect 220636 447924 220688 447976
rect 252100 447924 252152 447976
rect 337568 447924 337620 447976
rect 351184 447924 351236 447976
rect 459560 447924 459612 447976
rect 501236 447924 501288 447976
rect 548800 447924 548852 447976
rect 196992 447856 197044 447908
rect 221924 447856 221976 447908
rect 296076 447856 296128 447908
rect 405188 447856 405240 447908
rect 448520 447856 448572 447908
rect 522396 447856 522448 447908
rect 195612 447788 195664 447840
rect 223120 447788 223172 447840
rect 255688 447788 255740 447840
rect 503536 447788 503588 447840
rect 198648 447720 198700 447772
rect 213092 447720 213144 447772
rect 192760 447652 192812 447704
rect 204260 447652 204312 447704
rect 194508 447584 194560 447636
rect 205548 447584 205600 447636
rect 204536 447108 204588 447160
rect 449440 447108 449492 447160
rect 244556 446564 244608 446616
rect 338396 446564 338448 446616
rect 397460 446564 397512 446616
rect 466460 446564 466512 446616
rect 293040 446496 293092 446548
rect 436744 446496 436796 446548
rect 491024 446496 491076 446548
rect 543740 446496 543792 446548
rect 273168 446428 273220 446480
rect 494704 446428 494756 446480
rect 184204 446360 184256 446412
rect 452016 446360 452068 446412
rect 453672 446360 453724 446412
rect 524880 446360 524932 446412
rect 199844 445680 199896 445732
rect 226892 445680 226944 445732
rect 268384 445680 268436 445732
rect 341340 445680 341392 445732
rect 197176 445612 197228 445664
rect 225696 445612 225748 445664
rect 262128 445612 262180 445664
rect 339684 445612 339736 445664
rect 195888 445544 195940 445596
rect 228180 445544 228232 445596
rect 260840 445544 260892 445596
rect 339776 445544 339828 445596
rect 198464 445476 198516 445528
rect 230664 445476 230716 445528
rect 259644 445476 259696 445528
rect 339592 445476 339644 445528
rect 199568 445408 199620 445460
rect 231952 445408 232004 445460
rect 258356 445408 258408 445460
rect 341156 445408 341208 445460
rect 196624 445340 196676 445392
rect 229468 445340 229520 445392
rect 253296 445340 253348 445392
rect 337016 445340 337068 445392
rect 199660 445272 199712 445324
rect 234436 445272 234488 445324
rect 254584 445272 254636 445324
rect 338488 445272 338540 445324
rect 199476 445204 199528 445256
rect 233240 445204 233292 445256
rect 257068 445204 257120 445256
rect 341064 445204 341116 445256
rect 192852 445136 192904 445188
rect 235724 445136 235776 445188
rect 255872 445136 255924 445188
rect 341248 445136 341300 445188
rect 194232 445068 194284 445120
rect 237012 445068 237064 445120
rect 243268 445068 243320 445120
rect 338212 445068 338264 445120
rect 344284 445068 344336 445120
rect 460756 445068 460808 445120
rect 463608 445068 463660 445120
rect 529940 445068 529992 445120
rect 191656 445000 191708 445052
rect 238208 445000 238260 445052
rect 265624 445000 265676 445052
rect 498476 445000 498528 445052
rect 197084 444932 197136 444984
rect 224408 444932 224460 444984
rect 269672 444932 269724 444984
rect 342536 444932 342588 444984
rect 193036 444864 193088 444916
rect 211804 444864 211856 444916
rect 327540 444864 327592 444916
rect 399484 444864 399536 444916
rect 194416 444796 194468 444848
rect 210608 444796 210660 444848
rect 270960 444796 271012 444848
rect 340972 444796 341024 444848
rect 348424 443776 348476 443828
rect 456984 443776 457036 443828
rect 263508 443708 263560 443760
rect 499764 443708 499816 443760
rect 507124 443708 507176 443760
rect 551284 443708 551336 443760
rect 178776 443640 178828 443692
rect 439412 443640 439464 443692
rect 456708 443640 456760 443692
rect 526168 443640 526220 443692
rect 277216 442892 277268 442944
rect 337108 442892 337160 442944
rect 275928 442824 275980 442876
rect 339500 442824 339552 442876
rect 274732 442756 274784 442808
rect 338580 442756 338632 442808
rect 273444 442688 273496 442740
rect 339868 442688 339920 442740
rect 272156 442620 272208 442672
rect 340880 442620 340932 442672
rect 263416 442552 263468 442604
rect 336832 442552 336884 442604
rect 267188 442484 267240 442536
rect 342444 442484 342496 442536
rect 265900 442416 265952 442468
rect 342352 442416 342404 442468
rect 400956 442416 401008 442468
rect 434352 442416 434404 442468
rect 191748 442348 191800 442400
rect 239496 442348 239548 442400
rect 278688 442348 278740 442400
rect 492220 442348 492272 442400
rect 177304 442280 177356 442332
rect 450728 442280 450780 442332
rect 487068 442280 487120 442332
rect 541256 442280 541308 442332
rect 234528 442212 234580 442264
rect 514852 442212 514904 442264
rect 278504 442144 278556 442196
rect 337200 442144 337252 442196
rect 279700 442076 279752 442128
rect 337292 442076 337344 442128
rect 167920 441532 167972 441584
rect 443000 441532 443052 441584
rect 358084 441056 358136 441108
rect 454500 441056 454552 441108
rect 285588 440988 285640 441040
rect 471244 440988 471296 441040
rect 260748 440920 260800 440972
rect 501052 440920 501104 440972
rect 186964 440852 187016 440904
rect 448244 440852 448296 440904
rect 471888 440852 471940 440904
rect 533712 440852 533764 440904
rect 167828 440172 167880 440224
rect 437664 440172 437716 440224
rect 169760 440104 169812 440156
rect 438952 440104 439004 440156
rect 333796 439764 333848 439816
rect 409420 439764 409472 439816
rect 356704 439696 356756 439748
rect 458180 439696 458232 439748
rect 187792 439628 187844 439680
rect 444472 439628 444524 439680
rect 476764 439628 476816 439680
rect 535000 439628 535052 439680
rect 306288 439560 306340 439612
rect 478420 439560 478472 439612
rect 188344 439492 188396 439544
rect 444472 439492 444524 439544
rect 447048 439492 447100 439544
rect 521108 439492 521160 439544
rect 168012 438880 168064 438932
rect 169760 438880 169812 438932
rect 173256 438812 173308 438864
rect 187792 438812 187844 438864
rect 393964 438336 394016 438388
rect 462044 438336 462096 438388
rect 288348 438268 288400 438320
rect 485044 438268 485096 438320
rect 275836 438200 275888 438252
rect 493508 438200 493560 438252
rect 497464 438200 497516 438252
rect 545028 438200 545080 438252
rect 186964 438132 187016 438184
rect 432052 438132 432104 438184
rect 459468 438132 459520 438184
rect 527456 438132 527508 438184
rect 314936 436840 314988 436892
rect 409236 436840 409288 436892
rect 485136 436840 485188 436892
rect 538772 436840 538824 436892
rect 284208 436772 284260 436824
rect 489736 436772 489788 436824
rect 248236 436704 248288 436756
rect 507308 436704 507360 436756
rect 473360 435480 473412 435532
rect 548524 435480 548576 435532
rect 309048 435412 309100 435464
rect 477132 435412 477184 435464
rect 251088 435344 251140 435396
rect 506020 435344 506072 435396
rect 191564 434052 191616 434104
rect 426808 434052 426860 434104
rect 451188 434052 451240 434104
rect 523684 434052 523736 434104
rect 253848 433984 253900 434036
rect 504824 433984 504876 434036
rect 511908 433984 511960 434036
rect 553860 433984 553912 434036
rect 326252 432692 326304 432744
rect 398104 432692 398156 432744
rect 292304 432624 292356 432676
rect 409328 432624 409380 432676
rect 467104 432624 467156 432676
rect 531228 432624 531280 432676
rect 245568 432556 245620 432608
rect 508596 432556 508648 432608
rect 331312 431536 331364 431588
rect 340144 431536 340196 431588
rect 241980 431468 242032 431520
rect 336740 431468 336792 431520
rect 353944 431468 353996 431520
rect 455788 431468 455840 431520
rect 462228 431468 462280 431520
rect 528652 431468 528704 431520
rect 259368 431400 259420 431452
rect 502248 431400 502300 431452
rect 198556 431332 198608 431384
rect 465080 431332 465132 431384
rect 199200 431264 199252 431316
rect 468024 431264 468076 431316
rect 198372 431196 198424 431248
rect 467932 431196 467984 431248
rect 567936 430584 567988 430636
rect 579896 430584 579948 430636
rect 323768 430244 323820 430296
rect 391204 430244 391256 430296
rect 405004 430244 405056 430296
rect 463332 430244 463384 430296
rect 291108 430176 291160 430228
rect 447784 430176 447836 430228
rect 198740 430108 198792 430160
rect 459744 430108 459796 430160
rect 198924 430040 198976 430092
rect 461032 430040 461084 430092
rect 199016 429972 199068 430024
rect 462412 429972 462464 430024
rect 198648 429904 198700 429956
rect 462320 429904 462372 429956
rect 199108 429836 199160 429888
rect 466552 429836 466604 429888
rect 175372 429088 175424 429140
rect 451372 429088 451424 429140
rect 178040 429020 178092 429072
rect 452752 429020 452804 429072
rect 170312 428952 170364 429004
rect 171508 428952 171560 429004
rect 428464 428952 428516 429004
rect 303528 428680 303580 428732
rect 479616 428680 479668 428732
rect 198832 428612 198884 428664
rect 458272 428612 458324 428664
rect 198464 428544 198516 428596
rect 463792 428544 463844 428596
rect 177856 428476 177908 428528
rect 455512 428476 455564 428528
rect 178776 428408 178828 428460
rect 456892 428408 456944 428460
rect 474004 428408 474056 428460
rect 532424 428408 532476 428460
rect 173624 427796 173676 427848
rect 175372 427796 175424 427848
rect 177304 427796 177356 427848
rect 178040 427796 178092 427848
rect 173716 427728 173768 427780
rect 445852 427728 445904 427780
rect 180340 427660 180392 427712
rect 180800 427660 180852 427712
rect 447232 427660 447284 427712
rect 172152 427592 172204 427644
rect 198832 427592 198884 427644
rect 304908 427116 304960 427168
rect 409144 427116 409196 427168
rect 441528 427116 441580 427168
rect 518624 427116 518676 427168
rect 191748 427048 191800 427100
rect 448612 427048 448664 427100
rect 488448 427048 488500 427100
rect 542544 427048 542596 427100
rect 184204 426436 184256 426488
rect 392860 426436 392912 426488
rect 172336 426368 172388 426420
rect 172888 426368 172940 426420
rect 445760 426368 445812 426420
rect 173164 426300 173216 426352
rect 190460 426300 190512 426352
rect 191748 426300 191800 426352
rect 328736 425892 328788 425944
rect 396816 425892 396868 425944
rect 321192 425824 321244 425876
rect 400864 425824 400916 425876
rect 318708 425756 318760 425808
rect 406384 425756 406436 425808
rect 504364 425756 504416 425808
rect 550088 425756 550140 425808
rect 313648 425688 313700 425740
rect 405096 425688 405148 425740
rect 480904 425688 480956 425740
rect 536196 425688 536248 425740
rect 332508 425008 332560 425060
rect 342720 425008 342772 425060
rect 288532 424940 288584 424992
rect 341708 424940 341760 424992
rect 287244 424872 287296 424924
rect 342904 424872 342956 424924
rect 286048 424804 286100 424856
rect 342812 424804 342864 424856
rect 300768 424736 300820 424788
rect 480628 424736 480680 424788
rect 299388 424668 299440 424720
rect 481916 424668 481968 424720
rect 296628 424600 296680 424652
rect 483204 424600 483256 424652
rect 241428 424532 241480 424584
rect 510804 424532 510856 424584
rect 238668 424464 238720 424516
rect 512184 424464 512236 424516
rect 235908 424396 235960 424448
rect 513380 424396 513432 424448
rect 231768 424328 231820 424380
rect 516140 424328 516192 424380
rect 170128 423580 170180 423632
rect 440240 423580 440292 423632
rect 171416 423512 171468 423564
rect 437572 423512 437624 423564
rect 245752 423036 245804 423088
rect 338120 423036 338172 423088
rect 487804 423036 487856 423088
rect 539692 423036 539744 423088
rect 271788 422968 271840 423020
rect 495716 422968 495768 423020
rect 199384 422900 199436 422952
rect 213368 422900 213420 422952
rect 269028 422900 269080 422952
rect 497004 422900 497056 422952
rect 168104 422288 168156 422340
rect 171416 422288 171468 422340
rect 410524 422152 410576 422204
rect 425244 422152 425296 422204
rect 407856 422084 407908 422136
rect 435364 422084 435416 422136
rect 408132 422016 408184 422068
rect 436652 422016 436704 422068
rect 407948 421948 408000 422000
rect 440332 421948 440384 422000
rect 530584 421948 530636 422000
rect 545948 421948 546000 422000
rect 408040 421880 408092 421932
rect 441712 421880 441764 421932
rect 471244 421880 471296 421932
rect 488172 421880 488224 421932
rect 514668 421880 514720 421932
rect 554780 421880 554832 421932
rect 284760 421812 284812 421864
rect 342260 421812 342312 421864
rect 407764 421812 407816 421864
rect 446588 421812 446640 421864
rect 447784 421812 447836 421864
rect 485780 421812 485832 421864
rect 509148 421812 509200 421864
rect 552204 421812 552256 421864
rect 341524 421744 341576 421796
rect 427820 421744 427872 421796
rect 436744 421744 436796 421796
rect 484400 421744 484452 421796
rect 499488 421744 499540 421796
rect 547236 421744 547288 421796
rect 196624 421676 196676 421728
rect 397644 421676 397696 421728
rect 409788 421676 409840 421728
rect 470692 421676 470744 421728
rect 474648 421676 474700 421728
rect 546684 421676 546736 421728
rect 193864 421608 193916 421660
rect 400220 421608 400272 421660
rect 408316 421608 408368 421660
rect 471980 421608 472032 421660
rect 475844 421608 475896 421660
rect 547880 421608 547932 421660
rect 199568 421540 199620 421592
rect 407580 421540 407632 421592
rect 408408 421540 408460 421592
rect 465540 421540 465592 421592
rect 469588 421540 469640 421592
rect 546776 421540 546828 421592
rect 195244 421472 195296 421524
rect 403900 421472 403952 421524
rect 196992 421404 197044 421456
rect 408868 421404 408920 421456
rect 197084 421336 197136 421388
rect 415400 421336 415452 421388
rect 197176 421268 197228 421320
rect 416780 421268 416832 421320
rect 173164 421200 173216 421252
rect 393780 421200 393832 421252
rect 173256 421132 173308 421184
rect 398932 421132 398984 421184
rect 172152 421064 172204 421116
rect 406476 421064 406528 421116
rect 172244 420996 172296 421048
rect 412824 420996 412876 421048
rect 413284 420996 413336 421048
rect 420276 420996 420328 421048
rect 173532 420928 173584 420980
rect 414020 420928 414072 420980
rect 485044 420928 485096 420980
rect 487160 420928 487212 420980
rect 199476 420180 199528 420232
rect 213184 420180 213236 420232
rect 181444 419704 181496 419756
rect 402980 419704 403032 419756
rect 195520 419636 195572 419688
rect 418988 419636 419040 419688
rect 184388 419568 184440 419620
rect 410156 419568 410208 419620
rect 187516 419500 187568 419552
rect 417700 419500 417752 419552
rect 179052 419432 179104 419484
rect 197360 419432 197412 419484
rect 189816 416712 189868 416764
rect 197360 416712 197412 416764
rect 177580 415352 177632 415404
rect 197360 415352 197412 415404
rect 560208 415352 560260 415404
rect 580264 415352 580316 415404
rect 182916 413924 182968 413976
rect 197360 413924 197412 413976
rect 184480 412564 184532 412616
rect 197360 412564 197412 412616
rect 3424 411204 3476 411256
rect 28448 411204 28500 411256
rect 188528 411204 188580 411256
rect 197360 411204 197412 411256
rect 170956 409776 171008 409828
rect 197360 409776 197412 409828
rect 191288 409708 191340 409760
rect 197452 409708 197504 409760
rect 170220 408416 170272 408468
rect 171324 408416 171376 408468
rect 194048 408416 194100 408468
rect 197360 408416 197412 408468
rect 560116 408416 560168 408468
rect 577504 408416 577556 408468
rect 195428 407056 195480 407108
rect 197728 407056 197780 407108
rect 181628 405628 181680 405680
rect 197360 405628 197412 405680
rect 574836 404336 574888 404388
rect 580172 404336 580224 404388
rect 192484 404268 192536 404320
rect 197360 404268 197412 404320
rect 185676 401548 185728 401600
rect 197360 401548 197412 401600
rect 170864 400120 170916 400172
rect 197360 400120 197412 400172
rect 560024 400120 560076 400172
rect 570604 400120 570656 400172
rect 3240 398760 3292 398812
rect 28356 398760 28408 398812
rect 170772 398760 170824 398812
rect 197360 398760 197412 398812
rect 174636 398692 174688 398744
rect 197452 398692 197504 398744
rect 168840 398284 168892 398336
rect 169944 398284 169996 398336
rect 174728 397400 174780 397452
rect 197360 397400 197412 397452
rect 176200 395972 176252 396024
rect 197360 395972 197412 396024
rect 187148 394612 187200 394664
rect 197360 394612 197412 394664
rect 169484 393252 169536 393304
rect 174176 393252 174228 393304
rect 177488 393252 177540 393304
rect 197360 393252 197412 393304
rect 169116 391960 169168 392012
rect 169484 391960 169536 392012
rect 184296 391892 184348 391944
rect 197360 391892 197412 391944
rect 560208 391892 560260 391944
rect 578884 391892 578936 391944
rect 188436 390464 188488 390516
rect 197360 390464 197412 390516
rect 191196 389104 191248 389156
rect 197360 389104 197412 389156
rect 180064 387744 180116 387796
rect 197360 387744 197412 387796
rect 195336 386316 195388 386368
rect 197728 386316 197780 386368
rect 193956 386248 194008 386300
rect 197360 386248 197412 386300
rect 167736 384956 167788 385008
rect 197360 384956 197412 385008
rect 178960 383596 179012 383648
rect 197360 383596 197412 383648
rect 559196 383392 559248 383444
rect 560944 383392 560996 383444
rect 167644 382168 167696 382220
rect 197360 382168 197412 382220
rect 181536 380808 181588 380860
rect 197360 380808 197412 380860
rect 167552 379448 167604 379500
rect 197360 379448 197412 379500
rect 570604 378156 570656 378208
rect 580172 378156 580224 378208
rect 188712 378088 188764 378140
rect 197360 378088 197412 378140
rect 175004 376660 175056 376712
rect 197360 376660 197412 376712
rect 187424 375300 187476 375352
rect 197360 375300 197412 375352
rect 560208 375300 560260 375352
rect 567844 375300 567896 375352
rect 184756 373940 184808 373992
rect 197360 373940 197412 373992
rect 177764 372512 177816 372564
rect 197360 372512 197412 372564
rect 193772 372444 193824 372496
rect 197452 372444 197504 372496
rect 195152 371152 195204 371204
rect 197360 371152 197412 371204
rect 190000 369792 190052 369844
rect 197360 369792 197412 369844
rect 185860 368432 185912 368484
rect 197360 368432 197412 368484
rect 559196 367412 559248 367464
rect 565084 367412 565136 367464
rect 183100 367004 183152 367056
rect 197360 367004 197412 367056
rect 3424 365644 3476 365696
rect 197176 365644 197228 365696
rect 174912 365576 174964 365628
rect 197360 365576 197412 365628
rect 3424 365100 3476 365152
rect 197820 365100 197872 365152
rect 3608 365032 3660 365084
rect 199568 365032 199620 365084
rect 3516 364964 3568 365016
rect 200120 364964 200172 365016
rect 559564 364352 559616 364404
rect 579620 364352 579672 364404
rect 139216 364284 139268 364336
rect 168104 364284 168156 364336
rect 176384 364284 176436 364336
rect 197360 364284 197412 364336
rect 167184 364148 167236 364200
rect 178776 364148 178828 364200
rect 136548 364080 136600 364132
rect 168196 364080 168248 364132
rect 130936 363944 130988 363996
rect 172336 363944 172388 363996
rect 125508 363876 125560 363928
rect 173624 363876 173676 363928
rect 29644 363808 29696 363860
rect 42800 363808 42852 363860
rect 129648 363808 129700 363860
rect 180340 363808 180392 363860
rect 122748 363740 122800 363792
rect 177304 363740 177356 363792
rect 28632 363672 28684 363724
rect 42892 363672 42944 363724
rect 29736 363604 29788 363656
rect 46940 363604 46992 363656
rect 128268 363604 128320 363656
rect 190460 363604 190512 363656
rect 167736 363536 167788 363588
rect 170956 363536 171008 363588
rect 177856 363536 177908 363588
rect 148968 363468 149020 363520
rect 170312 363468 170364 363520
rect 136548 363332 136600 363384
rect 146944 363332 146996 363384
rect 137928 363264 137980 363316
rect 167828 363264 167880 363316
rect 29460 362924 29512 362976
rect 29644 362924 29696 362976
rect 151176 362924 151228 362976
rect 167092 362924 167144 362976
rect 169852 362924 169904 362976
rect 184940 362924 184992 362976
rect 187792 362924 187844 362976
rect 180156 362856 180208 362908
rect 197360 362856 197412 362908
rect 138296 362380 138348 362432
rect 180340 362380 180392 362432
rect 124128 362312 124180 362364
rect 170772 362312 170824 362364
rect 146944 362244 146996 362296
rect 168012 362244 168064 362296
rect 184296 362244 184348 362296
rect 108856 362176 108908 362228
rect 177304 362176 177356 362228
rect 167920 361496 167972 361548
rect 169760 361496 169812 361548
rect 179144 361496 179196 361548
rect 197360 361496 197412 361548
rect 181812 361428 181864 361480
rect 197452 361428 197504 361480
rect 150440 361088 150492 361140
rect 167184 361088 167236 361140
rect 171048 361088 171100 361140
rect 133144 361020 133196 361072
rect 167920 361020 167972 361072
rect 127624 360952 127676 361004
rect 170956 360952 171008 361004
rect 143356 360884 143408 360936
rect 167000 360884 167052 360936
rect 186964 360884 187016 360936
rect 193220 360884 193272 360936
rect 73160 360816 73212 360868
rect 176384 360816 176436 360868
rect 140320 360136 140372 360188
rect 193680 360136 193732 360188
rect 194600 360136 194652 360188
rect 560208 360136 560260 360188
rect 574744 360136 574796 360188
rect 125968 360068 126020 360120
rect 173808 360068 173860 360120
rect 176752 360068 176804 360120
rect 177672 360068 177724 360120
rect 197360 360068 197412 360120
rect 135904 359524 135956 359576
rect 174728 359524 174780 359576
rect 103152 359456 103204 359508
rect 167644 359456 167696 359508
rect 3332 358708 3384 358760
rect 195520 358708 195572 358760
rect 114376 358640 114428 358692
rect 172612 358640 172664 358692
rect 173808 358640 173860 358692
rect 188620 358640 188672 358692
rect 197360 358640 197412 358692
rect 132040 358096 132092 358148
rect 184940 358096 184992 358148
rect 63408 358028 63460 358080
rect 166264 358028 166316 358080
rect 173808 358028 173860 358080
rect 187884 358028 187936 358080
rect 184664 357348 184716 357400
rect 197360 357348 197412 357400
rect 132960 356872 133012 356924
rect 181812 356872 181864 356924
rect 136456 356804 136508 356856
rect 191840 356804 191892 356856
rect 119988 356736 120040 356788
rect 189172 356736 189224 356788
rect 95608 356668 95660 356720
rect 167828 356668 167880 356720
rect 109592 355988 109644 356040
rect 169852 355988 169904 356040
rect 170220 355988 170272 356040
rect 187240 355988 187292 356040
rect 197360 355988 197412 356040
rect 169852 355512 169904 355564
rect 174636 355512 174688 355564
rect 128268 355444 128320 355496
rect 178776 355444 178828 355496
rect 128176 355376 128228 355428
rect 187148 355376 187200 355428
rect 85672 355308 85724 355360
rect 185676 355308 185728 355360
rect 115756 354628 115808 354680
rect 171232 354628 171284 354680
rect 172428 354628 172480 354680
rect 191472 354356 191524 354408
rect 197360 354356 197412 354408
rect 172428 354152 172480 354204
rect 191196 354152 191248 354204
rect 129556 354084 129608 354136
rect 180064 354084 180116 354136
rect 125416 354016 125468 354068
rect 195428 354016 195480 354068
rect 88248 353948 88300 354000
rect 173716 353948 173768 354000
rect 180248 353200 180300 353252
rect 197360 353200 197412 353252
rect 111616 352588 111668 352640
rect 167736 352588 167788 352640
rect 75828 352520 75880 352572
rect 174912 352520 174964 352572
rect 176292 351840 176344 351892
rect 197360 351840 197412 351892
rect 559656 351840 559708 351892
rect 566464 351840 566516 351892
rect 130936 351364 130988 351416
rect 170864 351364 170916 351416
rect 124036 351296 124088 351348
rect 172336 351296 172388 351348
rect 118516 351228 118568 351280
rect 195336 351228 195388 351280
rect 198832 351228 198884 351280
rect 99288 351160 99340 351212
rect 181904 351160 181956 351212
rect 112996 350480 113048 350532
rect 173992 350480 174044 350532
rect 175188 350480 175240 350532
rect 185768 350480 185820 350532
rect 197360 350480 197412 350532
rect 175188 350004 175240 350056
rect 183560 350004 183612 350056
rect 137928 349936 137980 349988
rect 190460 349936 190512 349988
rect 115848 349868 115900 349920
rect 176292 349868 176344 349920
rect 93768 349800 93820 349852
rect 182916 349800 182968 349852
rect 174820 349052 174872 349104
rect 197360 349052 197412 349104
rect 192668 348984 192720 349036
rect 197452 348984 197504 349036
rect 148968 348508 149020 348560
rect 178960 348508 179012 348560
rect 113088 348440 113140 348492
rect 179052 348440 179104 348492
rect 78588 348372 78640 348424
rect 188344 348372 188396 348424
rect 108948 347692 109000 347744
rect 169852 347692 169904 347744
rect 168288 347624 168340 347676
rect 197360 347624 197412 347676
rect 169852 347216 169904 347268
rect 185032 347216 185084 347268
rect 129648 347148 129700 347200
rect 182180 347148 182232 347200
rect 118608 347080 118660 347132
rect 174820 347080 174872 347132
rect 100668 347012 100720 347064
rect 180248 347012 180300 347064
rect 3332 346332 3384 346384
rect 187516 346332 187568 346384
rect 117228 346264 117280 346316
rect 172520 346264 172572 346316
rect 173808 346264 173860 346316
rect 183008 346264 183060 346316
rect 197360 346264 197412 346316
rect 139216 345720 139268 345772
rect 189080 345720 189132 345772
rect 84108 345652 84160 345704
rect 172428 345652 172480 345704
rect 173808 345652 173860 345704
rect 198740 345652 198792 345704
rect 143448 344972 143500 345024
rect 179236 344972 179288 345024
rect 189908 344972 189960 345024
rect 197360 344972 197412 345024
rect 121276 344428 121328 344480
rect 173624 344428 173676 344480
rect 125508 344360 125560 344412
rect 186320 344360 186372 344412
rect 106188 344292 106240 344344
rect 167920 344292 167972 344344
rect 179236 344292 179288 344344
rect 186964 344292 187016 344344
rect 191380 343544 191432 343596
rect 197360 343544 197412 343596
rect 560208 343544 560260 343596
rect 570696 343544 570748 343596
rect 131028 342932 131080 342984
rect 177488 342932 177540 342984
rect 91008 342864 91060 342916
rect 184480 342864 184532 342916
rect 142068 342184 142120 342236
rect 187332 342184 187384 342236
rect 192576 342184 192628 342236
rect 197360 342184 197412 342236
rect 122748 341504 122800 341556
rect 176200 341504 176252 341556
rect 29828 340892 29880 340944
rect 46940 340892 46992 340944
rect 187332 340892 187384 340944
rect 187792 340892 187844 340944
rect 114468 340824 114520 340876
rect 171140 340824 171192 340876
rect 171692 340824 171744 340876
rect 181720 340824 181772 340876
rect 197360 340824 197412 340876
rect 171692 340416 171744 340468
rect 181628 340416 181680 340468
rect 135168 340348 135220 340400
rect 181536 340348 181588 340400
rect 68928 340280 68980 340332
rect 176844 340280 176896 340332
rect 29552 340212 29604 340264
rect 46204 340212 46256 340264
rect 66168 340212 66220 340264
rect 194876 340212 194928 340264
rect 3976 340144 4028 340196
rect 197084 340144 197136 340196
rect 28540 339532 28592 339584
rect 35164 339532 35216 339584
rect 60648 339396 60700 339448
rect 197360 339396 197412 339448
rect 121184 339328 121236 339380
rect 184572 339328 184624 339380
rect 184848 339328 184900 339380
rect 71688 338988 71740 339040
rect 168012 338988 168064 339040
rect 81348 338920 81400 338972
rect 187240 338920 187292 338972
rect 4068 338852 4120 338904
rect 172244 338852 172296 338904
rect 3884 338784 3936 338836
rect 173532 338784 173584 338836
rect 184848 338784 184900 338836
rect 196808 338784 196860 338836
rect 3792 338716 3844 338768
rect 196992 338716 197044 338768
rect 166264 338036 166316 338088
rect 197360 338036 197412 338088
rect 176844 336676 176896 336728
rect 197360 336676 197412 336728
rect 194876 336608 194928 336660
rect 197452 336608 197504 336660
rect 168012 335248 168064 335300
rect 197360 335248 197412 335300
rect 560208 335248 560260 335300
rect 578976 335248 579028 335300
rect 176384 333888 176436 333940
rect 197360 333888 197412 333940
rect 174912 332528 174964 332580
rect 197360 332528 197412 332580
rect 188344 331168 188396 331220
rect 197360 331168 197412 331220
rect 187240 329740 187292 329792
rect 197360 329740 197412 329792
rect 172428 328380 172480 328432
rect 197360 328380 197412 328432
rect 559932 328380 559984 328432
rect 565176 328380 565228 328432
rect 185676 327020 185728 327072
rect 197360 327020 197412 327072
rect 173716 325592 173768 325644
rect 197360 325592 197412 325644
rect 565084 324300 565136 324352
rect 580080 324300 580132 324352
rect 182916 324232 182968 324284
rect 197452 324232 197504 324284
rect 184480 324164 184532 324216
rect 197360 324164 197412 324216
rect 167828 322872 167880 322924
rect 197360 322872 197412 322924
rect 181904 321512 181956 321564
rect 197360 321512 197412 321564
rect 180248 320084 180300 320136
rect 197360 320084 197412 320136
rect 559380 320084 559432 320136
rect 566556 320084 566608 320136
rect 167644 318724 167696 318776
rect 197360 318724 197412 318776
rect 167920 317364 167972 317416
rect 197360 317364 197412 317416
rect 177304 315936 177356 315988
rect 197360 315936 197412 315988
rect 167736 314576 167788 314628
rect 197360 314576 197412 314628
rect 176292 313216 176344 313268
rect 197452 313216 197504 313268
rect 179052 313148 179104 313200
rect 197360 313148 197412 313200
rect 577504 311856 577556 311908
rect 580448 311856 580500 311908
rect 174820 311788 174872 311840
rect 197360 311788 197412 311840
rect 560208 311788 560260 311840
rect 577596 311788 577648 311840
rect 173624 310428 173676 310480
rect 197360 310428 197412 310480
rect 172336 309068 172388 309120
rect 197360 309068 197412 309120
rect 195428 307708 195480 307760
rect 197728 307708 197780 307760
rect 187148 306280 187200 306332
rect 197360 306280 197412 306332
rect 177488 304920 177540 304972
rect 197360 304920 197412 304972
rect 181812 303560 181864 303612
rect 197360 303560 197412 303612
rect 559288 303424 559340 303476
rect 561036 303424 561088 303476
rect 174728 302132 174780 302184
rect 197360 302132 197412 302184
rect 180340 300772 180392 300824
rect 197360 300772 197412 300824
rect 173532 299480 173584 299532
rect 197360 299480 197412 299532
rect 174728 298120 174780 298172
rect 197360 298120 197412 298172
rect 560944 298120 560996 298172
rect 580172 298120 580224 298172
rect 167644 296692 167696 296744
rect 197360 296692 197412 296744
rect 559012 296624 559064 296676
rect 580356 296624 580408 296676
rect 177304 295332 177356 295384
rect 197360 295332 197412 295384
rect 172244 293972 172296 294024
rect 197360 293972 197412 294024
rect 173624 292544 173676 292596
rect 197360 292544 197412 292596
rect 167736 291184 167788 291236
rect 197360 291184 197412 291236
rect 180248 289824 180300 289876
rect 197360 289824 197412 289876
rect 174820 288396 174872 288448
rect 197360 288396 197412 288448
rect 560208 288328 560260 288380
rect 567936 288328 567988 288380
rect 176292 287104 176344 287156
rect 197452 287104 197504 287156
rect 167920 287036 167972 287088
rect 197360 287036 197412 287088
rect 172336 285676 172388 285728
rect 197360 285676 197412 285728
rect 168012 284316 168064 284368
rect 197360 284316 197412 284368
rect 168104 282888 168156 282940
rect 197360 282888 197412 282940
rect 181720 281528 181772 281580
rect 197360 281528 197412 281580
rect 167828 280168 167880 280220
rect 197360 280168 197412 280220
rect 559932 280100 559984 280152
rect 574836 280100 574888 280152
rect 168196 278740 168248 278792
rect 197360 278740 197412 278792
rect 177488 277380 177540 277432
rect 197360 277380 197412 277432
rect 174912 276088 174964 276140
rect 197360 276088 197412 276140
rect 173716 276020 173768 276072
rect 197452 276020 197504 276072
rect 172428 274660 172480 274712
rect 197360 274660 197412 274712
rect 180340 273232 180392 273284
rect 197360 273232 197412 273284
rect 171048 271872 171100 271924
rect 197360 271872 197412 271924
rect 566464 271872 566516 271924
rect 579804 271872 579856 271924
rect 187148 270512 187200 270564
rect 197360 270512 197412 270564
rect 183008 267724 183060 267776
rect 197360 267724 197412 267776
rect 181812 266364 181864 266416
rect 197360 266364 197412 266416
rect 179052 264936 179104 264988
rect 197360 264936 197412 264988
rect 169208 264188 169260 264240
rect 182916 264188 182968 264240
rect 176384 263644 176436 263696
rect 197452 263644 197504 263696
rect 171692 263576 171744 263628
rect 197360 263576 197412 263628
rect 560208 263508 560260 263560
rect 570604 263508 570656 263560
rect 168288 262216 168340 262268
rect 197360 262216 197412 262268
rect 168564 261468 168616 261520
rect 195428 261468 195480 261520
rect 187240 260856 187292 260908
rect 197360 260856 197412 260908
rect 169852 258068 169904 258120
rect 197360 258068 197412 258120
rect 567844 258068 567896 258120
rect 580172 258068 580224 258120
rect 560024 256640 560076 256692
rect 578884 256640 578936 256692
rect 166724 254532 166776 254584
rect 197820 254532 197872 254584
rect 27528 253852 27580 253904
rect 197912 253852 197964 253904
rect 128084 253784 128136 253836
rect 179052 253784 179104 253836
rect 115664 253716 115716 253768
rect 171048 253716 171100 253768
rect 125508 253648 125560 253700
rect 181812 253648 181864 253700
rect 123024 253580 123076 253632
rect 183008 253580 183060 253632
rect 118332 253512 118384 253564
rect 187148 253512 187200 253564
rect 98276 253444 98328 253496
rect 167828 253444 167880 253496
rect 75552 253376 75604 253428
rect 167736 253376 167788 253428
rect 70676 253308 70728 253360
rect 172244 253308 172296 253360
rect 65708 253240 65760 253292
rect 167644 253240 167696 253292
rect 28356 253172 28408 253224
rect 29460 253172 29512 253224
rect 43352 253172 43404 253224
rect 60648 253172 60700 253224
rect 173532 253172 173584 253224
rect 130568 253104 130620 253156
rect 176384 253104 176436 253156
rect 132960 253036 133012 253088
rect 171692 253036 171744 253088
rect 27068 252492 27120 252544
rect 27252 252492 27304 252544
rect 28448 252492 28500 252544
rect 34520 252492 34572 252544
rect 198004 252492 198056 252544
rect 167000 252424 167052 252476
rect 197452 252424 197504 252476
rect 68192 252356 68244 252408
rect 177304 252356 177356 252408
rect 189264 252356 189316 252408
rect 190368 252356 190420 252408
rect 197360 252356 197412 252408
rect 78128 252288 78180 252340
rect 180248 252288 180300 252340
rect 73160 252220 73212 252272
rect 173624 252220 173676 252272
rect 83556 252152 83608 252204
rect 176292 252152 176344 252204
rect 95608 252084 95660 252136
rect 181720 252084 181772 252136
rect 85672 252016 85724 252068
rect 167920 252016 167972 252068
rect 90824 251948 90876 252000
rect 168012 251948 168064 252000
rect 93216 251880 93268 251932
rect 168104 251880 168156 251932
rect 100576 251812 100628 251864
rect 168196 251812 168248 251864
rect 175004 251812 175056 251864
rect 189264 251812 189316 251864
rect 120908 251744 120960 251796
rect 166724 251744 166776 251796
rect 167000 251744 167052 251796
rect 167828 251744 167880 251796
rect 135996 251676 136048 251728
rect 168288 251676 168340 251728
rect 151084 251608 151136 251660
rect 167000 251608 167052 251660
rect 63408 251540 63460 251592
rect 174728 251540 174780 251592
rect 81256 251132 81308 251184
rect 174820 251132 174872 251184
rect 88248 251064 88300 251116
rect 172336 251064 172388 251116
rect 103152 250996 103204 251048
rect 177488 250996 177540 251048
rect 106096 250928 106148 250980
rect 173716 250928 173768 250980
rect 113088 250860 113140 250912
rect 180340 250860 180392 250912
rect 108488 250792 108540 250844
rect 174912 250792 174964 250844
rect 110512 250724 110564 250776
rect 172428 250724 172480 250776
rect 138296 250656 138348 250708
rect 187240 250656 187292 250708
rect 129556 249704 129608 249756
rect 193588 249704 193640 249756
rect 114376 249636 114428 249688
rect 174544 249636 174596 249688
rect 175188 249636 175240 249688
rect 143356 249568 143408 249620
rect 176844 249568 176896 249620
rect 193588 249160 193640 249212
rect 194692 249160 194744 249212
rect 176844 249092 176896 249144
rect 177396 249092 177448 249144
rect 186412 249092 186464 249144
rect 175188 249024 175240 249076
rect 192024 249024 192076 249076
rect 114468 248344 114520 248396
rect 176108 248344 176160 248396
rect 560208 248344 560260 248396
rect 577504 248344 577556 248396
rect 132040 248276 132092 248328
rect 191104 248276 191156 248328
rect 126888 248208 126940 248260
rect 176660 248208 176712 248260
rect 176660 247120 176712 247172
rect 177396 247120 177448 247172
rect 176108 247052 176160 247104
rect 177304 247052 177356 247104
rect 191104 247052 191156 247104
rect 193404 247052 193456 247104
rect 28816 246984 28868 247036
rect 197360 246984 197412 247036
rect 124128 246916 124180 246968
rect 179420 246916 179472 246968
rect 140688 246304 140740 246356
rect 167644 246304 167696 246356
rect 179420 245624 179472 245676
rect 180248 245624 180300 245676
rect 28172 245556 28224 245608
rect 197360 245556 197412 245608
rect 122748 245488 122800 245540
rect 169852 245488 169904 245540
rect 169852 244876 169904 244928
rect 170680 244876 170732 244928
rect 180800 244876 180852 244928
rect 28540 244196 28592 244248
rect 197360 244196 197412 244248
rect 112996 244128 113048 244180
rect 172060 244128 172112 244180
rect 179144 244128 179196 244180
rect 143448 244060 143500 244112
rect 176016 244060 176068 244112
rect 176016 243516 176068 243568
rect 183652 243516 183704 243568
rect 28724 242836 28776 242888
rect 197360 242836 197412 242888
rect 119988 242768 120040 242820
rect 189724 242768 189776 242820
rect 190000 242768 190052 242820
rect 190000 242156 190052 242208
rect 196900 242156 196952 242208
rect 3240 241408 3292 241460
rect 184388 241408 184440 241460
rect 121276 241340 121328 241392
rect 173440 241340 173492 241392
rect 173808 241340 173860 241392
rect 173808 240728 173860 240780
rect 191104 240728 191156 240780
rect 115848 240048 115900 240100
rect 175280 240048 175332 240100
rect 129648 239980 129700 240032
rect 173900 239980 173952 240032
rect 560208 239572 560260 239624
rect 565084 239572 565136 239624
rect 182916 239368 182968 239420
rect 195980 239368 196032 239420
rect 173900 239232 173952 239284
rect 174728 239232 174780 239284
rect 195980 238892 196032 238944
rect 197360 238892 197412 238944
rect 107568 238688 107620 238740
rect 168196 238688 168248 238740
rect 128268 238620 128320 238672
rect 187700 238620 187752 238672
rect 47584 238008 47636 238060
rect 175004 238008 175056 238060
rect 178684 238008 178736 238060
rect 197360 238008 197412 238060
rect 168196 237396 168248 237448
rect 185584 237396 185636 237448
rect 117228 237328 117280 237380
rect 174084 237328 174136 237380
rect 142068 237260 142120 237312
rect 175924 237260 175976 237312
rect 175924 236716 175976 236768
rect 189264 236716 189316 236768
rect 28448 236648 28500 236700
rect 197452 236648 197504 236700
rect 174084 235968 174136 236020
rect 174544 235968 174596 236020
rect 118608 235900 118660 235952
rect 185952 235900 186004 235952
rect 195428 235900 195480 235952
rect 197728 235900 197780 235952
rect 139216 235832 139268 235884
rect 171968 235832 172020 235884
rect 172428 235832 172480 235884
rect 185952 235356 186004 235408
rect 195428 235356 195480 235408
rect 172428 235288 172480 235340
rect 188436 235288 188488 235340
rect 28908 235220 28960 235272
rect 197544 235220 197596 235272
rect 108948 234540 109000 234592
rect 169852 234540 169904 234592
rect 121184 234472 121236 234524
rect 172704 234472 172756 234524
rect 173348 234472 173400 234524
rect 131028 234404 131080 234456
rect 182088 234404 182140 234456
rect 183744 234404 183796 234456
rect 169852 233860 169904 233912
rect 170588 233860 170640 233912
rect 182824 233860 182876 233912
rect 179052 233248 179104 233300
rect 197360 233248 197412 233300
rect 110328 233180 110380 233232
rect 171784 233180 171836 233232
rect 172428 233180 172480 233232
rect 178040 233180 178092 233232
rect 178868 233180 178920 233232
rect 125508 233112 125560 233164
rect 172428 232568 172480 232620
rect 181720 232568 181772 232620
rect 178960 232500 179012 232552
rect 197360 232500 197412 232552
rect 565084 231820 565136 231872
rect 579804 231820 579856 231872
rect 111708 231752 111760 231804
rect 173072 231752 173124 231804
rect 180340 231752 180392 231804
rect 183008 231752 183060 231804
rect 183192 231752 183244 231804
rect 197360 231752 197412 231804
rect 559196 231684 559248 231736
rect 560944 231684 560996 231736
rect 148324 231072 148376 231124
rect 171140 231072 171192 231124
rect 183008 231072 183060 231124
rect 29828 230392 29880 230444
rect 47584 230392 47636 230444
rect 180156 229712 180208 229764
rect 197544 229712 197596 229764
rect 28724 229576 28776 229628
rect 29828 229576 29880 229628
rect 28540 229100 28592 229152
rect 29644 229032 29696 229084
rect 46756 229032 46808 229084
rect 50344 229032 50396 229084
rect 135168 229032 135220 229084
rect 168564 229032 168616 229084
rect 185032 229032 185084 229084
rect 198372 229032 198424 229084
rect 136456 228964 136508 229016
rect 170496 228964 170548 229016
rect 191196 228964 191248 229016
rect 198924 228964 198976 229016
rect 170496 228556 170548 228608
rect 177580 228556 177632 228608
rect 176108 228488 176160 228540
rect 185032 228488 185084 228540
rect 174636 228420 174688 228472
rect 191932 228420 191984 228472
rect 199108 228420 199160 228472
rect 3700 228352 3752 228404
rect 195244 228352 195296 228404
rect 29828 227740 29880 227792
rect 34520 227740 34572 227792
rect 35164 227740 35216 227792
rect 168564 227740 168616 227792
rect 187148 227740 187200 227792
rect 133788 227672 133840 227724
rect 187056 227672 187108 227724
rect 192484 227672 192536 227724
rect 198556 227672 198608 227724
rect 137928 227604 137980 227656
rect 171876 227604 171928 227656
rect 172428 227604 172480 227656
rect 136364 227536 136416 227588
rect 170220 227536 170272 227588
rect 170220 227128 170272 227180
rect 180892 227128 180944 227180
rect 172428 227060 172480 227112
rect 193956 227060 194008 227112
rect 3884 226992 3936 227044
rect 172152 226992 172204 227044
rect 187056 226312 187108 226364
rect 189356 226312 189408 226364
rect 183560 226244 183612 226296
rect 198464 226244 198516 226296
rect 171784 225564 171836 225616
rect 183560 225564 183612 225616
rect 181628 224204 181680 224256
rect 185032 224204 185084 224256
rect 197360 224204 197412 224256
rect 187884 223524 187936 223576
rect 199016 223524 199068 223576
rect 199568 223524 199620 223576
rect 560208 223524 560260 223576
rect 567844 223524 567896 223576
rect 171876 222844 171928 222896
rect 187884 222844 187936 222896
rect 193496 220804 193548 220856
rect 198924 220804 198976 220856
rect 184388 220056 184440 220108
rect 197360 220056 197412 220108
rect 195336 218764 195388 218816
rect 197912 218764 197964 218816
rect 174820 218696 174872 218748
rect 193496 218696 193548 218748
rect 559564 218016 559616 218068
rect 579896 218016 579948 218068
rect 189172 217948 189224 218000
rect 197360 217948 197412 218000
rect 171048 217268 171100 217320
rect 189172 217268 189224 217320
rect 170956 215908 171008 215960
rect 197360 215908 197412 215960
rect 198004 215908 198056 215960
rect 559196 215772 559248 215824
rect 566464 215772 566516 215824
rect 196808 215364 196860 215416
rect 197728 215364 197780 215416
rect 198096 215364 198148 215416
rect 176200 213936 176252 213988
rect 179420 213936 179472 213988
rect 197360 213936 197412 213988
rect 170772 213188 170824 213240
rect 178132 213188 178184 213240
rect 178132 212508 178184 212560
rect 197360 212508 197412 212560
rect 186320 212440 186372 212492
rect 197636 212440 197688 212492
rect 167920 211760 167972 211812
rect 186320 211760 186372 211812
rect 197636 211556 197688 211608
rect 197912 211556 197964 211608
rect 176660 211080 176712 211132
rect 197360 211080 197412 211132
rect 170772 210400 170824 210452
rect 176660 210400 176712 210452
rect 197360 210196 197412 210248
rect 197728 210196 197780 210248
rect 197728 210060 197780 210112
rect 198004 210060 198056 210112
rect 182916 209176 182968 209228
rect 197360 209176 197412 209228
rect 197728 209176 197780 209228
rect 197912 209176 197964 209228
rect 178776 209040 178828 209092
rect 180984 209040 181036 209092
rect 176200 208292 176252 208344
rect 182180 208292 182232 208344
rect 197360 208292 197412 208344
rect 560208 208292 560260 208344
rect 580264 208292 580316 208344
rect 180064 206320 180116 206372
rect 196072 206320 196124 206372
rect 197360 206320 197412 206372
rect 170956 206252 171008 206304
rect 180984 206252 181036 206304
rect 197728 206252 197780 206304
rect 170864 204892 170916 204944
rect 186320 204892 186372 204944
rect 186320 204280 186372 204332
rect 186504 204280 186556 204332
rect 197360 204280 197412 204332
rect 168104 204212 168156 204264
rect 169760 204212 169812 204264
rect 197728 204212 197780 204264
rect 184940 204144 184992 204196
rect 185400 204144 185452 204196
rect 197360 204144 197412 204196
rect 168012 203532 168064 203584
rect 185400 203532 185452 203584
rect 181536 202784 181588 202836
rect 187884 202784 187936 202836
rect 191288 202784 191340 202836
rect 197912 202784 197964 202836
rect 187884 201492 187936 201544
rect 197360 201492 197412 201544
rect 168196 200744 168248 200796
rect 191840 200744 191892 200796
rect 197360 200744 197412 200796
rect 184296 199384 184348 199436
rect 193312 199384 193364 199436
rect 197360 199384 197412 199436
rect 168288 197956 168340 198008
rect 190460 197956 190512 198008
rect 197360 197956 197412 198008
rect 189080 197276 189132 197328
rect 197360 197276 197412 197328
rect 173440 196596 173492 196648
rect 189080 196596 189132 196648
rect 194600 195916 194652 195968
rect 197360 195916 197412 195968
rect 181628 195236 181680 195288
rect 194600 195236 194652 195288
rect 187792 194488 187844 194540
rect 197360 194488 197412 194540
rect 174912 193808 174964 193860
rect 187792 193808 187844 193860
rect 177764 192448 177816 192500
rect 193220 192448 193272 192500
rect 197728 192448 197780 192500
rect 186964 191836 187016 191888
rect 190460 191836 190512 191888
rect 197360 191836 197412 191888
rect 560944 191836 560996 191888
rect 580172 191836 580224 191888
rect 560208 191700 560260 191752
rect 565084 191700 565136 191752
rect 185584 191088 185636 191140
rect 197360 191088 197412 191140
rect 182824 189728 182876 189780
rect 197360 189728 197412 189780
rect 181720 188300 181772 188352
rect 197360 188300 197412 188352
rect 181536 187688 181588 187740
rect 181720 187688 181772 187740
rect 180064 186940 180116 186992
rect 180340 186940 180392 186992
rect 197360 186940 197412 186992
rect 178684 185580 178736 185632
rect 179144 185580 179196 185632
rect 197360 185580 197412 185632
rect 560024 184832 560076 184884
rect 580264 184832 580316 184884
rect 177304 184152 177356 184204
rect 197360 184152 197412 184204
rect 170496 182792 170548 182844
rect 192024 182792 192076 182844
rect 197360 182792 197412 182844
rect 175280 182112 175332 182164
rect 175740 182112 175792 182164
rect 197360 182112 197412 182164
rect 170404 181432 170456 181484
rect 175740 181432 175792 181484
rect 174544 180072 174596 180124
rect 197360 180072 197412 180124
rect 195244 179460 195296 179512
rect 197360 179460 197412 179512
rect 168932 178644 168984 178696
rect 181720 178644 181772 178696
rect 196808 178236 196860 178288
rect 197912 178236 197964 178288
rect 169300 177352 169352 177404
rect 180340 177352 180392 177404
rect 173348 177284 173400 177336
rect 197360 177284 197412 177336
rect 560208 176604 560260 176656
rect 580172 176604 580224 176656
rect 168932 175992 168984 176044
rect 178224 175992 178276 176044
rect 169208 175924 169260 175976
rect 197636 175924 197688 175976
rect 191104 175652 191156 175704
rect 197360 175652 197412 175704
rect 182088 175176 182140 175228
rect 197360 175176 197412 175228
rect 168840 174564 168892 174616
rect 175004 174564 175056 174616
rect 170680 174496 170732 174548
rect 180800 174496 180852 174548
rect 182088 174496 182140 174548
rect 180248 173204 180300 173256
rect 197360 173204 197412 173256
rect 168748 173136 168800 173188
rect 194600 173136 194652 173188
rect 174636 172456 174688 172508
rect 178040 172456 178092 172508
rect 197360 172456 197412 172508
rect 168932 171776 168984 171828
rect 177856 171776 177908 171828
rect 169116 170484 169168 170536
rect 178960 170484 179012 170536
rect 177396 170416 177448 170468
rect 197360 170416 197412 170468
rect 169024 170348 169076 170400
rect 197544 170348 197596 170400
rect 187700 169668 187752 169720
rect 197360 169668 197412 169720
rect 178776 168988 178828 169040
rect 187700 168988 187752 169040
rect 194692 168308 194744 168360
rect 197544 168308 197596 168360
rect 559012 168240 559064 168292
rect 560944 168240 560996 168292
rect 184296 167696 184348 167748
rect 194692 167696 194744 167748
rect 174728 167628 174780 167680
rect 197360 167628 197412 167680
rect 184848 166948 184900 167000
rect 197360 166948 197412 167000
rect 177488 166268 177540 166320
rect 183744 166268 183796 166320
rect 184848 166268 184900 166320
rect 559564 165588 559616 165640
rect 580172 165588 580224 165640
rect 178868 164908 178920 164960
rect 193404 164908 193456 164960
rect 197360 164908 197412 164960
rect 169116 164840 169168 164892
rect 195980 164840 196032 164892
rect 188344 164160 188396 164212
rect 189356 164160 189408 164212
rect 197360 164160 197412 164212
rect 187148 162120 187200 162172
rect 197360 162120 197412 162172
rect 180800 161372 180852 161424
rect 197360 161372 197412 161424
rect 170588 160692 170640 160744
rect 180800 160692 180852 160744
rect 177580 159332 177632 159384
rect 197360 159332 197412 159384
rect 193956 158312 194008 158364
rect 197360 158312 197412 158364
rect 188436 156612 188488 156664
rect 197360 156612 197412 156664
rect 189080 155864 189132 155916
rect 189264 155864 189316 155916
rect 197544 155864 197596 155916
rect 167736 155252 167788 155304
rect 189080 155252 189132 155304
rect 167644 155184 167696 155236
rect 197360 155184 197412 155236
rect 184848 154504 184900 154556
rect 197360 154504 197412 154556
rect 175924 153824 175976 153876
rect 183652 153824 183704 153876
rect 184848 153824 184900 153876
rect 186320 153144 186372 153196
rect 197360 153144 197412 153196
rect 176016 152464 176068 152516
rect 186320 152464 186372 152516
rect 168748 151036 168800 151088
rect 179052 151036 179104 151088
rect 168564 150356 168616 150408
rect 197360 150424 197412 150476
rect 181720 149064 181772 149116
rect 187700 149064 187752 149116
rect 197360 149064 197412 149116
rect 180340 148996 180392 149048
rect 181904 148996 181956 149048
rect 180800 147636 180852 147688
rect 181904 147636 181956 147688
rect 197544 147636 197596 147688
rect 177672 147568 177724 147620
rect 178224 147568 178276 147620
rect 197360 147568 197412 147620
rect 175004 146208 175056 146260
rect 178040 146208 178092 146260
rect 178040 144916 178092 144968
rect 197360 144916 197412 144968
rect 560024 144848 560076 144900
rect 580264 144848 580316 144900
rect 191196 144712 191248 144764
rect 194600 144712 194652 144764
rect 197360 144712 197412 144764
rect 177856 144168 177908 144220
rect 194600 144168 194652 144220
rect 194600 143556 194652 143608
rect 197360 143556 197412 143608
rect 178960 142808 179012 142860
rect 186320 142808 186372 142860
rect 186320 142128 186372 142180
rect 197360 142128 197412 142180
rect 166172 141448 166224 141500
rect 197820 141448 197872 141500
rect 166264 141380 166316 141432
rect 197452 141380 197504 141432
rect 133144 141312 133196 141364
rect 168104 141312 168156 141364
rect 140044 141244 140096 141296
rect 181628 141244 181680 141296
rect 128544 141176 128596 141228
rect 176200 141176 176252 141228
rect 142344 141108 142396 141160
rect 190460 141108 190512 141160
rect 134248 141040 134300 141092
rect 187884 141040 187936 141092
rect 123760 140972 123812 141024
rect 178132 140972 178184 141024
rect 136548 140904 136600 140956
rect 193312 140904 193364 140956
rect 112168 140836 112220 140888
rect 171784 140836 171836 140888
rect 108488 140768 108540 140820
rect 176108 140768 176160 140820
rect 137928 140700 137980 140752
rect 168288 140700 168340 140752
rect 135352 140632 135404 140684
rect 168196 140632 168248 140684
rect 141240 140564 141292 140616
rect 174912 140564 174964 140616
rect 139032 140496 139084 140548
rect 173440 140496 173492 140548
rect 143448 140428 143500 140480
rect 177764 140428 177816 140480
rect 132040 140360 132092 140412
rect 168012 140360 168064 140412
rect 125968 140292 126020 140344
rect 170772 140292 170824 140344
rect 118976 140224 119028 140276
rect 171048 140224 171100 140276
rect 116768 140156 116820 140208
rect 184388 140156 184440 140208
rect 29828 140088 29880 140140
rect 35900 140088 35952 140140
rect 113272 140088 113324 140140
rect 185032 140088 185084 140140
rect 109592 140020 109644 140072
rect 191932 140020 191984 140072
rect 167828 139952 167880 140004
rect 197360 139952 197412 140004
rect 167000 139884 167052 139936
rect 197268 139884 197320 139936
rect 149520 139408 149572 139460
rect 167000 139408 167052 139460
rect 120356 139340 120408 139392
rect 191288 139340 191340 139392
rect 559564 139340 559616 139392
rect 580172 139340 580224 139392
rect 129648 139272 129700 139324
rect 196072 139272 196124 139324
rect 121368 139204 121420 139256
rect 182916 139204 182968 139256
rect 115480 139136 115532 139188
rect 174820 139136 174872 139188
rect 107384 139068 107436 139120
rect 166264 139068 166316 139120
rect 114376 139000 114428 139052
rect 171876 139000 171928 139052
rect 110880 138932 110932 138984
rect 169024 138932 169076 138984
rect 122656 138864 122708 138916
rect 179420 138864 179472 138916
rect 28816 138796 28868 138848
rect 43444 138796 43496 138848
rect 130752 138796 130804 138848
rect 186504 138796 186556 138848
rect 117872 138728 117924 138780
rect 169208 138728 169260 138780
rect 28632 138660 28684 138712
rect 43076 138660 43128 138712
rect 127716 138660 127768 138712
rect 170956 138660 171008 138712
rect 125232 138592 125284 138644
rect 167920 138592 167972 138644
rect 28356 138524 28408 138576
rect 28816 138524 28868 138576
rect 148416 138524 148468 138576
rect 166172 138524 166224 138576
rect 151084 138456 151136 138508
rect 167092 138456 167144 138508
rect 167092 138252 167144 138304
rect 167828 138252 167880 138304
rect 60648 137980 60700 138032
rect 117228 137980 117280 138032
rect 3332 137912 3384 137964
rect 181444 137912 181496 137964
rect 63224 137844 63276 137896
rect 197360 137844 197412 137896
rect 117228 137776 117280 137828
rect 197452 137776 197504 137828
rect 164884 136824 164936 136876
rect 168564 136824 168616 136876
rect 65800 136552 65852 136604
rect 197360 136552 197412 136604
rect 136456 135872 136508 135924
rect 194048 135872 194100 135924
rect 559288 135328 559340 135380
rect 560944 135328 560996 135380
rect 68928 135192 68980 135244
rect 197360 135192 197412 135244
rect 124128 134512 124180 134564
rect 178960 134512 179012 134564
rect 71044 133832 71096 133884
rect 197360 133832 197412 133884
rect 118424 133152 118476 133204
rect 180248 133152 180300 133204
rect 74448 132404 74500 132456
rect 197360 132404 197412 132456
rect 75828 132336 75880 132388
rect 197452 132336 197504 132388
rect 78588 131044 78640 131096
rect 197360 131044 197412 131096
rect 121368 130364 121420 130416
rect 181444 130364 181496 130416
rect 81348 129684 81400 129736
rect 197360 129684 197412 129736
rect 125416 129004 125468 129056
rect 174820 129004 174872 129056
rect 84108 128256 84160 128308
rect 197360 128256 197412 128308
rect 128268 127576 128320 127628
rect 177764 127576 177816 127628
rect 86868 126896 86920 126948
rect 197360 126896 197412 126948
rect 560944 126896 560996 126948
rect 580172 126896 580224 126948
rect 133788 126284 133840 126336
rect 167828 126284 167880 126336
rect 115848 126216 115900 126268
rect 184388 126216 184440 126268
rect 88248 125536 88300 125588
rect 197360 125536 197412 125588
rect 131028 124856 131080 124908
rect 174912 124856 174964 124908
rect 91008 124108 91060 124160
rect 197360 124108 197412 124160
rect 139308 123496 139360 123548
rect 180340 123496 180392 123548
rect 113088 123428 113140 123480
rect 171784 123428 171836 123480
rect 93768 122748 93820 122800
rect 197360 122748 197412 122800
rect 96528 121388 96580 121440
rect 197360 121388 197412 121440
rect 99288 120028 99340 120080
rect 197360 120028 197412 120080
rect 100668 119960 100720 120012
rect 197452 119960 197504 120012
rect 558920 118668 558972 118720
rect 561036 118668 561088 118720
rect 103428 118600 103480 118652
rect 197360 118600 197412 118652
rect 35900 117240 35952 117292
rect 164884 117240 164936 117292
rect 168564 117240 168616 117292
rect 28724 117172 28776 117224
rect 46940 117172 46992 117224
rect 106188 117172 106240 117224
rect 197360 117172 197412 117224
rect 28540 117104 28592 117156
rect 45836 117104 45888 117156
rect 108948 115880 109000 115932
rect 197360 115880 197412 115932
rect 3792 115336 3844 115388
rect 173256 115336 173308 115388
rect 3884 115268 3936 115320
rect 193864 115268 193916 115320
rect 3608 115200 3660 115252
rect 196716 115200 196768 115252
rect 111708 114452 111760 114504
rect 197360 114452 197412 114504
rect 3700 113840 3752 113892
rect 173164 113840 173216 113892
rect 4068 113772 4120 113824
rect 196624 113772 196676 113824
rect 171784 113092 171836 113144
rect 197360 113092 197412 113144
rect 561036 113092 561088 113144
rect 579804 113092 579856 113144
rect 559196 111800 559248 111852
rect 560944 111800 560996 111852
rect 184388 111732 184440 111784
rect 197360 111732 197412 111784
rect 180248 110372 180300 110424
rect 197360 110372 197412 110424
rect 178960 108944 179012 108996
rect 197544 108944 197596 108996
rect 181444 108876 181496 108928
rect 197360 108876 197412 108928
rect 174820 107584 174872 107636
rect 197452 107584 197504 107636
rect 177764 106224 177816 106276
rect 197360 106224 197412 106276
rect 174912 104796 174964 104848
rect 197360 104796 197412 104848
rect 560208 103776 560260 103828
rect 566464 103776 566516 103828
rect 167828 103436 167880 103488
rect 197360 103436 197412 103488
rect 194048 102076 194100 102128
rect 197360 102076 197412 102128
rect 180340 100648 180392 100700
rect 197360 100648 197412 100700
rect 559564 100648 559616 100700
rect 580172 100648 580224 100700
rect 167828 97996 167880 98048
rect 197360 97996 197412 98048
rect 559748 95208 559800 95260
rect 565084 95208 565136 95260
rect 178960 93848 179012 93900
rect 197360 93848 197412 93900
rect 167920 92488 167972 92540
rect 197360 92488 197412 92540
rect 176108 91060 176160 91112
rect 197360 91060 197412 91112
rect 177764 89700 177816 89752
rect 197360 89700 197412 89752
rect 176200 88340 176252 88392
rect 197360 88340 197412 88392
rect 174820 86980 174872 87032
rect 197360 86980 197412 87032
rect 560208 86980 560260 87032
rect 574836 86980 574888 87032
rect 560944 86912 560996 86964
rect 580172 86912 580224 86964
rect 173164 85552 173216 85604
rect 197360 85552 197412 85604
rect 169024 84192 169076 84244
rect 197360 84192 197412 84244
rect 168012 82832 168064 82884
rect 197360 82832 197412 82884
rect 174912 81472 174964 81524
rect 197452 81472 197504 81524
rect 173256 81404 173308 81456
rect 197360 81404 197412 81456
rect 175004 80044 175056 80096
rect 197360 80044 197412 80096
rect 169116 78684 169168 78736
rect 197360 78684 197412 78736
rect 560024 78684 560076 78736
rect 577504 78684 577556 78736
rect 168196 77256 168248 77308
rect 197360 77256 197412 77308
rect 171784 75896 171836 75948
rect 197360 75896 197412 75948
rect 168104 74536 168156 74588
rect 197360 74536 197412 74588
rect 169208 73176 169260 73228
rect 197360 73176 197412 73228
rect 565084 73108 565136 73160
rect 580172 73108 580224 73160
rect 559196 71816 559248 71868
rect 560944 71816 560996 71868
rect 173440 71748 173492 71800
rect 197360 71748 197412 71800
rect 176292 70388 176344 70440
rect 197360 70388 197412 70440
rect 168840 69640 168892 69692
rect 187700 69640 187752 69692
rect 168840 66172 168892 66224
rect 180800 66172 180852 66224
rect 168840 64812 168892 64864
rect 177672 64812 177724 64864
rect 168932 64132 168984 64184
rect 191196 64132 191248 64184
rect 170956 63520 171008 63572
rect 197360 63520 197412 63572
rect 560208 63520 560260 63572
rect 570604 63520 570656 63572
rect 169392 63452 169444 63504
rect 178040 63452 178092 63504
rect 168840 61344 168892 61396
rect 194600 61344 194652 61396
rect 172060 60732 172112 60784
rect 197360 60732 197412 60784
rect 566464 60664 566516 60716
rect 580172 60664 580224 60716
rect 169300 59372 169352 59424
rect 197544 59372 197596 59424
rect 168840 59304 168892 59356
rect 186320 59304 186372 59356
rect 560944 58624 560996 58676
rect 580356 58624 580408 58676
rect 196624 57808 196676 57860
rect 201500 58012 201552 58064
rect 202052 58012 202104 58064
rect 181444 57740 181496 57792
rect 206744 57876 206796 57928
rect 211804 57740 211856 57792
rect 214656 57740 214708 57792
rect 224132 57740 224184 57792
rect 471244 57740 471296 57792
rect 477684 57740 477736 57792
rect 480904 57740 480956 57792
rect 487068 57740 487120 57792
rect 502432 57740 502484 57792
rect 508044 57740 508096 57792
rect 171968 57672 172020 57724
rect 203156 57672 203208 57724
rect 214564 57672 214616 57724
rect 175096 57604 175148 57656
rect 217600 57604 217652 57656
rect 171876 57536 171928 57588
rect 214748 57536 214800 57588
rect 407212 57672 407264 57724
rect 407764 57672 407816 57724
rect 419540 57672 419592 57724
rect 420092 57672 420144 57724
rect 420920 57672 420972 57724
rect 421564 57672 421616 57724
rect 423680 57672 423732 57724
rect 424508 57672 424560 57724
rect 425060 57672 425112 57724
rect 425980 57672 426032 57724
rect 438124 57672 438176 57724
rect 439228 57672 439280 57724
rect 467104 57672 467156 57724
rect 475476 57672 475528 57724
rect 478144 57672 478196 57724
rect 484860 57672 484912 57724
rect 487804 57672 487856 57724
rect 495716 57672 495768 57724
rect 503720 57672 503772 57724
rect 508780 57672 508832 57724
rect 522580 57672 522632 57724
rect 525892 57672 525944 57724
rect 541348 57672 541400 57724
rect 556344 57672 556396 57724
rect 227720 57604 227772 57656
rect 228180 57604 228232 57656
rect 229100 57604 229152 57656
rect 229652 57604 229704 57656
rect 233240 57604 233292 57656
rect 233884 57604 233936 57656
rect 237380 57604 237432 57656
rect 238300 57604 238352 57656
rect 242900 57604 242952 57656
rect 243452 57604 243504 57656
rect 244280 57604 244332 57656
rect 244924 57604 244976 57656
rect 247040 57604 247092 57656
rect 247684 57604 247736 57656
rect 250536 57604 250588 57656
rect 253112 57604 253164 57656
rect 254860 57604 254912 57656
rect 255320 57604 255372 57656
rect 259460 57604 259512 57656
rect 260012 57604 260064 57656
rect 260840 57604 260892 57656
rect 261484 57604 261536 57656
rect 276020 57604 276072 57656
rect 276756 57604 276808 57656
rect 278044 57604 278096 57656
rect 279240 57604 279292 57656
rect 289820 57604 289872 57656
rect 290556 57604 290608 57656
rect 296720 57604 296772 57656
rect 297732 57604 297784 57656
rect 302240 57604 302292 57656
rect 302700 57604 302752 57656
rect 303620 57604 303672 57656
rect 304172 57604 304224 57656
rect 307760 57604 307812 57656
rect 308588 57604 308640 57656
rect 318800 57604 318852 57656
rect 319444 57604 319496 57656
rect 320180 57604 320232 57656
rect 320916 57604 320968 57656
rect 324320 57604 324372 57656
rect 325148 57604 325200 57656
rect 325700 57604 325752 57656
rect 326620 57604 326672 57656
rect 329840 57604 329892 57656
rect 330300 57604 330352 57656
rect 331220 57604 331272 57656
rect 331772 57604 331824 57656
rect 333980 57604 334032 57656
rect 334716 57604 334768 57656
rect 345020 57604 345072 57656
rect 345572 57604 345624 57656
rect 346492 57604 346544 57656
rect 347044 57604 347096 57656
rect 349160 57604 349212 57656
rect 349804 57604 349856 57656
rect 350632 57604 350684 57656
rect 351276 57604 351328 57656
rect 362960 57604 363012 57656
rect 363604 57604 363656 57656
rect 367100 57604 367152 57656
rect 368020 57604 368072 57656
rect 374000 57604 374052 57656
rect 374460 57604 374512 57656
rect 378140 57604 378192 57656
rect 378876 57604 378928 57656
rect 389180 57604 389232 57656
rect 389732 57604 389784 57656
rect 391940 57604 391992 57656
rect 392676 57604 392728 57656
rect 393412 57604 393464 57656
rect 393964 57604 394016 57656
rect 394700 57604 394752 57656
rect 395436 57604 395488 57656
rect 396080 57604 396132 57656
rect 396908 57604 396960 57656
rect 400220 57604 400272 57656
rect 445760 57604 445812 57656
rect 446404 57604 446456 57656
rect 447968 57604 448020 57656
rect 452660 57604 452712 57656
rect 453396 57604 453448 57656
rect 458916 57604 458968 57656
rect 460296 57604 460348 57656
rect 462320 57604 462372 57656
rect 462780 57604 462832 57656
rect 463700 57604 463752 57656
rect 464252 57604 464304 57656
rect 464344 57604 464396 57656
rect 250260 57536 250312 57588
rect 254584 57536 254636 57588
rect 263232 57536 263284 57588
rect 393320 57536 393372 57588
rect 441436 57536 441488 57588
rect 441620 57536 441672 57588
rect 442540 57536 442592 57588
rect 458824 57536 458876 57588
rect 471888 57536 471940 57588
rect 474004 57604 474056 57656
rect 476212 57604 476264 57656
rect 479800 57604 479852 57656
rect 486424 57604 486476 57656
rect 489276 57604 489328 57656
rect 489368 57604 489420 57656
rect 494980 57604 495032 57656
rect 477500 57536 477552 57588
rect 492864 57536 492916 57588
rect 177672 57468 177724 57520
rect 222016 57468 222068 57520
rect 224224 57468 224276 57520
rect 241520 57468 241572 57520
rect 247684 57468 247736 57520
rect 273444 57468 273496 57520
rect 386420 57468 386472 57520
rect 437112 57468 437164 57520
rect 467196 57468 467248 57520
rect 484124 57468 484176 57520
rect 488540 57468 488592 57520
rect 499396 57604 499448 57656
rect 505284 57604 505336 57656
rect 509516 57604 509568 57656
rect 513380 57604 513432 57656
rect 514300 57604 514352 57656
rect 514760 57604 514812 57656
rect 515772 57604 515824 57656
rect 524420 57604 524472 57656
rect 525156 57604 525208 57656
rect 534080 57604 534132 57656
rect 534540 57604 534592 57656
rect 536288 57604 536340 57656
rect 537484 57604 537536 57656
rect 538220 57604 538272 57656
rect 538956 57604 539008 57656
rect 539600 57604 539652 57656
rect 540244 57604 540296 57656
rect 543740 57604 543792 57656
rect 544660 57604 544712 57656
rect 550640 57604 550692 57656
rect 551284 57604 551336 57656
rect 554780 57604 554832 57656
rect 555516 57604 555568 57656
rect 504456 57536 504508 57588
rect 509332 57536 509384 57588
rect 512368 57536 512420 57588
rect 529756 57536 529808 57588
rect 534724 57536 534776 57588
rect 552204 57536 552256 57588
rect 567844 57536 567896 57588
rect 497004 57468 497056 57520
rect 498292 57468 498344 57520
rect 505928 57468 505980 57520
rect 510804 57468 510856 57520
rect 513104 57468 513156 57520
rect 542820 57468 542872 57520
rect 558184 57468 558236 57520
rect 170772 57400 170824 57452
rect 245844 57400 245896 57452
rect 246304 57400 246356 57452
rect 251640 57400 251692 57452
rect 254676 57400 254728 57452
rect 284668 57400 284720 57452
rect 284944 57400 284996 57452
rect 295892 57400 295944 57452
rect 377404 57400 377456 57452
rect 430580 57400 430632 57452
rect 459560 57400 459612 57452
rect 482008 57400 482060 57452
rect 485044 57400 485096 57452
rect 489368 57400 489420 57452
rect 494060 57400 494112 57452
rect 502984 57400 503036 57452
rect 535552 57400 535604 57452
rect 547144 57400 547196 57452
rect 549352 57400 549404 57452
rect 566464 57400 566516 57452
rect 188528 57332 188580 57384
rect 269764 57332 269816 57384
rect 271144 57332 271196 57384
rect 287152 57332 287204 57384
rect 287704 57332 287756 57384
rect 289360 57332 289412 57384
rect 350540 57332 350592 57384
rect 415400 57332 415452 57384
rect 440884 57332 440936 57384
rect 175188 57264 175240 57316
rect 258908 57264 258960 57316
rect 267004 57264 267056 57316
rect 272708 57264 272760 57316
rect 273904 57264 273956 57316
rect 293684 57264 293736 57316
rect 343640 57264 343692 57316
rect 410984 57264 411036 57316
rect 436100 57264 436152 57316
rect 467472 57264 467524 57316
rect 468484 57332 468536 57384
rect 468944 57264 468996 57316
rect 470600 57264 470652 57316
rect 482284 57332 482336 57384
rect 493600 57332 493652 57384
rect 500224 57332 500276 57384
rect 502248 57332 502300 57384
rect 529020 57332 529072 57384
rect 530584 57332 530636 57384
rect 543556 57332 543608 57384
rect 560300 57332 560352 57384
rect 170864 57196 170916 57248
rect 254308 57196 254360 57248
rect 258816 57196 258868 57248
rect 291476 57196 291528 57248
rect 338764 57196 338816 57248
rect 406660 57196 406712 57248
rect 407120 57196 407172 57248
rect 450084 57196 450136 57248
rect 454684 57196 454736 57248
rect 456616 57196 456668 57248
rect 456800 57196 456852 57248
rect 480536 57196 480588 57248
rect 486332 57264 486384 57316
rect 490196 57264 490248 57316
rect 500776 57264 500828 57316
rect 545764 57264 545816 57316
rect 564440 57264 564492 57316
rect 484400 57196 484452 57248
rect 496820 57196 496872 57248
rect 498200 57196 498252 57248
rect 505192 57196 505244 57248
rect 556620 57196 556672 57248
rect 582380 57196 582432 57248
rect 488632 57128 488684 57180
rect 264244 57060 264296 57112
rect 266176 57060 266228 57112
rect 518900 57060 518952 57112
rect 520280 57060 520332 57112
rect 531964 57060 532016 57112
rect 538864 57060 538916 57112
rect 231124 56924 231176 56976
rect 232872 56924 232924 56976
rect 277400 56788 277452 56840
rect 278228 56788 278280 56840
rect 523316 56788 523368 56840
rect 527180 56788 527232 56840
rect 499764 56720 499816 56772
rect 506572 56720 506624 56772
rect 506480 56652 506532 56704
rect 510620 56652 510672 56704
rect 233884 56584 233936 56636
rect 239404 56584 239456 56636
rect 410524 56584 410576 56636
rect 413192 56584 413244 56636
rect 443000 56584 443052 56636
rect 444012 56584 444064 56636
rect 447784 56584 447836 56636
rect 452292 56584 452344 56636
rect 476764 56584 476816 56636
rect 482744 56584 482796 56636
rect 508504 56584 508556 56636
rect 510252 56584 510304 56636
rect 527272 56244 527324 56296
rect 528100 56244 528152 56296
rect 269764 55972 269816 56024
rect 362500 55972 362552 56024
rect 258724 55904 258776 55956
rect 355232 55904 355284 55956
rect 364340 55904 364392 55956
rect 423312 55904 423364 55956
rect 426440 55904 426492 55956
rect 461676 55904 461728 55956
rect 171232 55836 171284 55888
rect 305276 55836 305328 55888
rect 308404 55836 308456 55888
rect 382740 55836 382792 55888
rect 383660 55836 383712 55888
rect 435640 55836 435692 55888
rect 448704 55836 448756 55888
rect 474740 55836 474792 55888
rect 483020 55836 483072 55888
rect 496452 55836 496504 55888
rect 533436 55836 533488 55888
rect 543832 55836 543884 55888
rect 546408 55836 546460 55888
rect 564532 55836 564584 55888
rect 471980 55564 472032 55616
rect 472900 55564 472952 55616
rect 456892 55428 456944 55480
rect 457812 55428 457864 55480
rect 454040 55360 454092 55412
rect 454868 55360 454920 55412
rect 346400 54680 346452 54732
rect 411904 54680 411956 54732
rect 276664 54612 276716 54664
rect 359004 54612 359056 54664
rect 244924 54544 244976 54596
rect 349252 54544 349304 54596
rect 440240 54544 440292 54596
rect 469956 54544 470008 54596
rect 487252 54544 487304 54596
rect 498384 54544 498436 54596
rect 178040 54476 178092 54528
rect 309140 54476 309192 54528
rect 311164 54476 311216 54528
rect 389272 54476 389324 54528
rect 405740 54476 405792 54528
rect 448520 54476 448572 54528
rect 476212 54476 476264 54528
rect 491484 54476 491536 54528
rect 552480 54476 552532 54528
rect 574744 54476 574796 54528
rect 298744 53252 298796 53304
rect 381544 53252 381596 53304
rect 268384 53184 268436 53236
rect 361580 53184 361632 53236
rect 226432 53116 226484 53168
rect 338672 53116 338724 53168
rect 412640 53116 412692 53168
rect 452752 53116 452804 53168
rect 200304 53048 200356 53100
rect 322020 53048 322072 53100
rect 367192 53048 367244 53100
rect 425152 53048 425204 53100
rect 444380 53048 444432 53100
rect 472072 53048 472124 53100
rect 473360 53048 473412 53100
rect 489920 53048 489972 53100
rect 554872 53048 554924 53100
rect 578884 53048 578936 53100
rect 285036 51892 285088 51944
rect 372712 51892 372764 51944
rect 266360 51824 266412 51876
rect 363052 51824 363104 51876
rect 209780 51756 209832 51808
rect 328552 51756 328604 51808
rect 379612 51756 379664 51808
rect 432144 51756 432196 51808
rect 184940 51688 184992 51740
rect 313280 51688 313332 51740
rect 360200 51688 360252 51740
rect 421012 51688 421064 51740
rect 430672 51688 430724 51740
rect 463792 51688 463844 51740
rect 554780 51688 554832 51740
rect 580264 51688 580316 51740
rect 309140 50464 309192 50516
rect 389180 50464 389232 50516
rect 238024 50396 238076 50448
rect 345112 50396 345164 50448
rect 218704 50328 218756 50380
rect 331312 50328 331364 50380
rect 374092 50328 374144 50380
rect 429200 50328 429252 50380
rect 433432 50328 433484 50380
rect 465540 50328 465592 50380
rect 330484 49172 330536 49224
rect 394700 49172 394752 49224
rect 313280 49104 313332 49156
rect 392032 49104 392084 49156
rect 226984 49036 227036 49088
rect 333152 49036 333204 49088
rect 173532 48968 173584 49020
rect 226524 48968 226576 49020
rect 233332 48968 233384 49020
rect 342260 48968 342312 49020
rect 394700 48968 394752 49020
rect 441712 48968 441764 49020
rect 455420 48968 455472 49020
rect 478972 48968 479024 49020
rect 334624 47744 334676 47796
rect 399484 47744 399536 47796
rect 257344 47676 257396 47728
rect 351920 47676 351972 47728
rect 407396 47676 407448 47728
rect 448612 47676 448664 47728
rect 220820 47608 220872 47660
rect 335360 47608 335412 47660
rect 218244 47540 218296 47592
rect 334072 47540 334124 47592
rect 339684 47540 339736 47592
rect 407212 47540 407264 47592
rect 447876 47540 447928 47592
rect 471980 47540 472032 47592
rect 574836 46860 574888 46912
rect 580172 46860 580224 46912
rect 276756 46316 276808 46368
rect 366180 46316 366232 46368
rect 416964 46316 417016 46368
rect 455512 46316 455564 46368
rect 240784 46248 240836 46300
rect 339500 46248 339552 46300
rect 179420 46180 179472 46232
rect 309876 46180 309928 46232
rect 353392 46180 353444 46232
rect 416872 46180 416924 46232
rect 250444 45024 250496 45076
rect 340972 45024 341024 45076
rect 280160 44956 280212 45008
rect 371240 44956 371292 45008
rect 191840 44888 191892 44940
rect 317420 44888 317472 44940
rect 450544 44888 450596 44940
rect 473452 44888 473504 44940
rect 172520 44820 172572 44872
rect 305000 44820 305052 44872
rect 340972 44820 341024 44872
rect 408592 44820 408644 44872
rect 409880 44820 409932 44872
rect 451372 44820 451424 44872
rect 317420 43596 317472 43648
rect 394792 43596 394844 43648
rect 236644 43528 236696 43580
rect 343824 43528 343876 43580
rect 216772 43460 216824 43512
rect 332600 43460 332652 43512
rect 193220 43392 193272 43444
rect 318892 43392 318944 43444
rect 348424 43392 348476 43444
rect 401692 43392 401744 43444
rect 414112 43392 414164 43444
rect 452660 43392 452712 43444
rect 287152 42236 287204 42288
rect 375472 42236 375524 42288
rect 247776 42168 247828 42220
rect 347872 42168 347924 42220
rect 194600 42100 194652 42152
rect 318800 42100 318852 42152
rect 176660 42032 176712 42084
rect 307852 42032 307904 42084
rect 351920 42032 351972 42084
rect 415492 42032 415544 42084
rect 428004 42032 428056 42084
rect 462412 42032 462464 42084
rect 304264 40876 304316 40928
rect 378232 40876 378284 40928
rect 245752 40808 245804 40860
rect 350724 40808 350776 40860
rect 198740 40740 198792 40792
rect 321560 40740 321612 40792
rect 183560 40672 183612 40724
rect 311900 40672 311952 40724
rect 342260 40672 342312 40724
rect 409972 40672 410024 40724
rect 240876 39448 240928 39500
rect 346584 39448 346636 39500
rect 205732 39380 205784 39432
rect 325792 39380 325844 39432
rect 327724 39380 327776 39432
rect 393504 39380 393556 39432
rect 397644 39380 397696 39432
rect 443092 39380 443144 39432
rect 186320 39312 186372 39364
rect 314752 39312 314804 39364
rect 335360 39312 335412 39364
rect 405832 39312 405884 39364
rect 297364 38020 297416 38072
rect 380900 38020 380952 38072
rect 259644 37952 259696 38004
rect 358820 37952 358872 38004
rect 231216 37884 231268 37936
rect 339592 37884 339644 37936
rect 356704 37884 356756 37936
rect 408500 37884 408552 37936
rect 289912 36660 289964 36712
rect 376852 36660 376904 36712
rect 254768 36592 254820 36644
rect 352012 36592 352064 36644
rect 209964 36524 210016 36576
rect 328460 36524 328512 36576
rect 378232 36524 378284 36576
rect 431960 36524 432012 36576
rect 316684 35368 316736 35420
rect 383844 35368 383896 35420
rect 236736 35300 236788 35352
rect 336832 35300 336884 35352
rect 201684 35232 201736 35284
rect 323032 35232 323084 35284
rect 384304 35232 384356 35284
rect 434720 35232 434772 35284
rect 190460 35164 190512 35216
rect 316224 35164 316276 35216
rect 332600 35164 332652 35216
rect 403164 35164 403216 35216
rect 250628 33872 250680 33924
rect 347780 33872 347832 33924
rect 172152 33804 172204 33856
rect 212632 33804 212684 33856
rect 217324 33804 217376 33856
rect 331220 33804 331272 33856
rect 365812 33804 365864 33856
rect 423772 33804 423824 33856
rect 207204 33736 207256 33788
rect 325700 33736 325752 33788
rect 328460 33736 328512 33788
rect 401600 33736 401652 33788
rect 320364 32580 320416 32632
rect 396172 32580 396224 32632
rect 264336 32512 264388 32564
rect 356060 32512 356112 32564
rect 228364 32444 228416 32496
rect 338120 32444 338172 32496
rect 195980 32376 196032 32428
rect 320272 32376 320324 32428
rect 396172 32376 396224 32428
rect 441620 32376 441672 32428
rect 169392 31220 169444 31272
rect 276112 31220 276164 31272
rect 283012 31220 283064 31272
rect 372804 31220 372856 31272
rect 208584 31152 208636 31204
rect 327080 31152 327132 31204
rect 189080 31084 189132 31136
rect 316040 31084 316092 31136
rect 382372 31084 382424 31136
rect 433524 31084 433576 31136
rect 168380 31016 168432 31068
rect 303712 31016 303764 31068
rect 318064 31016 318116 31068
rect 386604 31016 386656 31068
rect 433984 31016 434036 31068
rect 465080 31016 465132 31068
rect 143172 29860 143224 29912
rect 198188 29860 198240 29912
rect 135812 29792 135864 29844
rect 198096 29792 198148 29844
rect 128360 29724 128412 29776
rect 198556 29724 198608 29776
rect 237564 29724 237616 29776
rect 345020 29724 345072 29776
rect 127624 29656 127676 29708
rect 198372 29656 198424 29708
rect 211252 29656 211304 29708
rect 329932 29656 329984 29708
rect 370504 29656 370556 29708
rect 425060 29656 425112 29708
rect 124036 29588 124088 29640
rect 198280 29588 198332 29640
rect 204904 29588 204956 29640
rect 324412 29588 324464 29640
rect 331220 29588 331272 29640
rect 402980 29588 403032 29640
rect 429200 29588 429252 29640
rect 462320 29588 462372 29640
rect 166172 29520 166224 29572
rect 198648 29520 198700 29572
rect 166264 29452 166316 29504
rect 198464 29452 198516 29504
rect 166356 29384 166408 29436
rect 198004 29384 198056 29436
rect 130568 29044 130620 29096
rect 170956 29044 171008 29096
rect 138940 28976 138992 29028
rect 188436 28976 188488 29028
rect 134248 28908 134300 28960
rect 186964 28908 187016 28960
rect 143264 28840 143316 28892
rect 197912 28840 197964 28892
rect 103152 28772 103204 28824
rect 168196 28772 168248 28824
rect 90732 28704 90784 28756
rect 168012 28704 168064 28756
rect 88064 28636 88116 28688
rect 169024 28636 169076 28688
rect 83096 28568 83148 28620
rect 174820 28568 174872 28620
rect 80704 28500 80756 28552
rect 176200 28500 176252 28552
rect 78128 28432 78180 28484
rect 177764 28432 177816 28484
rect 75552 28364 75604 28416
rect 176108 28364 176160 28416
rect 60648 28296 60700 28348
rect 167828 28296 167880 28348
rect 244464 28296 244516 28348
rect 349160 28296 349212 28348
rect 68192 28228 68244 28280
rect 178960 28228 179012 28280
rect 224316 28228 224368 28280
rect 335452 28228 335504 28280
rect 389180 28228 389232 28280
rect 437572 28228 437624 28280
rect 128544 28160 128596 28212
rect 174728 28160 174780 28212
rect 135904 28092 135956 28144
rect 172060 28092 172112 28144
rect 138296 28024 138348 28076
rect 169300 28024 169352 28076
rect 28632 27548 28684 27600
rect 42800 27548 42852 27600
rect 120632 27548 120684 27600
rect 127624 27548 127676 27600
rect 132776 27548 132828 27600
rect 143264 27548 143316 27600
rect 150624 27548 150676 27600
rect 167092 27548 167144 27600
rect 28816 27480 28868 27532
rect 43628 27480 43680 27532
rect 143448 27480 143500 27532
rect 176016 27480 176068 27532
rect 118424 27412 118476 27464
rect 115664 27344 115716 27396
rect 124036 27344 124088 27396
rect 132040 27412 132092 27464
rect 178868 27412 178920 27464
rect 176292 27344 176344 27396
rect 124128 27276 124180 27328
rect 180156 27276 180208 27328
rect 129648 27208 129700 27260
rect 184296 27208 184348 27260
rect 126336 27140 126388 27192
rect 177396 27140 177448 27192
rect 123760 27072 123812 27124
rect 166264 27072 166316 27124
rect 128176 27004 128228 27056
rect 166172 27004 166224 27056
rect 214748 27004 214800 27056
rect 329840 27004 329892 27056
rect 112168 26936 112220 26988
rect 149060 26936 149112 26988
rect 150072 26936 150124 26988
rect 167000 26936 167052 26988
rect 204444 26936 204496 26988
rect 324320 26936 324372 26988
rect 324964 26936 325016 26988
rect 390652 26936 390704 26988
rect 110328 26868 110380 26920
rect 143356 26868 143408 26920
rect 143448 26868 143500 26920
rect 175924 26868 175976 26920
rect 193312 26868 193364 26920
rect 317512 26868 317564 26920
rect 327080 26868 327132 26920
rect 400312 26868 400364 26920
rect 418344 26868 418396 26920
rect 454684 26868 454736 26920
rect 64880 26800 64932 26852
rect 135812 26800 135864 26852
rect 140136 26800 140188 26852
rect 167644 26800 167696 26852
rect 141240 26732 141292 26784
rect 167736 26732 167788 26784
rect 63224 26664 63276 26716
rect 166356 26664 166408 26716
rect 71596 26596 71648 26648
rect 143172 26596 143224 26648
rect 98276 26188 98328 26240
rect 175004 26188 175056 26240
rect 100208 26120 100260 26172
rect 169116 26120 169168 26172
rect 105544 26052 105596 26104
rect 171784 26052 171836 26104
rect 142160 25984 142212 26036
rect 271144 25984 271196 26036
rect 157340 25916 157392 25968
rect 295432 25916 295484 25968
rect 154580 25848 154632 25900
rect 294052 25848 294104 25900
rect 128360 25780 128412 25832
rect 278044 25780 278096 25832
rect 114560 25712 114612 25764
rect 270592 25712 270644 25764
rect 104900 25644 104952 25696
rect 263692 25644 263744 25696
rect 60740 25576 60792 25628
rect 236092 25576 236144 25628
rect 294604 25576 294656 25628
rect 364524 25576 364576 25628
rect 60832 25508 60884 25560
rect 237472 25508 237524 25560
rect 271236 25508 271288 25560
rect 362960 25508 363012 25560
rect 363052 25508 363104 25560
rect 422300 25508 422352 25560
rect 431960 25508 432012 25560
rect 463700 25508 463752 25560
rect 111524 25440 111576 25492
rect 169208 25440 169260 25492
rect 112904 25372 112956 25424
rect 173440 25372 173492 25424
rect 108028 25304 108080 25356
rect 168104 25304 168156 25356
rect 147680 24760 147732 24812
rect 171140 24760 171192 24812
rect 86592 24692 86644 24744
rect 173164 24692 173216 24744
rect 92756 24624 92808 24676
rect 174912 24624 174964 24676
rect 162860 24556 162912 24608
rect 299572 24556 299624 24608
rect 146300 24488 146352 24540
rect 290004 24488 290056 24540
rect 140780 24420 140832 24472
rect 285772 24420 285824 24472
rect 111800 24352 111852 24404
rect 267832 24352 267884 24404
rect 89720 24284 89772 24336
rect 254860 24284 254912 24336
rect 85580 24216 85632 24268
rect 251272 24216 251324 24268
rect 46940 24148 46992 24200
rect 229192 24148 229244 24200
rect 10324 24080 10376 24132
rect 204352 24080 204404 24132
rect 290464 24080 290516 24132
rect 360384 24080 360436 24132
rect 392032 24080 392084 24132
rect 440332 24080 440384 24132
rect 454224 24080 454276 24132
rect 477592 24080 477644 24132
rect 135352 24012 135404 24064
rect 177580 24012 177632 24064
rect 73988 23944 74040 23996
rect 167920 23944 167972 23996
rect 95240 23876 95292 23928
rect 173256 23876 173308 23928
rect 106280 23400 106332 23452
rect 185584 23400 185636 23452
rect 88340 23332 88392 23384
rect 170864 23332 170916 23384
rect 165620 23264 165672 23316
rect 301044 23264 301096 23316
rect 167000 23196 167052 23248
rect 302332 23196 302384 23248
rect 164240 23128 164292 23180
rect 300860 23128 300912 23180
rect 139400 23060 139452 23112
rect 285680 23060 285732 23112
rect 107660 22992 107712 23044
rect 264244 22992 264296 23044
rect 69020 22924 69072 22976
rect 242992 22924 243044 22976
rect 53840 22856 53892 22908
rect 233424 22856 233476 22908
rect 37280 22788 37332 22840
rect 222292 22788 222344 22840
rect 306564 22788 306616 22840
rect 387892 22788 387944 22840
rect 2780 22720 2832 22772
rect 201592 22720 201644 22772
rect 286324 22720 286376 22772
rect 368572 22720 368624 22772
rect 385132 22720 385184 22772
rect 436192 22720 436244 22772
rect 440332 22720 440384 22772
rect 469220 22720 469272 22772
rect 118240 22652 118292 22704
rect 195244 22652 195296 22704
rect 110972 22584 111024 22636
rect 180064 22584 180116 22636
rect 120816 22516 120868 22568
rect 173348 22516 173400 22568
rect 108764 22040 108816 22092
rect 182824 22040 182876 22092
rect 120080 21972 120132 22024
rect 191104 21972 191156 22024
rect 149060 21904 149112 21956
rect 258816 21904 258868 21956
rect 158720 21836 158772 21888
rect 296812 21836 296864 21888
rect 132500 21768 132552 21820
rect 280344 21768 280396 21820
rect 126980 21700 127032 21752
rect 277492 21700 277544 21752
rect 4160 21632 4212 21684
rect 171968 21632 172020 21684
rect 185032 21632 185084 21684
rect 313372 21632 313424 21684
rect 62120 21564 62172 21616
rect 237380 21564 237432 21616
rect 57980 21496 58032 21548
rect 234712 21496 234764 21548
rect 360844 21496 360896 21548
rect 419632 21496 419684 21548
rect 34520 21428 34572 21480
rect 220912 21428 220964 21480
rect 316040 21428 316092 21480
rect 393412 21428 393464 21480
rect 16580 21360 16632 21412
rect 209872 21360 209924 21412
rect 278044 21360 278096 21412
rect 368480 21360 368532 21412
rect 415400 21360 415452 21412
rect 454132 21360 454184 21412
rect 117136 21292 117188 21344
rect 174544 21292 174596 21344
rect 3424 20612 3476 20664
rect 184204 20612 184256 20664
rect 577504 20612 577556 20664
rect 579620 20612 579672 20664
rect 138020 20476 138072 20528
rect 254676 20476 254728 20528
rect 182180 20408 182232 20460
rect 310612 20408 310664 20460
rect 150440 20340 150492 20392
rect 291292 20340 291344 20392
rect 147680 20272 147732 20324
rect 289820 20272 289872 20324
rect 96620 20204 96672 20256
rect 259552 20204 259604 20256
rect 38660 20136 38712 20188
rect 214656 20136 214708 20188
rect 51080 20068 51132 20120
rect 230572 20068 230624 20120
rect 48320 20000 48372 20052
rect 229100 20000 229152 20052
rect 324320 20000 324372 20052
rect 397552 20000 397604 20052
rect 22100 19932 22152 19984
rect 214012 19932 214064 19984
rect 253940 19932 253992 19984
rect 354680 19932 354732 19984
rect 402980 19932 403032 19984
rect 447232 19932 447284 19984
rect 151820 19116 151872 19168
rect 273904 19116 273956 19168
rect 161480 19048 161532 19100
rect 299480 19048 299532 19100
rect 135260 18980 135312 19032
rect 282920 18980 282972 19032
rect 23480 18912 23532 18964
rect 171876 18912 171928 18964
rect 175280 18912 175332 18964
rect 306472 18912 306524 18964
rect 127072 18844 127124 18896
rect 277400 18844 277452 18896
rect 84200 18776 84252 18828
rect 246304 18776 246356 18828
rect 69112 18708 69164 18760
rect 241612 18708 241664 18760
rect 357624 18708 357676 18760
rect 418436 18708 418488 18760
rect 44180 18640 44232 18692
rect 227812 18640 227864 18692
rect 302332 18640 302384 18692
rect 385040 18640 385092 18692
rect 26240 18572 26292 18624
rect 215392 18572 215444 18624
rect 273352 18572 273404 18624
rect 367284 18572 367336 18624
rect 423772 18572 423824 18624
rect 458916 18572 458968 18624
rect 530032 18572 530084 18624
rect 539784 18572 539836 18624
rect 118700 17756 118752 17808
rect 247684 17756 247736 17808
rect 160192 17688 160244 17740
rect 296720 17688 296772 17740
rect 160100 17620 160152 17672
rect 298100 17620 298152 17672
rect 143540 17552 143592 17604
rect 287244 17552 287296 17604
rect 136640 17484 136692 17536
rect 284300 17484 284352 17536
rect 131120 17416 131172 17468
rect 280252 17416 280304 17468
rect 67640 17348 67692 17400
rect 224224 17348 224276 17400
rect 93860 17280 93912 17332
rect 256884 17280 256936 17332
rect 299480 17280 299532 17332
rect 382280 17280 382332 17332
rect 422300 17280 422352 17332
rect 458180 17280 458232 17332
rect 33140 17212 33192 17264
rect 219532 17212 219584 17264
rect 280804 17212 280856 17264
rect 369952 17212 370004 17264
rect 371240 17212 371292 17264
rect 426624 17212 426676 17264
rect 153752 16396 153804 16448
rect 293960 16396 294012 16448
rect 144736 16328 144788 16380
rect 288532 16328 288584 16380
rect 135352 16260 135404 16312
rect 281632 16260 281684 16312
rect 125600 16192 125652 16244
rect 276020 16192 276072 16244
rect 102140 16124 102192 16176
rect 254584 16124 254636 16176
rect 116400 16056 116452 16108
rect 270684 16056 270736 16108
rect 86408 15988 86460 16040
rect 250536 15988 250588 16040
rect 334624 15988 334676 16040
rect 404544 15988 404596 16040
rect 40224 15920 40276 15972
rect 223672 15920 223724 15972
rect 294512 15920 294564 15972
rect 379704 15920 379756 15972
rect 7656 15852 7708 15904
rect 204260 15852 204312 15904
rect 270776 15852 270828 15904
rect 365720 15852 365772 15904
rect 398932 15852 398984 15904
rect 444472 15852 444524 15904
rect 120632 14900 120684 14952
rect 273536 14900 273588 14952
rect 117320 14832 117372 14884
rect 271972 14832 272024 14884
rect 110512 14764 110564 14816
rect 266544 14764 266596 14816
rect 106464 14696 106516 14748
rect 265072 14696 265124 14748
rect 99840 14628 99892 14680
rect 260932 14628 260984 14680
rect 92480 14560 92532 14612
rect 256700 14560 256752 14612
rect 338672 14560 338724 14612
rect 407304 14560 407356 14612
rect 46664 14492 46716 14544
rect 227720 14492 227772 14544
rect 273904 14492 273956 14544
rect 353484 14492 353536 14544
rect 25320 14424 25372 14476
rect 215300 14424 215352 14476
rect 277952 14424 278004 14476
rect 369860 14424 369912 14476
rect 420184 14424 420236 14476
rect 456984 14424 457036 14476
rect 475752 14424 475804 14476
rect 491300 14424 491352 14476
rect 543924 14424 543976 14476
rect 562048 14424 562100 14476
rect 81624 13540 81676 13592
rect 214564 13540 214616 13592
rect 109040 13472 109092 13524
rect 266452 13472 266504 13524
rect 102232 13404 102284 13456
rect 262312 13404 262364 13456
rect 94688 13336 94740 13388
rect 258172 13336 258224 13388
rect 91560 13268 91612 13320
rect 255412 13268 255464 13320
rect 87512 13200 87564 13252
rect 252652 13200 252704 13252
rect 349160 13200 349212 13252
rect 412732 13200 412784 13252
rect 80888 13132 80940 13184
rect 248512 13132 248564 13184
rect 297456 13132 297508 13184
rect 374184 13132 374236 13184
rect 77392 13064 77444 13116
rect 247132 13064 247184 13116
rect 294696 13064 294748 13116
rect 378140 13064 378192 13116
rect 421012 13064 421064 13116
rect 456892 13064 456944 13116
rect 56784 12180 56836 12232
rect 234620 12180 234672 12232
rect 50160 12112 50212 12164
rect 230480 12112 230532 12164
rect 41880 12044 41932 12096
rect 224960 12044 225012 12096
rect 31944 11976 31996 12028
rect 219440 11976 219492 12028
rect 18604 11908 18656 11960
rect 208492 11908 208544 11960
rect 234620 11908 234672 11960
rect 343732 11908 343784 11960
rect 9680 11840 9732 11892
rect 205824 11840 205876 11892
rect 231032 11840 231084 11892
rect 340880 11840 340932 11892
rect 6000 11772 6052 11824
rect 202972 11772 203024 11824
rect 223580 11772 223632 11824
rect 336740 11772 336792 11824
rect 337384 11772 337436 11824
rect 397460 11772 397512 11824
rect 113824 11704 113876 11756
rect 200120 11704 200172 11756
rect 219992 11704 220044 11756
rect 333980 11704 334032 11756
rect 345296 11704 345348 11756
rect 411260 11704 411312 11756
rect 423864 11704 423916 11756
rect 459652 11704 459704 11756
rect 160100 11636 160152 11688
rect 161296 11636 161348 11688
rect 188528 10888 188580 10940
rect 314844 10888 314896 10940
rect 180984 10820 181036 10872
rect 310520 10820 310572 10872
rect 95792 10752 95844 10804
rect 175188 10752 175240 10804
rect 177580 10752 177632 10804
rect 307760 10752 307812 10804
rect 75000 10684 75052 10736
rect 170772 10684 170824 10736
rect 173900 10684 173952 10736
rect 306380 10684 306432 10736
rect 170312 10616 170364 10668
rect 303620 10616 303672 10668
rect 111616 10548 111668 10600
rect 267740 10548 267792 10600
rect 104072 10480 104124 10532
rect 263600 10480 263652 10532
rect 64328 10412 64380 10464
rect 233884 10412 233936 10464
rect 36728 10344 36780 10396
rect 222200 10344 222252 10396
rect 349252 10344 349304 10396
rect 414020 10344 414072 10396
rect 442632 10344 442684 10396
rect 470692 10344 470744 10396
rect 17960 10276 18012 10328
rect 211160 10276 211212 10328
rect 314752 10276 314804 10328
rect 391940 10276 391992 10328
rect 409144 10276 409196 10328
rect 449992 10276 450044 10328
rect 473912 10276 473964 10328
rect 490012 10276 490064 10328
rect 490104 10276 490156 10328
rect 499672 10276 499724 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 78588 9392 78640 9444
rect 247040 9392 247092 9444
rect 66720 9324 66772 9376
rect 240140 9324 240192 9376
rect 59636 9256 59688 9308
rect 236000 9256 236052 9308
rect 286600 9256 286652 9308
rect 375380 9256 375432 9308
rect 56048 9188 56100 9240
rect 233240 9188 233292 9240
rect 261760 9188 261812 9240
rect 360292 9188 360344 9240
rect 52552 9120 52604 9172
rect 231952 9120 232004 9172
rect 258264 9120 258316 9172
rect 357532 9120 357584 9172
rect 31300 9052 31352 9104
rect 218152 9052 218204 9104
rect 251180 9052 251232 9104
rect 353300 9052 353352 9104
rect 27712 8984 27764 9036
rect 216864 8984 216916 9036
rect 247592 8984 247644 9036
rect 350632 8984 350684 9036
rect 416688 8984 416740 9036
rect 454040 8984 454092 9036
rect 480536 8984 480588 9036
rect 494152 8984 494204 9036
rect 13544 8916 13596 8968
rect 207112 8916 207164 8968
rect 240508 8916 240560 8968
rect 346492 8916 346544 8968
rect 359924 8916 359976 8968
rect 419540 8916 419592 8968
rect 459192 8916 459244 8968
rect 480444 8916 480496 8968
rect 532700 8916 532752 8968
rect 543188 8916 543240 8968
rect 550732 8916 550784 8968
rect 572720 8916 572772 8968
rect 151912 8100 151964 8152
rect 292672 8100 292724 8152
rect 145932 8032 145984 8084
rect 287704 8032 287756 8084
rect 134156 7964 134208 8016
rect 281540 7964 281592 8016
rect 325608 7964 325660 8016
rect 398840 7964 398892 8016
rect 130568 7896 130620 7948
rect 278872 7896 278924 7948
rect 322112 7896 322164 7948
rect 396080 7896 396132 7948
rect 123484 7828 123536 7880
rect 274732 7828 274784 7880
rect 307944 7828 307996 7880
rect 387984 7828 388036 7880
rect 122288 7760 122340 7812
rect 274640 7760 274692 7812
rect 311440 7760 311492 7812
rect 390560 7760 390612 7812
rect 72608 7692 72660 7744
rect 244372 7692 244424 7744
rect 304356 7692 304408 7744
rect 386512 7692 386564 7744
rect 14740 7624 14792 7676
rect 208400 7624 208452 7676
rect 300768 7624 300820 7676
rect 383752 7624 383804 7676
rect 435548 7624 435600 7676
rect 466552 7624 466604 7676
rect 4068 7556 4120 7608
rect 201500 7556 201552 7608
rect 293684 7556 293736 7608
rect 379520 7556 379572 7608
rect 402520 7556 402572 7608
rect 445852 7556 445904 7608
rect 462780 7556 462832 7608
rect 483112 7556 483164 7608
rect 540980 7556 541032 7608
rect 558552 7556 558604 7608
rect 374092 7488 374144 7540
rect 375288 7488 375340 7540
rect 570604 6808 570656 6860
rect 580172 6808 580224 6860
rect 98644 6604 98696 6656
rect 259552 6604 259604 6656
rect 83280 6536 83332 6588
rect 249892 6536 249944 6588
rect 76196 6468 76248 6520
rect 246028 6468 246080 6520
rect 79692 6400 79744 6452
rect 248420 6400 248472 6452
rect 71504 6332 71556 6384
rect 242900 6332 242952 6384
rect 288992 6332 289044 6384
rect 376760 6332 376812 6384
rect 44272 6264 44324 6316
rect 226616 6264 226668 6316
rect 285404 6264 285456 6316
rect 374000 6264 374052 6316
rect 381176 6264 381228 6316
rect 433340 6264 433392 6316
rect 30104 6196 30156 6248
rect 218060 6196 218112 6248
rect 274824 6196 274876 6248
rect 367100 6196 367152 6248
rect 377680 6196 377732 6248
rect 430764 6196 430816 6248
rect 466276 6196 466328 6248
rect 484492 6196 484544 6248
rect 536932 6196 536984 6248
rect 551468 6196 551520 6248
rect 21824 6128 21876 6180
rect 212724 6128 212776 6180
rect 257068 6128 257120 6180
rect 357532 6128 357584 6180
rect 367008 6128 367060 6180
rect 423680 6128 423732 6180
rect 437940 6128 437992 6180
rect 467932 6128 467984 6180
rect 495900 6128 495952 6180
rect 503812 6128 503864 6180
rect 547972 6128 548024 6180
rect 569132 6128 569184 6180
rect 197912 5312 197964 5364
rect 320180 5312 320232 5364
rect 156604 5244 156656 5296
rect 284944 5244 284996 5296
rect 118792 5176 118844 5228
rect 267004 5176 267056 5228
rect 101036 5108 101088 5160
rect 260840 5108 260892 5160
rect 399024 5108 399076 5160
rect 443000 5108 443052 5160
rect 73804 5040 73856 5092
rect 244280 5040 244332 5092
rect 391848 5040 391900 5092
rect 438952 5040 439004 5092
rect 65524 4972 65576 5024
rect 238852 4972 238904 5024
rect 388260 4972 388312 5024
rect 437480 4972 437532 5024
rect 53748 4904 53800 4956
rect 231124 4904 231176 4956
rect 374184 4904 374236 4956
rect 427912 4904 427964 4956
rect 12348 4836 12400 4888
rect 207020 4836 207072 4888
rect 268844 4836 268896 4888
rect 364432 4836 364484 4888
rect 370596 4836 370648 4888
rect 426532 4836 426584 4888
rect 469864 4836 469916 4888
rect 487160 4836 487212 4888
rect 547144 4836 547196 4888
rect 547880 4836 547932 4888
rect 1676 4768 1728 4820
rect 200212 4768 200264 4820
rect 201500 4768 201552 4820
rect 322940 4768 322992 4820
rect 356336 4768 356388 4820
rect 418160 4768 418212 4820
rect 452108 4768 452160 4820
rect 476304 4768 476356 4820
rect 492312 4768 492364 4820
rect 501052 4768 501104 4820
rect 539692 4768 539744 4820
rect 554964 4768 555016 4820
rect 15936 4088 15988 4140
rect 18604 4088 18656 4140
rect 265348 4088 265400 4140
rect 269764 4088 269816 4140
rect 296076 4088 296128 4140
rect 297364 4088 297416 4140
rect 376484 4088 376536 4140
rect 377404 4088 377456 4140
rect 383568 4088 383620 4140
rect 384304 4088 384356 4140
rect 479340 4088 479392 4140
rect 482284 4088 482336 4140
rect 527272 4088 527324 4140
rect 527916 4088 527968 4140
rect 537484 4088 537536 4140
rect 549076 4088 549128 4140
rect 135260 4020 135312 4072
rect 136456 4020 136508 4072
rect 151820 4020 151872 4072
rect 153016 4020 153068 4072
rect 241704 4020 241756 4072
rect 250628 4020 250680 4072
rect 523040 4020 523092 4072
rect 529020 4020 529072 4072
rect 536840 4020 536892 4072
rect 550272 4020 550324 4072
rect 124680 3952 124732 4004
rect 169392 3952 169444 4004
rect 538220 3952 538272 4004
rect 553768 3952 553820 4004
rect 114008 3884 114060 3936
rect 188620 3884 188672 3936
rect 534724 3884 534776 3936
rect 538404 3884 538456 3936
rect 539600 3884 539652 3936
rect 556160 3884 556212 3936
rect 43076 3816 43128 3868
rect 173532 3816 173584 3868
rect 276020 3816 276072 3868
rect 278044 3816 278096 3868
rect 409880 3816 409932 3868
rect 410524 3816 410576 3868
rect 525800 3816 525852 3868
rect 532516 3816 532568 3868
rect 546500 3816 546552 3868
rect 566832 3816 566884 3868
rect 35992 3748 36044 3800
rect 177672 3748 177724 3800
rect 284300 3748 284352 3800
rect 297456 3748 297508 3800
rect 390652 3748 390704 3800
rect 438124 3748 438176 3800
rect 456892 3748 456944 3800
rect 464344 3748 464396 3800
rect 529940 3748 529992 3800
rect 28908 3680 28960 3732
rect 175096 3680 175148 3732
rect 260656 3680 260708 3732
rect 276664 3680 276716 3732
rect 298468 3680 298520 3732
rect 308404 3680 308456 3732
rect 316224 3680 316276 3732
rect 327724 3680 327776 3732
rect 372896 3680 372948 3732
rect 427820 3680 427872 3732
rect 443828 3680 443880 3732
rect 458824 3680 458876 3732
rect 465172 3680 465224 3732
rect 478236 3680 478288 3732
rect 527364 3680 527416 3732
rect 534908 3680 534960 3732
rect 20628 3612 20680 3664
rect 172152 3612 172204 3664
rect 225144 3612 225196 3664
rect 236736 3612 236788 3664
rect 252376 3612 252428 3664
rect 273904 3612 273956 3664
rect 277124 3612 277176 3664
rect 286324 3612 286376 3664
rect 19432 3544 19484 3596
rect 181444 3544 181496 3596
rect 193220 3544 193272 3596
rect 194416 3544 194468 3596
rect 196624 3544 196676 3596
rect 203892 3544 203944 3596
rect 204904 3544 204956 3596
rect 214472 3544 214524 3596
rect 218704 3544 218756 3596
rect 8760 3476 8812 3528
rect 10324 3476 10376 3528
rect 11152 3476 11204 3528
rect 213368 3476 213420 3528
rect 214748 3476 214800 3528
rect 215668 3476 215720 3528
rect 217324 3476 217376 3528
rect 218060 3476 218112 3528
rect 226984 3544 227036 3596
rect 228732 3544 228784 3596
rect 240784 3544 240836 3596
rect 244096 3544 244148 3596
rect 244924 3544 244976 3596
rect 222752 3476 222804 3528
rect 224316 3476 224368 3528
rect 226340 3476 226392 3528
rect 228364 3476 228416 3528
rect 235816 3476 235868 3528
rect 236644 3476 236696 3528
rect 250444 3544 250496 3596
rect 255872 3544 255924 3596
rect 264336 3544 264388 3596
rect 270040 3544 270092 3596
rect 294604 3612 294656 3664
rect 319720 3612 319772 3664
rect 330484 3612 330536 3664
rect 341064 3612 341116 3664
rect 356704 3612 356756 3664
rect 292580 3544 292632 3596
rect 294696 3544 294748 3596
rect 572 3408 624 3460
rect 113824 3408 113876 3460
rect 118700 3408 118752 3460
rect 119896 3408 119948 3460
rect 168380 3408 168432 3460
rect 169576 3408 169628 3460
rect 69020 3340 69072 3392
rect 69940 3340 69992 3392
rect 102140 3340 102192 3392
rect 103336 3340 103388 3392
rect 168380 3272 168432 3324
rect 229836 3272 229888 3324
rect 231216 3272 231268 3324
rect 232228 3340 232280 3392
rect 249984 3476 250036 3528
rect 254768 3476 254820 3528
rect 262956 3476 263008 3528
rect 290464 3476 290516 3528
rect 291384 3476 291436 3528
rect 304264 3544 304316 3596
rect 305552 3544 305604 3596
rect 318156 3544 318208 3596
rect 330392 3544 330444 3596
rect 297272 3476 297324 3528
rect 298744 3476 298796 3528
rect 301964 3476 302016 3528
rect 316684 3476 316736 3528
rect 323308 3476 323360 3528
rect 337384 3476 337436 3528
rect 337476 3476 337528 3528
rect 338764 3476 338816 3528
rect 340972 3476 341024 3528
rect 342168 3476 342220 3528
rect 348056 3544 348108 3596
rect 348424 3476 348476 3528
rect 349252 3476 349304 3528
rect 350448 3476 350500 3528
rect 355232 3544 355284 3596
rect 358728 3544 358780 3596
rect 360844 3544 360896 3596
rect 362316 3612 362368 3664
rect 420920 3612 420972 3664
rect 439136 3612 439188 3664
rect 440884 3612 440936 3664
rect 449808 3612 449860 3664
rect 467104 3612 467156 3664
rect 417056 3544 417108 3596
rect 423772 3544 423824 3596
rect 424968 3544 425020 3596
rect 426164 3544 426216 3596
rect 441620 3544 441672 3596
rect 237012 3340 237064 3392
rect 238024 3340 238076 3392
rect 302240 3408 302292 3460
rect 309048 3408 309100 3460
rect 311164 3408 311216 3460
rect 312636 3408 312688 3460
rect 324964 3408 325016 3460
rect 333888 3408 333940 3460
rect 404360 3408 404412 3460
rect 267740 3340 267792 3392
rect 271236 3340 271288 3392
rect 281908 3340 281960 3392
rect 285036 3340 285088 3392
rect 326804 3340 326856 3392
rect 334716 3340 334768 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 407120 3476 407172 3528
rect 408408 3476 408460 3528
rect 411904 3476 411956 3528
rect 447784 3544 447836 3596
rect 446220 3476 446272 3528
rect 447876 3476 447928 3528
rect 404820 3408 404872 3460
rect 446404 3408 446456 3460
rect 409880 3340 409932 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 441620 3340 441672 3392
rect 460940 3544 460992 3596
rect 461584 3544 461636 3596
rect 467472 3544 467524 3596
rect 468484 3544 468536 3596
rect 468668 3612 468720 3664
rect 480904 3612 480956 3664
rect 525984 3612 526036 3664
rect 533712 3612 533764 3664
rect 543740 3748 543792 3800
rect 563244 3748 563296 3800
rect 566464 3748 566516 3800
rect 570328 3748 570380 3800
rect 547972 3680 548024 3732
rect 568028 3680 568080 3732
rect 539600 3612 539652 3664
rect 550640 3612 550692 3664
rect 573916 3612 573968 3664
rect 456800 3476 456852 3528
rect 458088 3476 458140 3528
rect 450912 3408 450964 3460
rect 239312 3272 239364 3324
rect 240876 3272 240928 3324
rect 253480 3272 253532 3324
rect 258724 3272 258776 3324
rect 272432 3272 272484 3324
rect 276756 3272 276808 3324
rect 453304 3340 453356 3392
rect 471244 3476 471296 3528
rect 472256 3544 472308 3596
rect 486424 3544 486476 3596
rect 493508 3544 493560 3596
rect 500224 3544 500276 3596
rect 501788 3544 501840 3596
rect 506756 3544 506808 3596
rect 508872 3544 508924 3596
rect 510712 3544 510764 3596
rect 534172 3544 534224 3596
rect 545488 3544 545540 3596
rect 549260 3544 549312 3596
rect 571524 3544 571576 3596
rect 574744 3544 574796 3596
rect 576308 3544 576360 3596
rect 476764 3476 476816 3528
rect 481732 3476 481784 3528
rect 485044 3476 485096 3528
rect 506480 3476 506532 3528
rect 508504 3476 508556 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 518992 3476 519044 3528
rect 521844 3476 521896 3528
rect 524420 3476 524472 3528
rect 531320 3476 531372 3528
rect 534080 3476 534132 3528
rect 474004 3408 474056 3460
rect 486424 3408 486476 3460
rect 496912 3408 496964 3460
rect 521660 3408 521712 3460
rect 525432 3408 525484 3460
rect 527916 3408 527968 3460
rect 536104 3408 536156 3460
rect 538864 3476 538916 3528
rect 541992 3476 542044 3528
rect 553400 3476 553452 3528
rect 577412 3476 577464 3528
rect 578884 3476 578936 3528
rect 581000 3476 581052 3528
rect 546684 3408 546736 3460
rect 553492 3408 553544 3460
rect 578608 3408 578660 3460
rect 482836 3340 482888 3392
rect 487804 3340 487856 3392
rect 538312 3340 538364 3392
rect 552664 3340 552716 3392
rect 558184 3272 558236 3324
rect 559748 3272 559800 3324
rect 580264 3272 580316 3324
rect 582196 3272 582248 3324
rect 242900 3204 242952 3256
rect 247776 3204 247828 3256
rect 463976 3204 464028 3256
rect 467196 3204 467248 3256
rect 517612 3204 517664 3256
rect 519544 3204 519596 3256
rect 520464 3204 520516 3256
rect 524236 3204 524288 3256
rect 369400 3136 369452 3188
rect 370504 3136 370556 3188
rect 447416 3136 447468 3188
rect 450544 3136 450596 3188
rect 512460 3136 512512 3188
rect 513472 3136 513524 3188
rect 520372 3136 520424 3188
rect 523040 3136 523092 3188
rect 524512 3136 524564 3188
rect 530124 3136 530176 3188
rect 248788 3068 248840 3120
rect 257344 3068 257396 3120
rect 279516 3000 279568 3052
rect 280804 3000 280856 3052
rect 530584 3000 530636 3052
rect 537208 3000 537260 3052
rect 433248 2932 433300 2984
rect 434076 2932 434128 2984
rect 567844 2932 567896 2984
rect 575112 2932 575164 2984
rect 264152 2864 264204 2916
rect 268384 2864 268436 2916
rect 316040 960 316092 1012
rect 317328 960 317380 1012
<< metal2 >>
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 2962 619168 3018 619177
rect 2962 619103 3018 619112
rect 2976 618322 3004 619103
rect 2964 618316 3016 618322
rect 2964 618258 3016 618264
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 3160 579698 3188 579935
rect 3148 579692 3200 579698
rect 3148 579634 3200 579640
rect 3436 567194 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 571985 3556 658135
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3620 573374 3648 632023
rect 21364 618316 21416 618322
rect 21364 618258 21416 618264
rect 3698 606112 3754 606121
rect 3698 606047 3754 606056
rect 3712 576854 3740 606047
rect 3712 576826 3832 576854
rect 3608 573368 3660 573374
rect 3608 573310 3660 573316
rect 3514 571976 3570 571985
rect 3514 571911 3570 571920
rect 3436 567166 3556 567194
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3528 565146 3556 567166
rect 3516 565140 3568 565146
rect 3516 565082 3568 565088
rect 3804 563718 3832 576826
rect 3792 563712 3844 563718
rect 3792 563654 3844 563660
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3436 450945 3464 527847
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 18604 514820 18656 514826
rect 3516 514762 3568 514768
rect 18604 514762 18656 514768
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3528 475590 3556 475623
rect 3516 475584 3568 475590
rect 3516 475526 3568 475532
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3422 450936 3478 450945
rect 3422 450871 3478 450880
rect 18616 450566 18644 514762
rect 21376 450673 21404 618258
rect 21362 450664 21418 450673
rect 21362 450599 21418 450608
rect 18604 450560 18656 450566
rect 23492 450537 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40512 700369 40540 703520
rect 72988 700398 73016 703520
rect 89180 700505 89208 703520
rect 89166 700496 89222 700505
rect 89166 700431 89222 700440
rect 72976 700392 73028 700398
rect 40498 700360 40554 700369
rect 72976 700334 73028 700340
rect 40498 700295 40554 700304
rect 105464 698970 105492 703520
rect 137848 700466 137876 703520
rect 154132 700641 154160 703520
rect 154118 700632 154174 700641
rect 154118 700567 154174 700576
rect 170324 700534 170352 703520
rect 170312 700528 170364 700534
rect 170312 700470 170364 700476
rect 177304 700528 177356 700534
rect 177304 700470 177356 700476
rect 137836 700460 137888 700466
rect 137836 700402 137888 700408
rect 105452 698964 105504 698970
rect 105452 698906 105504 698912
rect 28724 675028 28776 675034
rect 28724 674970 28776 674976
rect 28632 674960 28684 674966
rect 28632 674902 28684 674908
rect 28170 669216 28226 669225
rect 28170 669151 28226 669160
rect 27434 609376 27490 609385
rect 27434 609311 27490 609320
rect 27342 607744 27398 607753
rect 27342 607679 27398 607688
rect 27158 604888 27214 604897
rect 27158 604823 27214 604832
rect 27066 494320 27122 494329
rect 27066 494255 27122 494264
rect 18604 450502 18656 450508
rect 23478 450528 23534 450537
rect 23478 450463 23534 450472
rect 3332 450016 3384 450022
rect 3332 449958 3384 449964
rect 3344 449585 3372 449958
rect 3516 449948 3568 449954
rect 3516 449890 3568 449896
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3528 423609 3556 449890
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3424 411256 3476 411262
rect 3424 411198 3476 411204
rect 3436 410553 3464 411198
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3240 398812 3292 398818
rect 3240 398754 3292 398760
rect 3252 397497 3280 398754
rect 3238 397488 3294 397497
rect 3238 397423 3294 397432
rect 27080 382401 27108 494255
rect 27172 494057 27200 604823
rect 27250 603664 27306 603673
rect 27250 603599 27306 603608
rect 27158 494048 27214 494057
rect 27158 493983 27214 493992
rect 27264 491609 27292 603599
rect 27356 495689 27384 607679
rect 27448 497321 27476 609311
rect 27526 606384 27582 606393
rect 27526 606319 27582 606328
rect 27434 497312 27490 497321
rect 27434 497247 27490 497256
rect 27342 495680 27398 495689
rect 27342 495615 27398 495624
rect 27250 491600 27306 491609
rect 27250 491535 27306 491544
rect 27158 386336 27214 386345
rect 27158 386271 27214 386280
rect 27172 385393 27200 386271
rect 27158 385384 27214 385393
rect 27158 385319 27214 385328
rect 27066 382392 27122 382401
rect 27066 382327 27122 382336
rect 27066 379808 27122 379817
rect 27066 379743 27122 379752
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 365702 3464 371311
rect 3424 365696 3476 365702
rect 3424 365638 3476 365644
rect 3424 365152 3476 365158
rect 3424 365094 3476 365100
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3332 137964 3384 137970
rect 3332 137906 3384 137912
rect 3344 136785 3372 137906
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3436 32473 3464 365094
rect 3608 365084 3660 365090
rect 3608 365026 3660 365032
rect 3516 365016 3568 365022
rect 3516 364958 3568 364964
rect 3528 58585 3556 364958
rect 3620 201929 3648 365026
rect 3976 340196 4028 340202
rect 3976 340138 4028 340144
rect 3698 340096 3754 340105
rect 3698 340031 3754 340040
rect 3712 254153 3740 340031
rect 3884 338836 3936 338842
rect 3884 338778 3936 338784
rect 3792 338768 3844 338774
rect 3792 338710 3844 338716
rect 3804 267209 3832 338710
rect 3896 293185 3924 338778
rect 3988 306241 4016 340138
rect 4068 338904 4120 338910
rect 4068 338846 4120 338852
rect 4080 319297 4108 338846
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 3974 306232 4030 306241
rect 3974 306167 4030 306176
rect 3882 293176 3938 293185
rect 3882 293111 3938 293120
rect 27080 269113 27108 379743
rect 27172 273329 27200 385319
rect 27264 379681 27292 491535
rect 27356 383761 27384 495615
rect 27448 386345 27476 497247
rect 27540 494329 27568 606319
rect 27526 494320 27582 494329
rect 27526 494255 27582 494264
rect 27526 494048 27582 494057
rect 27526 493983 27582 493992
rect 27540 492833 27568 493983
rect 27526 492824 27582 492833
rect 27526 492759 27582 492768
rect 27434 386336 27490 386345
rect 27434 386271 27490 386280
rect 27342 383752 27398 383761
rect 27342 383687 27398 383696
rect 27250 379672 27306 379681
rect 27250 379607 27306 379616
rect 27158 273320 27214 273329
rect 27158 273255 27214 273264
rect 27066 269104 27122 269113
rect 27066 269039 27122 269048
rect 3790 267200 3846 267209
rect 3790 267135 3846 267144
rect 3698 254144 3754 254153
rect 3698 254079 3754 254088
rect 27172 252657 27200 273255
rect 27356 271697 27384 383687
rect 27434 382392 27490 382401
rect 27434 382327 27490 382336
rect 27342 271688 27398 271697
rect 27342 271623 27398 271632
rect 27250 269104 27306 269113
rect 27250 269039 27306 269048
rect 27158 252648 27214 252657
rect 27158 252583 27214 252592
rect 27068 252544 27120 252550
rect 26974 252512 27030 252521
rect 27068 252486 27120 252492
rect 26974 252447 27030 252456
rect 26988 251569 27016 252447
rect 26974 251560 27030 251569
rect 26974 251495 27030 251504
rect 3700 228404 3752 228410
rect 3700 228346 3752 228352
rect 3606 201920 3662 201929
rect 3606 201855 3662 201864
rect 3712 149841 3740 228346
rect 3974 227080 4030 227089
rect 3884 227044 3936 227050
rect 3974 227015 4030 227024
rect 3884 226986 3936 226992
rect 3790 226944 3846 226953
rect 3790 226879 3846 226888
rect 3804 162897 3832 226879
rect 3896 188873 3924 226986
rect 3988 214985 4016 227015
rect 3974 214976 4030 214985
rect 3974 214911 4030 214920
rect 3882 188864 3938 188873
rect 3882 188799 3938 188808
rect 3790 162888 3846 162897
rect 3790 162823 3846 162832
rect 26988 158409 27016 251495
rect 26974 158400 27030 158409
rect 26974 158335 27030 158344
rect 27080 156913 27108 252486
rect 27172 161401 27200 252583
rect 27264 252550 27292 269039
rect 27356 253881 27384 271623
rect 27448 270337 27476 382327
rect 27540 380905 27568 492759
rect 27526 380896 27582 380905
rect 27526 380831 27582 380840
rect 27540 379817 27568 380831
rect 27526 379808 27582 379817
rect 27526 379743 27582 379752
rect 27526 379672 27582 379681
rect 27526 379607 27582 379616
rect 27434 270328 27490 270337
rect 27434 270263 27490 270272
rect 27342 253872 27398 253881
rect 27342 253807 27398 253816
rect 27252 252544 27304 252550
rect 27252 252486 27304 252492
rect 27158 161392 27214 161401
rect 27158 161327 27214 161336
rect 27172 160177 27200 161327
rect 27158 160168 27214 160177
rect 27158 160103 27214 160112
rect 27356 159769 27384 253807
rect 27448 252521 27476 270263
rect 27540 267617 27568 379607
rect 27526 267608 27582 267617
rect 27526 267543 27582 267552
rect 27540 253910 27568 267543
rect 27528 253904 27580 253910
rect 27528 253846 27580 253852
rect 27434 252512 27490 252521
rect 27434 252447 27490 252456
rect 27434 160168 27490 160177
rect 27434 160103 27490 160112
rect 27342 159760 27398 159769
rect 27342 159695 27398 159704
rect 27250 158400 27306 158409
rect 27250 158335 27306 158344
rect 27066 156904 27122 156913
rect 27066 156839 27122 156848
rect 3698 149832 3754 149841
rect 3698 149767 3754 149776
rect 3792 115388 3844 115394
rect 3792 115330 3844 115336
rect 3608 115252 3660 115258
rect 3608 115194 3660 115200
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3620 45529 3648 115194
rect 3700 113892 3752 113898
rect 3700 113834 3752 113840
rect 3712 71641 3740 113834
rect 3804 84697 3832 115330
rect 3884 115320 3936 115326
rect 3884 115262 3936 115268
rect 3896 97617 3924 115262
rect 4068 113824 4120 113830
rect 4068 113766 4120 113772
rect 4080 110673 4108 113766
rect 4066 110664 4122 110673
rect 4066 110599 4122 110608
rect 3882 97608 3938 97617
rect 3882 97543 3938 97552
rect 3790 84688 3846 84697
rect 3790 84623 3846 84632
rect 3698 71632 3754 71641
rect 3698 71567 3754 71576
rect 3606 45520 3662 45529
rect 3606 45455 3662 45464
rect 27080 44985 27108 156839
rect 27158 155680 27214 155689
rect 27158 155615 27214 155624
rect 27066 44976 27122 44985
rect 27066 44911 27122 44920
rect 27172 43761 27200 155615
rect 27264 46481 27292 158335
rect 27356 47841 27384 159695
rect 27448 49473 27476 160103
rect 27540 155689 27568 253846
rect 28184 245614 28212 669151
rect 28540 586628 28592 586634
rect 28540 586570 28592 586576
rect 28448 586560 28500 586566
rect 28448 586502 28500 586508
rect 28264 553444 28316 553450
rect 28264 553386 28316 553392
rect 28276 450809 28304 553386
rect 28460 475318 28488 586502
rect 28552 475522 28580 586570
rect 28644 562018 28672 674902
rect 28736 562630 28764 674970
rect 34520 674960 34572 674966
rect 34518 674928 34520 674937
rect 46204 674960 46256 674966
rect 34572 674928 34574 674937
rect 28816 674892 28868 674898
rect 34518 674863 34574 674872
rect 46202 674928 46204 674937
rect 46256 674928 46258 674937
rect 46202 674863 46258 674872
rect 46938 674928 46994 674937
rect 46938 674863 46940 674872
rect 28816 674834 28868 674840
rect 46992 674863 46994 674872
rect 46940 674834 46992 674840
rect 28724 562624 28776 562630
rect 28724 562566 28776 562572
rect 28828 562358 28856 674834
rect 169022 626920 169078 626929
rect 169022 626855 169078 626864
rect 168562 618216 168618 618225
rect 168562 618151 168618 618160
rect 43074 587888 43130 587897
rect 43074 587823 43130 587832
rect 43534 587888 43590 587897
rect 43534 587823 43590 587832
rect 60646 587888 60702 587897
rect 60646 587823 60702 587832
rect 62946 587888 63002 587897
rect 62946 587823 63002 587832
rect 68926 587888 68982 587897
rect 68926 587823 68982 587832
rect 74446 587888 74502 587897
rect 74446 587823 74502 587832
rect 83830 587888 83886 587897
rect 83830 587823 83886 587832
rect 86406 587888 86462 587897
rect 86406 587823 86462 587832
rect 88246 587888 88302 587897
rect 88246 587823 88302 587832
rect 95238 587888 95294 587897
rect 95238 587823 95294 587832
rect 99194 587888 99250 587897
rect 99194 587823 99250 587832
rect 100574 587888 100630 587897
rect 100574 587823 100630 587832
rect 103150 587888 103206 587897
rect 103150 587823 103206 587832
rect 105082 587888 105138 587897
rect 105082 587823 105138 587832
rect 106278 587888 106334 587897
rect 106278 587823 106334 587832
rect 107750 587888 107806 587897
rect 107750 587823 107806 587832
rect 109498 587888 109554 587897
rect 109498 587823 109554 587832
rect 110510 587888 110566 587897
rect 110510 587823 110566 587832
rect 111614 587888 111670 587897
rect 111614 587823 111670 587832
rect 112534 587888 112590 587897
rect 112534 587823 112590 587832
rect 113086 587888 113142 587897
rect 113086 587823 113142 587832
rect 113822 587888 113878 587897
rect 113822 587823 113878 587832
rect 114834 587888 114890 587897
rect 114834 587823 114890 587832
rect 117134 587888 117190 587897
rect 117134 587823 117190 587832
rect 119802 587888 119858 587897
rect 119802 587823 119858 587832
rect 120262 587888 120318 587897
rect 120262 587823 120318 587832
rect 120538 587888 120594 587897
rect 120538 587823 120594 587832
rect 122654 587888 122710 587897
rect 122654 587823 122710 587832
rect 122838 587888 122894 587897
rect 122838 587823 122894 587832
rect 125046 587888 125102 587897
rect 125046 587823 125102 587832
rect 126886 587888 126942 587897
rect 126886 587823 126942 587832
rect 129370 587888 129426 587897
rect 129370 587823 129426 587832
rect 129646 587888 129702 587897
rect 129646 587823 129702 587832
rect 130566 587888 130622 587897
rect 130566 587823 130622 587832
rect 131118 587888 131174 587897
rect 131118 587823 131174 587832
rect 132590 587888 132646 587897
rect 132590 587823 132646 587832
rect 133142 587888 133198 587897
rect 133142 587823 133198 587832
rect 136454 587888 136510 587897
rect 136454 587823 136510 587832
rect 137926 587888 137982 587897
rect 137926 587823 137982 587832
rect 139306 587888 139362 587897
rect 139306 587823 139362 587832
rect 140134 587888 140190 587897
rect 140134 587823 140190 587832
rect 142710 587888 142766 587897
rect 142710 587823 142766 587832
rect 143446 587888 143502 587897
rect 143446 587823 143502 587832
rect 147678 587888 147734 587897
rect 147678 587823 147734 587832
rect 149518 587888 149574 587897
rect 149518 587823 149574 587832
rect 150714 587888 150770 587897
rect 150714 587823 150770 587832
rect 43088 586634 43116 587823
rect 43076 586628 43128 586634
rect 43076 586570 43128 586576
rect 43548 586566 43576 587823
rect 43536 586560 43588 586566
rect 43536 586502 43588 586508
rect 29736 563168 29788 563174
rect 29736 563110 29788 563116
rect 35714 563136 35770 563145
rect 29644 563100 29696 563106
rect 29644 563042 29696 563048
rect 28816 562352 28868 562358
rect 28816 562294 28868 562300
rect 29656 562018 29684 563042
rect 29748 562630 29776 563110
rect 35714 563071 35716 563080
rect 35768 563071 35770 563080
rect 46754 563136 46810 563145
rect 46754 563071 46756 563080
rect 35716 563042 35768 563048
rect 46808 563071 46810 563080
rect 46756 563042 46808 563048
rect 29736 562624 29788 562630
rect 29736 562566 29788 562572
rect 28632 562012 28684 562018
rect 28632 561954 28684 561960
rect 29644 562012 29696 562018
rect 29644 561954 29696 561960
rect 28814 557152 28870 557161
rect 28814 557087 28870 557096
rect 28724 501016 28776 501022
rect 28724 500958 28776 500964
rect 28540 475516 28592 475522
rect 28540 475458 28592 475464
rect 28448 475312 28500 475318
rect 28448 475254 28500 475260
rect 28460 474706 28488 475254
rect 28448 474700 28500 474706
rect 28448 474642 28500 474648
rect 28552 470594 28580 475458
rect 28552 470566 28672 470594
rect 28540 451988 28592 451994
rect 28540 451930 28592 451936
rect 28262 450800 28318 450809
rect 28262 450735 28318 450744
rect 28356 450152 28408 450158
rect 28356 450094 28408 450100
rect 28368 398818 28396 450094
rect 28448 450084 28500 450090
rect 28448 450026 28500 450032
rect 28460 411262 28488 450026
rect 28448 411256 28500 411262
rect 28448 411198 28500 411204
rect 28356 398812 28408 398818
rect 28356 398754 28408 398760
rect 28552 339590 28580 451930
rect 28644 363730 28672 470566
rect 28736 450634 28764 500958
rect 28724 450628 28776 450634
rect 28724 450570 28776 450576
rect 28722 445224 28778 445233
rect 28722 445159 28778 445168
rect 28632 363724 28684 363730
rect 28632 363666 28684 363672
rect 28540 339584 28592 339590
rect 28540 339526 28592 339532
rect 28552 335354 28580 339526
rect 28460 335326 28580 335354
rect 28356 253224 28408 253230
rect 28356 253166 28408 253172
rect 28172 245608 28224 245614
rect 28172 245550 28224 245556
rect 27526 155680 27582 155689
rect 27526 155615 27582 155624
rect 28368 138582 28396 253166
rect 28460 252550 28488 335326
rect 28538 333160 28594 333169
rect 28538 333095 28594 333104
rect 28448 252544 28500 252550
rect 28448 252486 28500 252492
rect 28552 244254 28580 333095
rect 28644 252385 28672 363666
rect 28630 252376 28686 252385
rect 28630 252311 28686 252320
rect 28540 244248 28592 244254
rect 28540 244190 28592 244196
rect 28448 236700 28500 236706
rect 28448 236642 28500 236648
rect 28460 221241 28488 236642
rect 28540 229152 28592 229158
rect 28540 229094 28592 229100
rect 28446 221232 28502 221241
rect 28446 221167 28502 221176
rect 28356 138576 28408 138582
rect 28356 138518 28408 138524
rect 28552 117162 28580 229094
rect 28644 138718 28672 252311
rect 28736 242894 28764 445159
rect 28828 247042 28856 557087
rect 29656 475386 29684 561954
rect 29644 475380 29696 475386
rect 29644 475322 29696 475328
rect 29644 474700 29696 474706
rect 29644 474642 29696 474648
rect 29552 452600 29604 452606
rect 29552 452542 29604 452548
rect 29564 451926 29592 452542
rect 29552 451920 29604 451926
rect 29552 451862 29604 451868
rect 29460 362976 29512 362982
rect 29460 362918 29512 362924
rect 29472 253230 29500 362918
rect 29564 340270 29592 451862
rect 29656 363866 29684 474642
rect 29748 452606 29776 562566
rect 60660 562358 60688 587823
rect 62960 584458 62988 587823
rect 64878 586528 64934 586537
rect 64878 586463 64934 586472
rect 62948 584452 63000 584458
rect 62948 584394 63000 584400
rect 64892 580310 64920 586463
rect 64880 580304 64932 580310
rect 64880 580246 64932 580252
rect 68940 573442 68968 587823
rect 71686 586392 71742 586401
rect 71686 586327 71742 586336
rect 68928 573436 68980 573442
rect 68928 573378 68980 573384
rect 71700 572014 71728 586327
rect 71688 572008 71740 572014
rect 71688 571950 71740 571956
rect 74460 566506 74488 587823
rect 75826 586392 75882 586401
rect 75826 586327 75882 586336
rect 78586 586392 78642 586401
rect 78586 586327 78642 586336
rect 81346 586392 81402 586401
rect 81346 586327 81402 586336
rect 74448 566500 74500 566506
rect 74448 566442 74500 566448
rect 75840 565214 75868 586327
rect 75828 565208 75880 565214
rect 75828 565150 75880 565156
rect 78600 563786 78628 586327
rect 81360 574802 81388 586327
rect 83844 578950 83872 587823
rect 83832 578944 83884 578950
rect 83832 578886 83884 578892
rect 86420 577522 86448 587823
rect 86408 577516 86460 577522
rect 86408 577458 86460 577464
rect 81348 574796 81400 574802
rect 81348 574738 81400 574744
rect 88260 570654 88288 587823
rect 91006 586392 91062 586401
rect 91006 586327 91062 586336
rect 93766 586392 93822 586401
rect 93766 586327 93822 586336
rect 88248 570648 88300 570654
rect 88248 570590 88300 570596
rect 91020 569226 91048 586327
rect 93780 576162 93808 586327
rect 95252 581670 95280 587823
rect 99208 587450 99236 587823
rect 99196 587444 99248 587450
rect 99196 587386 99248 587392
rect 100588 586702 100616 587823
rect 100576 586696 100628 586702
rect 100576 586638 100628 586644
rect 103164 586634 103192 587823
rect 103152 586628 103204 586634
rect 103152 586570 103204 586576
rect 105096 585818 105124 587823
rect 105084 585812 105136 585818
rect 105084 585754 105136 585760
rect 95240 581664 95292 581670
rect 106292 581641 106320 587823
rect 107764 581777 107792 587823
rect 108946 586392 109002 586401
rect 108946 586327 109002 586336
rect 107750 581768 107806 581777
rect 107750 581703 107806 581712
rect 95240 581606 95292 581612
rect 106278 581632 106334 581641
rect 106278 581567 106334 581576
rect 93768 576156 93820 576162
rect 93768 576098 93820 576104
rect 91008 569220 91060 569226
rect 91008 569162 91060 569168
rect 108960 567866 108988 586327
rect 109512 584594 109540 587823
rect 109500 584588 109552 584594
rect 109500 584530 109552 584536
rect 110524 584526 110552 587823
rect 110512 584520 110564 584526
rect 111628 584497 111656 587823
rect 110512 584462 110564 584468
rect 111614 584488 111670 584497
rect 111614 584423 111670 584432
rect 112548 584361 112576 587823
rect 112534 584352 112590 584361
rect 112534 584287 112590 584296
rect 113100 576230 113128 587823
rect 113836 584662 113864 587823
rect 114374 587752 114430 587761
rect 114374 587687 114430 587696
rect 114558 587752 114614 587761
rect 114558 587687 114614 587696
rect 113824 584656 113876 584662
rect 114388 584633 114416 587687
rect 113824 584598 113876 584604
rect 114374 584624 114430 584633
rect 114374 584559 114430 584568
rect 114572 577590 114600 587687
rect 114848 584730 114876 587823
rect 117148 584798 117176 587823
rect 118606 586392 118662 586401
rect 118606 586327 118662 586336
rect 117136 584792 117188 584798
rect 117136 584734 117188 584740
rect 114836 584724 114888 584730
rect 114836 584666 114888 584672
rect 114560 577584 114612 577590
rect 114560 577526 114612 577532
rect 113088 576224 113140 576230
rect 113088 576166 113140 576172
rect 118620 574870 118648 586327
rect 119816 584769 119844 587823
rect 120170 587752 120226 587761
rect 120170 587687 120226 587696
rect 119802 584760 119858 584769
rect 119802 584695 119858 584704
rect 120184 579018 120212 587687
rect 120276 584905 120304 587823
rect 120552 585070 120580 587823
rect 120540 585064 120592 585070
rect 120540 585006 120592 585012
rect 120262 584896 120318 584905
rect 122668 584866 122696 587823
rect 120262 584831 120318 584840
rect 122656 584860 122708 584866
rect 122656 584802 122708 584808
rect 122852 581738 122880 587823
rect 125060 585002 125088 587823
rect 126900 586770 126928 587823
rect 126888 586764 126940 586770
rect 126888 586706 126940 586712
rect 125506 586392 125562 586401
rect 125506 586327 125562 586336
rect 128266 586392 128322 586401
rect 128266 586327 128322 586336
rect 125048 584996 125100 585002
rect 125048 584938 125100 584944
rect 122840 581732 122892 581738
rect 122840 581674 122892 581680
rect 120172 579012 120224 579018
rect 120172 578954 120224 578960
rect 118608 574864 118660 574870
rect 118608 574806 118660 574812
rect 125520 570722 125548 586327
rect 125508 570716 125560 570722
rect 125508 570658 125560 570664
rect 128280 569498 128308 586327
rect 129384 584934 129412 587823
rect 129660 586838 129688 587823
rect 129648 586832 129700 586838
rect 129648 586774 129700 586780
rect 130580 585138 130608 587823
rect 131026 587752 131082 587761
rect 131026 587687 131082 587696
rect 130568 585132 130620 585138
rect 130568 585074 130620 585080
rect 129372 584928 129424 584934
rect 129372 584870 129424 584876
rect 128268 569492 128320 569498
rect 128268 569434 128320 569440
rect 131040 567934 131068 587687
rect 131132 584390 131160 587823
rect 131120 584384 131172 584390
rect 131120 584326 131172 584332
rect 132604 583030 132632 587823
rect 133156 586906 133184 587823
rect 133144 586900 133196 586906
rect 133144 586842 133196 586848
rect 136468 584322 136496 587823
rect 137940 587110 137968 587823
rect 137928 587104 137980 587110
rect 136546 587072 136602 587081
rect 137928 587046 137980 587052
rect 139030 587072 139086 587081
rect 136546 587007 136602 587016
rect 139030 587007 139032 587016
rect 136560 586974 136588 587007
rect 139084 587007 139086 587016
rect 139032 586978 139084 586984
rect 136548 586968 136600 586974
rect 136548 586910 136600 586916
rect 139320 585886 139348 587823
rect 140148 587178 140176 587823
rect 142724 587246 142752 587823
rect 143460 587314 143488 587823
rect 143448 587308 143500 587314
rect 143448 587250 143500 587256
rect 142712 587240 142764 587246
rect 142712 587182 142764 587188
rect 140136 587172 140188 587178
rect 140136 587114 140188 587120
rect 142066 586392 142122 586401
rect 142066 586327 142122 586336
rect 139308 585880 139360 585886
rect 139308 585822 139360 585828
rect 136456 584316 136508 584322
rect 136456 584258 136508 584264
rect 132592 583024 132644 583030
rect 132592 582966 132644 582972
rect 131028 567928 131080 567934
rect 131028 567870 131080 567876
rect 108948 567860 109000 567866
rect 108948 567802 109000 567808
rect 142080 563854 142108 586327
rect 147692 584254 147720 587823
rect 149532 587382 149560 587823
rect 149520 587376 149572 587382
rect 149520 587318 149572 587324
rect 150728 586566 150756 587823
rect 167000 587308 167052 587314
rect 167000 587250 167052 587256
rect 150716 586560 150768 586566
rect 150716 586502 150768 586508
rect 147680 584248 147732 584254
rect 147680 584190 147732 584196
rect 142068 563848 142120 563854
rect 142068 563790 142120 563796
rect 78588 563780 78640 563786
rect 78588 563722 78640 563728
rect 29828 562352 29880 562358
rect 29828 562294 29880 562300
rect 48044 562352 48096 562358
rect 48044 562294 48096 562300
rect 60648 562352 60700 562358
rect 60648 562294 60700 562300
rect 29736 452600 29788 452606
rect 29736 452542 29788 452548
rect 29840 451246 29868 562294
rect 48056 561785 48084 562294
rect 48042 561776 48098 561785
rect 48042 561711 48098 561720
rect 115478 477864 115534 477873
rect 115478 477799 115534 477808
rect 122654 477864 122710 477873
rect 122654 477799 122710 477808
rect 63406 476096 63462 476105
rect 63406 476031 63462 476040
rect 66166 476096 66222 476105
rect 66166 476031 66222 476040
rect 84106 476096 84162 476105
rect 84106 476031 84162 476040
rect 86866 476096 86922 476105
rect 86866 476031 86922 476040
rect 96526 476096 96582 476105
rect 96526 476031 96582 476040
rect 106186 476096 106242 476105
rect 106186 476031 106242 476040
rect 112994 476096 113050 476105
rect 112994 476031 113050 476040
rect 42798 475552 42854 475561
rect 42798 475487 42800 475496
rect 42852 475487 42854 475496
rect 42800 475458 42852 475464
rect 42798 475416 42854 475425
rect 34520 475380 34572 475386
rect 42798 475351 42800 475360
rect 34520 475322 34572 475328
rect 42852 475351 42854 475360
rect 42800 475322 42852 475328
rect 34532 452577 34560 475322
rect 60646 474872 60702 474881
rect 60646 474807 60648 474816
rect 60700 474807 60702 474816
rect 60648 474778 60700 474784
rect 63420 456074 63448 476031
rect 63408 456068 63460 456074
rect 63408 456010 63460 456016
rect 34518 452568 34574 452577
rect 34518 452503 34574 452512
rect 34532 451994 34560 452503
rect 66180 451994 66208 476031
rect 68926 474872 68982 474881
rect 68926 474807 68982 474816
rect 71686 474872 71742 474881
rect 71686 474807 71742 474816
rect 74446 474872 74502 474881
rect 74446 474807 74502 474816
rect 75826 474872 75882 474881
rect 75826 474807 75882 474816
rect 78586 474872 78642 474881
rect 78586 474807 78642 474816
rect 81346 474872 81402 474881
rect 81346 474807 81402 474816
rect 68940 464370 68968 474807
rect 68928 464364 68980 464370
rect 68928 464306 68980 464312
rect 71700 454714 71728 474807
rect 74460 465730 74488 474807
rect 75840 468518 75868 474807
rect 75828 468512 75880 468518
rect 75828 468454 75880 468460
rect 78600 467158 78628 474807
rect 78588 467152 78640 467158
rect 78588 467094 78640 467100
rect 74448 465724 74500 465730
rect 74448 465666 74500 465672
rect 81360 461650 81388 474807
rect 84120 469878 84148 476031
rect 86880 471306 86908 476031
rect 88246 474872 88302 474881
rect 88246 474807 88302 474816
rect 91006 474872 91062 474881
rect 91006 474807 91062 474816
rect 93766 474872 93822 474881
rect 93766 474807 93822 474816
rect 86868 471300 86920 471306
rect 86868 471242 86920 471248
rect 84108 469872 84160 469878
rect 84108 469814 84160 469820
rect 81348 461644 81400 461650
rect 81348 461586 81400 461592
rect 88260 460222 88288 474807
rect 88248 460216 88300 460222
rect 88248 460158 88300 460164
rect 91020 458862 91048 474807
rect 93780 472666 93808 474807
rect 96540 474026 96568 476031
rect 99286 474872 99342 474881
rect 99286 474807 99342 474816
rect 100666 474872 100722 474881
rect 100666 474807 100722 474816
rect 103426 474872 103482 474881
rect 103426 474807 103482 474816
rect 96528 474020 96580 474026
rect 96528 473962 96580 473968
rect 93768 472660 93820 472666
rect 93768 472602 93820 472608
rect 91008 458856 91060 458862
rect 91008 458798 91060 458804
rect 99300 457502 99328 474807
rect 100680 464438 100708 474807
rect 100668 464432 100720 464438
rect 100668 464374 100720 464380
rect 103440 461718 103468 474807
rect 106200 467226 106228 476031
rect 108854 475008 108910 475017
rect 108854 474943 108910 474952
rect 110326 475008 110382 475017
rect 110326 474943 110328 474952
rect 107566 474872 107622 474881
rect 107566 474807 107622 474816
rect 106188 467220 106240 467226
rect 106188 467162 106240 467168
rect 103428 461712 103480 461718
rect 103428 461654 103480 461660
rect 99288 457496 99340 457502
rect 99288 457438 99340 457444
rect 107580 456249 107608 474807
rect 108868 468586 108896 474943
rect 110380 474943 110382 474952
rect 111614 475008 111670 475017
rect 111614 474943 111670 474952
rect 110328 474914 110380 474920
rect 108946 474872 109002 474881
rect 108946 474807 109002 474816
rect 108856 468580 108908 468586
rect 108856 468522 108908 468528
rect 107566 456240 107622 456249
rect 107566 456175 107622 456184
rect 108960 454753 108988 474807
rect 111628 469946 111656 474943
rect 111706 474872 111762 474881
rect 111706 474807 111762 474816
rect 111616 469940 111668 469946
rect 111616 469882 111668 469888
rect 111720 456113 111748 474807
rect 113008 471374 113036 476031
rect 115492 475046 115520 477799
rect 121182 475552 121238 475561
rect 121182 475487 121238 475496
rect 115480 475040 115532 475046
rect 114374 475008 114430 475017
rect 115480 474982 115532 474988
rect 118606 475008 118662 475017
rect 114374 474943 114430 474952
rect 118606 474943 118662 474952
rect 113086 474872 113142 474881
rect 113086 474807 113142 474816
rect 112996 471368 113048 471374
rect 112996 471310 113048 471316
rect 111706 456104 111762 456113
rect 111706 456039 111762 456048
rect 113100 454850 113128 474807
rect 113088 454844 113140 454850
rect 113088 454786 113140 454792
rect 114388 454782 114416 474943
rect 114466 474872 114522 474881
rect 114466 474807 114522 474816
rect 115754 474872 115810 474881
rect 115754 474807 115810 474816
rect 117226 474872 117282 474881
rect 117226 474807 117282 474816
rect 118514 474872 118570 474881
rect 118514 474807 118570 474816
rect 114376 454776 114428 454782
rect 108946 454744 109002 454753
rect 71688 454708 71740 454714
rect 114376 454718 114428 454724
rect 108946 454679 109002 454688
rect 71688 454650 71740 454656
rect 114480 453490 114508 474807
rect 115768 467294 115796 474807
rect 115756 467288 115808 467294
rect 115756 467230 115808 467236
rect 117240 453626 117268 474807
rect 118528 458930 118556 474807
rect 118516 458924 118568 458930
rect 118516 458866 118568 458872
rect 117228 453620 117280 453626
rect 117228 453562 117280 453568
rect 114468 453484 114520 453490
rect 114468 453426 114520 453432
rect 118620 453422 118648 474943
rect 121196 474910 121224 475487
rect 121366 475008 121422 475017
rect 121366 474943 121422 474952
rect 121184 474904 121236 474910
rect 119986 474872 120042 474881
rect 121184 474846 121236 474852
rect 121274 474872 121330 474881
rect 119986 474807 120042 474816
rect 121274 474807 121330 474816
rect 118608 453416 118660 453422
rect 118608 453358 118660 453364
rect 120000 453354 120028 474807
rect 121288 468654 121316 474807
rect 121380 474774 121408 474943
rect 121368 474768 121420 474774
rect 121368 474710 121420 474716
rect 122668 470594 122696 477799
rect 165434 476232 165490 476241
rect 165434 476167 165490 476176
rect 129554 476096 129610 476105
rect 129554 476031 129610 476040
rect 132406 476096 132462 476105
rect 132406 476031 132462 476040
rect 133786 476096 133842 476105
rect 133786 476031 133842 476040
rect 143354 476096 143410 476105
rect 143354 476031 143410 476040
rect 148322 476096 148378 476105
rect 148322 476031 148378 476040
rect 124034 475824 124090 475833
rect 124034 475759 124090 475768
rect 122668 470566 122788 470594
rect 121276 468648 121328 468654
rect 121276 468590 121328 468596
rect 122760 453762 122788 470566
rect 124048 470014 124076 475759
rect 126886 475280 126942 475289
rect 126886 475215 126888 475224
rect 126940 475215 126942 475224
rect 126888 475186 126940 475192
rect 128266 475144 128322 475153
rect 128266 475079 128268 475088
rect 128320 475079 128322 475088
rect 128268 475050 128320 475056
rect 129568 474910 129596 476031
rect 129646 475416 129702 475425
rect 129646 475351 129702 475360
rect 129660 475318 129688 475351
rect 129648 475312 129700 475318
rect 129648 475254 129700 475260
rect 131026 475280 131082 475289
rect 131026 475215 131082 475224
rect 131040 475182 131068 475215
rect 131028 475176 131080 475182
rect 131028 475118 131080 475124
rect 129004 474904 129056 474910
rect 124126 474872 124182 474881
rect 124126 474807 124182 474816
rect 125506 474872 125562 474881
rect 125506 474807 125562 474816
rect 128266 474872 128322 474881
rect 129004 474846 129056 474852
rect 129556 474904 129608 474910
rect 129556 474846 129608 474852
rect 131026 474872 131082 474881
rect 128266 474807 128322 474816
rect 124036 470008 124088 470014
rect 124036 469950 124088 469956
rect 122748 453756 122800 453762
rect 122748 453698 122800 453704
rect 124140 453694 124168 474807
rect 125520 457570 125548 474807
rect 126244 474768 126296 474774
rect 126244 474710 126296 474716
rect 125508 457564 125560 457570
rect 125508 457506 125560 457512
rect 126256 453830 126284 474710
rect 128280 460290 128308 474807
rect 128268 460284 128320 460290
rect 128268 460226 128320 460232
rect 129016 453898 129044 474846
rect 131026 474807 131082 474816
rect 131040 471442 131068 474807
rect 131028 471436 131080 471442
rect 131028 471378 131080 471384
rect 129004 453892 129056 453898
rect 129004 453834 129056 453840
rect 126244 453824 126296 453830
rect 126244 453766 126296 453772
rect 124128 453688 124180 453694
rect 124128 453630 124180 453636
rect 132420 453558 132448 476031
rect 133694 475144 133750 475153
rect 133694 475079 133750 475088
rect 133708 472734 133736 475079
rect 133696 472728 133748 472734
rect 133696 472670 133748 472676
rect 132408 453552 132460 453558
rect 132408 453494 132460 453500
rect 119988 453348 120040 453354
rect 119988 453290 120040 453296
rect 133800 452062 133828 476031
rect 141790 475824 141846 475833
rect 141790 475759 141846 475768
rect 141804 475386 141832 475759
rect 141792 475380 141844 475386
rect 141792 475322 141844 475328
rect 139306 475280 139362 475289
rect 139306 475215 139362 475224
rect 136454 475008 136510 475017
rect 136454 474943 136510 474952
rect 135166 474872 135222 474881
rect 135166 474807 135222 474816
rect 136362 474872 136418 474881
rect 136362 474807 136418 474816
rect 135180 456754 135208 474807
rect 136376 474094 136404 474807
rect 136364 474088 136416 474094
rect 136364 474030 136416 474036
rect 136468 470594 136496 474943
rect 136546 474872 136602 474881
rect 136546 474807 136602 474816
rect 137926 474872 137982 474881
rect 137926 474807 137982 474816
rect 139214 474872 139270 474881
rect 139214 474807 139270 474816
rect 136560 474230 136588 474807
rect 136548 474224 136600 474230
rect 136548 474166 136600 474172
rect 137284 474224 137336 474230
rect 137284 474166 137336 474172
rect 136468 470566 136588 470594
rect 136560 464506 136588 470566
rect 136548 464500 136600 464506
rect 136548 464442 136600 464448
rect 135168 456748 135220 456754
rect 135168 456690 135220 456696
rect 137296 452130 137324 474166
rect 137940 456142 137968 474807
rect 137928 456136 137980 456142
rect 137928 456078 137980 456084
rect 139228 452198 139256 474807
rect 139320 474162 139348 475215
rect 140686 474872 140742 474881
rect 140686 474807 140742 474816
rect 139308 474156 139360 474162
rect 139308 474098 139360 474104
rect 140700 452606 140728 474807
rect 143368 472802 143396 476031
rect 143446 474872 143502 474881
rect 143446 474807 143502 474816
rect 143356 472796 143408 472802
rect 143356 472738 143408 472744
rect 143460 453966 143488 474807
rect 148336 454918 148364 476031
rect 151358 475552 151414 475561
rect 151358 475487 151414 475496
rect 151372 475454 151400 475487
rect 151360 475448 151412 475454
rect 151360 475390 151412 475396
rect 151728 475448 151780 475454
rect 151728 475390 151780 475396
rect 150346 474872 150402 474881
rect 150346 474807 150402 474816
rect 150360 454986 150388 474807
rect 150348 454980 150400 454986
rect 150348 454922 150400 454928
rect 148324 454912 148376 454918
rect 148324 454854 148376 454860
rect 143448 453960 143500 453966
rect 143448 453902 143500 453908
rect 140688 452600 140740 452606
rect 140688 452542 140740 452548
rect 151740 452266 151768 475390
rect 151728 452260 151780 452266
rect 151728 452202 151780 452208
rect 139216 452192 139268 452198
rect 139216 452134 139268 452140
rect 137284 452124 137336 452130
rect 137284 452066 137336 452072
rect 133788 452056 133840 452062
rect 133788 451998 133840 452004
rect 34520 451988 34572 451994
rect 34520 451930 34572 451936
rect 66168 451988 66220 451994
rect 66168 451930 66220 451936
rect 45652 451920 45704 451926
rect 45650 451888 45652 451897
rect 45704 451888 45706 451897
rect 45650 451823 45706 451832
rect 48042 451344 48098 451353
rect 48042 451279 48098 451288
rect 48056 451246 48084 451279
rect 29828 451240 29880 451246
rect 29828 451182 29880 451188
rect 48044 451240 48096 451246
rect 48044 451182 48096 451188
rect 29840 431954 29868 451182
rect 165448 449993 165476 476167
rect 165528 476128 165580 476134
rect 165528 476070 165580 476076
rect 165540 450702 165568 476070
rect 166724 475584 166776 475590
rect 166724 475526 166776 475532
rect 165528 450696 165580 450702
rect 165528 450638 165580 450644
rect 165434 449984 165490 449993
rect 165434 449919 165490 449928
rect 166736 449274 166764 475526
rect 166724 449268 166776 449274
rect 166724 449210 166776 449216
rect 29748 431926 29868 431954
rect 29644 363860 29696 363866
rect 29644 363802 29696 363808
rect 29656 362982 29684 363802
rect 29748 363662 29776 431926
rect 139216 364336 139268 364342
rect 42890 364304 42946 364313
rect 42890 364239 42946 364248
rect 112994 364304 113050 364313
rect 112994 364239 113050 364248
rect 115754 364304 115810 364313
rect 115754 364239 115810 364248
rect 132958 364304 133014 364313
rect 132958 364239 133014 364248
rect 136546 364304 136602 364313
rect 139216 364278 139268 364284
rect 143354 364304 143410 364313
rect 136546 364239 136602 364248
rect 42798 364168 42854 364177
rect 42798 364103 42854 364112
rect 42812 363866 42840 364103
rect 42800 363860 42852 363866
rect 42800 363802 42852 363808
rect 42904 363730 42932 364239
rect 63406 364168 63462 364177
rect 63406 364103 63462 364112
rect 66166 364168 66222 364177
rect 66166 364103 66222 364112
rect 73158 364168 73214 364177
rect 73158 364103 73214 364112
rect 75826 364168 75882 364177
rect 75826 364103 75882 364112
rect 84106 364168 84162 364177
rect 84106 364103 84162 364112
rect 85670 364168 85726 364177
rect 85670 364103 85726 364112
rect 93766 364168 93822 364177
rect 93766 364103 93822 364112
rect 95606 364168 95662 364177
rect 95606 364103 95662 364112
rect 103150 364168 103206 364177
rect 103150 364103 103206 364112
rect 106186 364168 106242 364177
rect 106186 364103 106242 364112
rect 109590 364168 109646 364177
rect 109590 364103 109646 364112
rect 42892 363724 42944 363730
rect 42892 363666 42944 363672
rect 29736 363656 29788 363662
rect 29736 363598 29788 363604
rect 46940 363656 46992 363662
rect 46940 363598 46992 363604
rect 29644 362976 29696 362982
rect 29644 362918 29696 362924
rect 46952 340950 46980 363598
rect 60646 363080 60702 363089
rect 60646 363015 60702 363024
rect 29828 340944 29880 340950
rect 29828 340886 29880 340892
rect 46940 340944 46992 340950
rect 46940 340886 46992 340892
rect 29552 340264 29604 340270
rect 29552 340206 29604 340212
rect 29564 335354 29592 340206
rect 29564 335326 29684 335354
rect 29460 253224 29512 253230
rect 29460 253166 29512 253172
rect 28816 247036 28868 247042
rect 28816 246978 28868 246984
rect 28724 242888 28776 242894
rect 28724 242830 28776 242836
rect 28908 235272 28960 235278
rect 28908 235214 28960 235220
rect 28724 229628 28776 229634
rect 28724 229570 28776 229576
rect 28632 138712 28684 138718
rect 28632 138654 28684 138660
rect 28540 117156 28592 117162
rect 28540 117098 28592 117104
rect 27434 49464 27490 49473
rect 27434 49399 27490 49408
rect 27342 47832 27398 47841
rect 27342 47767 27398 47776
rect 27250 46472 27306 46481
rect 27250 46407 27306 46416
rect 27158 43752 27214 43761
rect 27158 43687 27214 43696
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 28644 27606 28672 138654
rect 28736 117230 28764 229570
rect 28816 138848 28868 138854
rect 28816 138790 28868 138796
rect 28828 138582 28856 138790
rect 28816 138576 28868 138582
rect 28816 138518 28868 138524
rect 28724 117224 28776 117230
rect 28724 117166 28776 117172
rect 28632 27600 28684 27606
rect 28632 27542 28684 27548
rect 28828 27538 28856 138518
rect 28920 109313 28948 235214
rect 29656 229090 29684 335326
rect 29840 230450 29868 340886
rect 46952 340785 46980 340886
rect 46938 340776 46994 340785
rect 46938 340711 46994 340720
rect 46204 340264 46256 340270
rect 46202 340232 46204 340241
rect 46256 340232 46258 340241
rect 46202 340167 46258 340176
rect 35164 339584 35216 339590
rect 35162 339552 35164 339561
rect 35216 339552 35218 339561
rect 35162 339487 35218 339496
rect 60660 339454 60688 363015
rect 63420 358086 63448 364103
rect 63408 358080 63460 358086
rect 63408 358022 63460 358028
rect 66180 340270 66208 364103
rect 68926 363080 68982 363089
rect 68926 363015 68982 363024
rect 71686 363080 71742 363089
rect 71686 363015 71742 363024
rect 68940 340338 68968 363015
rect 68928 340332 68980 340338
rect 68928 340274 68980 340280
rect 66168 340264 66220 340270
rect 66168 340206 66220 340212
rect 60648 339448 60700 339454
rect 60648 339390 60700 339396
rect 71700 339046 71728 363015
rect 73172 360874 73200 364103
rect 73160 360868 73212 360874
rect 73160 360810 73212 360816
rect 75840 352578 75868 364103
rect 78586 363080 78642 363089
rect 78586 363015 78642 363024
rect 81346 363080 81402 363089
rect 81346 363015 81402 363024
rect 75828 352572 75880 352578
rect 75828 352514 75880 352520
rect 78600 348430 78628 363015
rect 78588 348424 78640 348430
rect 78588 348366 78640 348372
rect 71688 339040 71740 339046
rect 71688 338982 71740 338988
rect 81360 338978 81388 363015
rect 84120 345710 84148 364103
rect 85684 355366 85712 364103
rect 88246 363080 88302 363089
rect 88246 363015 88302 363024
rect 91006 363080 91062 363089
rect 91006 363015 91062 363024
rect 85672 355360 85724 355366
rect 85672 355302 85724 355308
rect 88260 354006 88288 363015
rect 88248 354000 88300 354006
rect 88248 353942 88300 353948
rect 84108 345704 84160 345710
rect 84108 345646 84160 345652
rect 91020 342922 91048 363015
rect 93780 349858 93808 364103
rect 95620 356726 95648 364103
rect 99286 363080 99342 363089
rect 99286 363015 99342 363024
rect 100666 363080 100722 363089
rect 100666 363015 100722 363024
rect 95608 356720 95660 356726
rect 95608 356662 95660 356668
rect 99300 351218 99328 363015
rect 99288 351212 99340 351218
rect 99288 351154 99340 351160
rect 93768 349852 93820 349858
rect 93768 349794 93820 349800
rect 100680 347070 100708 363015
rect 103164 359514 103192 364103
rect 103152 359508 103204 359514
rect 103152 359450 103204 359456
rect 100668 347064 100720 347070
rect 100668 347006 100720 347012
rect 106200 344350 106228 364103
rect 108854 363352 108910 363361
rect 108854 363287 108910 363296
rect 107566 363080 107622 363089
rect 107566 363015 107622 363024
rect 107580 353297 107608 363015
rect 108868 362234 108896 363287
rect 108946 363080 109002 363089
rect 108946 363015 109002 363024
rect 108856 362228 108908 362234
rect 108856 362170 108908 362176
rect 107566 353288 107622 353297
rect 107566 353223 107622 353232
rect 108960 347750 108988 363015
rect 109604 356046 109632 364103
rect 111614 363216 111670 363225
rect 111614 363151 111670 363160
rect 109592 356040 109644 356046
rect 109592 355982 109644 355988
rect 111628 352646 111656 363151
rect 111706 363080 111762 363089
rect 111706 363015 111762 363024
rect 111616 352640 111668 352646
rect 111616 352582 111668 352588
rect 108948 347744 109000 347750
rect 108948 347686 109000 347692
rect 106188 344344 106240 344350
rect 106188 344286 106240 344292
rect 111720 343641 111748 363015
rect 113008 350538 113036 364239
rect 113086 364168 113142 364177
rect 113086 364103 113142 364112
rect 114466 364168 114522 364177
rect 114466 364103 114522 364112
rect 112996 350532 113048 350538
rect 112996 350474 113048 350480
rect 113100 348498 113128 364103
rect 114374 363080 114430 363089
rect 114374 363015 114430 363024
rect 114388 358698 114416 363015
rect 114376 358692 114428 358698
rect 114376 358634 114428 358640
rect 113088 348492 113140 348498
rect 113088 348434 113140 348440
rect 111706 343632 111762 343641
rect 111706 343567 111762 343576
rect 91008 342916 91060 342922
rect 91008 342858 91060 342864
rect 114480 340882 114508 364103
rect 115768 354686 115796 364239
rect 115846 364168 115902 364177
rect 115846 364103 115902 364112
rect 124034 364168 124090 364177
rect 124034 364103 124090 364112
rect 125966 364168 126022 364177
rect 125966 364103 126022 364112
rect 129554 364168 129610 364177
rect 129554 364103 129610 364112
rect 132038 364168 132094 364177
rect 132038 364103 132094 364112
rect 115756 354680 115808 354686
rect 115756 354622 115808 354628
rect 115860 349926 115888 364103
rect 122746 363896 122802 363905
rect 122746 363831 122802 363840
rect 122760 363798 122788 363831
rect 122748 363792 122800 363798
rect 122748 363734 122800 363740
rect 119986 363352 120042 363361
rect 119986 363287 120042 363296
rect 118514 363216 118570 363225
rect 118514 363151 118570 363160
rect 117226 363080 117282 363089
rect 117226 363015 117282 363024
rect 115848 349920 115900 349926
rect 115848 349862 115900 349868
rect 117240 346322 117268 363015
rect 118528 351286 118556 363151
rect 118606 363080 118662 363089
rect 118606 363015 118662 363024
rect 118516 351280 118568 351286
rect 118516 351222 118568 351228
rect 118620 347138 118648 363015
rect 120000 356794 120028 363287
rect 121274 363216 121330 363225
rect 121274 363151 121330 363160
rect 121182 363080 121238 363089
rect 121182 363015 121238 363024
rect 119988 356788 120040 356794
rect 119988 356730 120040 356736
rect 118608 347132 118660 347138
rect 118608 347074 118660 347080
rect 117228 346316 117280 346322
rect 117228 346258 117280 346264
rect 114468 340876 114520 340882
rect 114468 340818 114520 340824
rect 121196 339386 121224 363015
rect 121288 344486 121316 363151
rect 121276 344480 121328 344486
rect 121276 344422 121328 344428
rect 122760 341562 122788 363734
rect 124048 351354 124076 364103
rect 125508 363928 125560 363934
rect 125508 363870 125560 363876
rect 124126 363488 124182 363497
rect 124126 363423 124182 363432
rect 124140 362370 124168 363423
rect 125520 363225 125548 363870
rect 125506 363216 125562 363225
rect 125506 363151 125562 363160
rect 125414 363080 125470 363089
rect 125414 363015 125470 363024
rect 124128 362364 124180 362370
rect 124128 362306 124180 362312
rect 125428 354074 125456 363015
rect 125416 354068 125468 354074
rect 125416 354010 125468 354016
rect 124036 351348 124088 351354
rect 124036 351290 124088 351296
rect 125520 344418 125548 363151
rect 125980 360126 126008 364103
rect 127622 364032 127678 364041
rect 127622 363967 127678 363976
rect 127636 361010 127664 363967
rect 128266 363760 128322 363769
rect 128266 363695 128322 363704
rect 128280 363662 128308 363695
rect 128268 363656 128320 363662
rect 128268 363598 128320 363604
rect 128174 363080 128230 363089
rect 128174 363015 128230 363024
rect 127624 361004 127676 361010
rect 127624 360946 127676 360952
rect 125968 360120 126020 360126
rect 125968 360062 126020 360068
rect 128188 355434 128216 363015
rect 128280 355502 128308 363598
rect 128268 355496 128320 355502
rect 128268 355438 128320 355444
rect 128176 355428 128228 355434
rect 128176 355370 128228 355376
rect 129568 354142 129596 364103
rect 130936 363996 130988 364002
rect 130936 363938 130988 363944
rect 129648 363860 129700 363866
rect 129648 363802 129700 363808
rect 129660 363089 129688 363802
rect 130948 363225 130976 363938
rect 130934 363216 130990 363225
rect 130934 363151 130990 363160
rect 129646 363080 129702 363089
rect 129646 363015 129702 363024
rect 129556 354136 129608 354142
rect 129556 354078 129608 354084
rect 129660 347206 129688 363015
rect 130948 351422 130976 363151
rect 131026 363080 131082 363089
rect 131026 363015 131082 363024
rect 130936 351416 130988 351422
rect 130936 351358 130988 351364
rect 129648 347200 129700 347206
rect 129648 347142 129700 347148
rect 125508 344412 125560 344418
rect 125508 344354 125560 344360
rect 131040 342990 131068 363015
rect 132052 358154 132080 364103
rect 132040 358148 132092 358154
rect 132040 358090 132092 358096
rect 132972 356930 133000 364239
rect 133142 364168 133198 364177
rect 133142 364103 133198 364112
rect 135902 364168 135958 364177
rect 136560 364138 136588 364239
rect 135902 364103 135958 364112
rect 136548 364132 136600 364138
rect 133156 361078 133184 364103
rect 135166 363760 135222 363769
rect 135166 363695 135222 363704
rect 135180 363089 135208 363695
rect 135166 363080 135222 363089
rect 135166 363015 135222 363024
rect 133144 361072 133196 361078
rect 133144 361014 133196 361020
rect 132960 356924 133012 356930
rect 132960 356866 133012 356872
rect 131028 342984 131080 342990
rect 131028 342926 131080 342932
rect 122748 341556 122800 341562
rect 122748 341498 122800 341504
rect 135180 340406 135208 363015
rect 135916 359582 135944 364103
rect 136548 364074 136600 364080
rect 136560 364018 136588 364074
rect 136468 363990 136588 364018
rect 135904 359576 135956 359582
rect 135904 359518 135956 359524
rect 136468 356862 136496 363990
rect 136546 363896 136602 363905
rect 136546 363831 136602 363840
rect 136560 363390 136588 363831
rect 138294 363488 138350 363497
rect 138294 363423 138350 363432
rect 136548 363384 136600 363390
rect 136548 363326 136600 363332
rect 137928 363316 137980 363322
rect 137928 363258 137980 363264
rect 137940 363089 137968 363258
rect 137926 363080 137982 363089
rect 137926 363015 137982 363024
rect 136456 356856 136508 356862
rect 136456 356798 136508 356804
rect 137940 349994 137968 363015
rect 138308 362438 138336 363423
rect 139228 363089 139256 364278
rect 143354 364239 143410 364248
rect 139214 363080 139270 363089
rect 139214 363015 139270 363024
rect 140318 363080 140374 363089
rect 140318 363015 140374 363024
rect 142066 363080 142122 363089
rect 142066 363015 142122 363024
rect 138296 362432 138348 362438
rect 138296 362374 138348 362380
rect 137928 349988 137980 349994
rect 137928 349930 137980 349936
rect 139228 345778 139256 363015
rect 140332 360194 140360 363015
rect 140320 360188 140372 360194
rect 140320 360130 140372 360136
rect 139216 345772 139268 345778
rect 139216 345714 139268 345720
rect 142080 342242 142108 363015
rect 143368 360942 143396 364239
rect 143446 364168 143502 364177
rect 143446 364103 143502 364112
rect 150346 364168 150402 364177
rect 150402 364126 150480 364154
rect 150346 364103 150402 364112
rect 143356 360936 143408 360942
rect 143356 360878 143408 360884
rect 143460 345030 143488 364103
rect 148968 363520 149020 363526
rect 148968 363462 149020 363468
rect 146944 363384 146996 363390
rect 146944 363326 146996 363332
rect 146956 362302 146984 363326
rect 148980 363089 149008 363462
rect 148966 363080 149022 363089
rect 148966 363015 149022 363024
rect 146944 362296 146996 362302
rect 146944 362238 146996 362244
rect 148980 348566 149008 363015
rect 150452 361146 150480 364126
rect 151174 363624 151230 363633
rect 151174 363559 151230 363568
rect 151188 362982 151216 363559
rect 151176 362976 151228 362982
rect 151176 362918 151228 362924
rect 150440 361140 150492 361146
rect 150440 361082 150492 361088
rect 167012 360942 167040 587250
rect 168104 587240 168156 587246
rect 168104 587182 168156 587188
rect 168012 587172 168064 587178
rect 168012 587114 168064 587120
rect 167828 587104 167880 587110
rect 167828 587046 167880 587052
rect 167092 586560 167144 586566
rect 167092 586502 167144 586508
rect 167104 475454 167132 586502
rect 167184 585064 167236 585070
rect 167184 585006 167236 585012
rect 167196 476134 167224 585006
rect 167644 584316 167696 584322
rect 167644 584258 167696 584264
rect 167184 476128 167236 476134
rect 167184 476070 167236 476076
rect 167092 475448 167144 475454
rect 167092 475390 167144 475396
rect 167552 474836 167604 474842
rect 167552 474778 167604 474784
rect 167276 452600 167328 452606
rect 167276 452542 167328 452548
rect 167288 451926 167316 452542
rect 167276 451920 167328 451926
rect 167274 451888 167276 451897
rect 167328 451888 167330 451897
rect 167274 451823 167330 451832
rect 167288 451797 167316 451823
rect 167564 379506 167592 474778
rect 167656 382226 167684 584258
rect 167736 567928 167788 567934
rect 167736 567870 167788 567876
rect 167748 385014 167776 567870
rect 167840 440230 167868 587046
rect 167920 586900 167972 586906
rect 167920 586842 167972 586848
rect 167932 441590 167960 586842
rect 168024 450906 168052 587114
rect 168012 450900 168064 450906
rect 168012 450842 168064 450848
rect 168116 450770 168144 587182
rect 168196 563848 168248 563854
rect 168196 563790 168248 563796
rect 168208 450838 168236 563790
rect 168378 514992 168434 515001
rect 168378 514927 168434 514936
rect 168288 457564 168340 457570
rect 168288 457506 168340 457512
rect 168196 450832 168248 450838
rect 168196 450774 168248 450780
rect 168104 450764 168156 450770
rect 168104 450706 168156 450712
rect 167920 441584 167972 441590
rect 167920 441526 167972 441532
rect 167828 440224 167880 440230
rect 167828 440166 167880 440172
rect 167736 385008 167788 385014
rect 167736 384950 167788 384956
rect 167734 382392 167790 382401
rect 167734 382327 167790 382336
rect 167644 382220 167696 382226
rect 167644 382162 167696 382168
rect 167552 379500 167604 379506
rect 167552 379442 167604 379448
rect 167184 364200 167236 364206
rect 167182 364168 167184 364177
rect 167236 364168 167238 364177
rect 167182 364103 167238 364112
rect 167748 363594 167776 382327
rect 167736 363588 167788 363594
rect 167736 363530 167788 363536
rect 167840 363322 167868 440166
rect 167828 363316 167880 363322
rect 167828 363258 167880 363264
rect 167092 362976 167144 362982
rect 167092 362918 167144 362924
rect 167000 360936 167052 360942
rect 167000 360878 167052 360884
rect 167104 360618 167132 362918
rect 167932 361554 167960 441526
rect 168012 438932 168064 438938
rect 168012 438874 168064 438880
rect 168024 362302 168052 438874
rect 168194 423600 168250 423609
rect 168194 423535 168250 423544
rect 168104 422340 168156 422346
rect 168104 422282 168156 422288
rect 168116 364342 168144 422282
rect 168104 364336 168156 364342
rect 168104 364278 168156 364284
rect 168208 364138 168236 423535
rect 168196 364132 168248 364138
rect 168196 364074 168248 364080
rect 168012 362296 168064 362302
rect 168012 362238 168064 362244
rect 167920 361548 167972 361554
rect 167920 361490 167972 361496
rect 167184 361140 167236 361146
rect 167184 361082 167236 361088
rect 167012 360590 167132 360618
rect 166264 358080 166316 358086
rect 166264 358022 166316 358028
rect 148968 348560 149020 348566
rect 148968 348502 149020 348508
rect 143448 345024 143500 345030
rect 143448 344966 143500 344972
rect 142068 342236 142120 342242
rect 142068 342178 142120 342184
rect 135168 340400 135220 340406
rect 135168 340342 135220 340348
rect 121184 339380 121236 339386
rect 121184 339322 121236 339328
rect 81348 338972 81400 338978
rect 81348 338914 81400 338920
rect 166276 338094 166304 358022
rect 166264 338088 166316 338094
rect 166264 338030 166316 338036
rect 166724 254584 166776 254590
rect 166724 254526 166776 254532
rect 128084 253836 128136 253842
rect 128084 253778 128136 253784
rect 115664 253768 115716 253774
rect 60646 253736 60702 253745
rect 60646 253671 60702 253680
rect 65706 253736 65762 253745
rect 65706 253671 65762 253680
rect 70674 253736 70730 253745
rect 70674 253671 70730 253680
rect 75550 253736 75606 253745
rect 75550 253671 75606 253680
rect 98274 253736 98330 253745
rect 98274 253671 98330 253680
rect 115662 253736 115664 253745
rect 128096 253745 128124 253778
rect 115716 253736 115718 253745
rect 115662 253671 115718 253680
rect 118330 253736 118386 253745
rect 118330 253671 118386 253680
rect 123022 253736 123078 253745
rect 123022 253671 123078 253680
rect 125506 253736 125562 253745
rect 125506 253671 125508 253680
rect 43350 253600 43406 253609
rect 43350 253535 43406 253544
rect 43364 253230 43392 253535
rect 60660 253230 60688 253671
rect 65720 253298 65748 253671
rect 70688 253366 70716 253671
rect 75564 253434 75592 253671
rect 98288 253502 98316 253671
rect 118344 253570 118372 253671
rect 123036 253638 123064 253671
rect 125560 253671 125562 253680
rect 128082 253736 128138 253745
rect 128082 253671 128138 253680
rect 125508 253642 125560 253648
rect 123024 253632 123076 253638
rect 123024 253574 123076 253580
rect 130566 253600 130622 253609
rect 118332 253564 118384 253570
rect 130566 253535 130622 253544
rect 136454 253600 136510 253609
rect 136454 253535 136510 253544
rect 118332 253506 118384 253512
rect 98276 253496 98328 253502
rect 98276 253438 98328 253444
rect 75552 253428 75604 253434
rect 75552 253370 75604 253376
rect 70676 253360 70728 253366
rect 70676 253302 70728 253308
rect 65708 253292 65760 253298
rect 65708 253234 65760 253240
rect 43352 253224 43404 253230
rect 43352 253166 43404 253172
rect 60648 253224 60700 253230
rect 60648 253166 60700 253172
rect 34520 252544 34572 252550
rect 34520 252486 34572 252492
rect 29828 230444 29880 230450
rect 29828 230386 29880 230392
rect 29840 229634 29868 230386
rect 29828 229628 29880 229634
rect 29828 229570 29880 229576
rect 29644 229084 29696 229090
rect 29644 229026 29696 229032
rect 34532 227798 34560 252486
rect 43364 251433 43392 253166
rect 130580 253162 130608 253535
rect 132958 253464 133014 253473
rect 132958 253399 133014 253408
rect 130568 253156 130620 253162
rect 130568 253098 130620 253104
rect 132972 253094 133000 253399
rect 132960 253088 133012 253094
rect 132960 253030 133012 253036
rect 63406 252512 63462 252521
rect 63406 252447 63462 252456
rect 68190 252512 68246 252521
rect 68190 252447 68246 252456
rect 73158 252512 73214 252521
rect 73158 252447 73214 252456
rect 78126 252512 78182 252521
rect 78126 252447 78182 252456
rect 81254 252512 81310 252521
rect 81254 252447 81310 252456
rect 83554 252512 83610 252521
rect 83554 252447 83610 252456
rect 85670 252512 85726 252521
rect 85670 252447 85726 252456
rect 88246 252512 88302 252521
rect 88246 252447 88302 252456
rect 90822 252512 90878 252521
rect 90822 252447 90878 252456
rect 93214 252512 93270 252521
rect 93214 252447 93270 252456
rect 95606 252512 95662 252521
rect 95606 252447 95662 252456
rect 100574 252512 100630 252521
rect 100574 252447 100630 252456
rect 103150 252512 103206 252521
rect 103150 252447 103206 252456
rect 106094 252512 106150 252521
rect 106094 252447 106150 252456
rect 108486 252512 108542 252521
rect 108486 252447 108542 252456
rect 110510 252512 110566 252521
rect 110510 252447 110566 252456
rect 113086 252512 113142 252521
rect 113086 252447 113142 252456
rect 115846 252512 115902 252521
rect 115846 252447 115902 252456
rect 120906 252512 120962 252521
rect 120906 252447 120962 252456
rect 135994 252512 136050 252521
rect 135994 252447 136050 252456
rect 63420 251598 63448 252447
rect 68204 252414 68232 252447
rect 68192 252408 68244 252414
rect 68192 252350 68244 252356
rect 73172 252278 73200 252447
rect 78140 252346 78168 252447
rect 78128 252340 78180 252346
rect 78128 252282 78180 252288
rect 73160 252272 73212 252278
rect 73160 252214 73212 252220
rect 63408 251592 63460 251598
rect 63408 251534 63460 251540
rect 43350 251424 43406 251433
rect 43350 251359 43406 251368
rect 81268 251190 81296 252447
rect 83568 252210 83596 252447
rect 83556 252204 83608 252210
rect 83556 252146 83608 252152
rect 85684 252074 85712 252447
rect 85672 252068 85724 252074
rect 85672 252010 85724 252016
rect 81256 251184 81308 251190
rect 81256 251126 81308 251132
rect 88260 251122 88288 252447
rect 90836 252006 90864 252447
rect 90824 252000 90876 252006
rect 90824 251942 90876 251948
rect 93228 251938 93256 252447
rect 95620 252142 95648 252447
rect 95608 252136 95660 252142
rect 95608 252078 95660 252084
rect 93216 251932 93268 251938
rect 93216 251874 93268 251880
rect 100588 251870 100616 252447
rect 100576 251864 100628 251870
rect 100576 251806 100628 251812
rect 88248 251116 88300 251122
rect 88248 251058 88300 251064
rect 103164 251054 103192 252447
rect 103152 251048 103204 251054
rect 103152 250990 103204 250996
rect 106108 250986 106136 252447
rect 107566 251288 107622 251297
rect 107566 251223 107622 251232
rect 106096 250980 106148 250986
rect 106096 250922 106148 250928
rect 50342 250472 50398 250481
rect 50342 250407 50398 250416
rect 47584 238060 47636 238066
rect 47584 238002 47636 238008
rect 47596 230450 47624 238002
rect 47584 230444 47636 230450
rect 47584 230386 47636 230392
rect 46756 229084 46808 229090
rect 46756 229026 46808 229032
rect 29828 227792 29880 227798
rect 29828 227734 29880 227740
rect 34520 227792 34572 227798
rect 35164 227792 35216 227798
rect 34520 227734 34572 227740
rect 35162 227760 35164 227769
rect 46768 227769 46796 229026
rect 47596 227769 47624 230386
rect 50356 229090 50384 250407
rect 107580 238746 107608 251223
rect 108500 250850 108528 252447
rect 110326 252376 110382 252385
rect 110326 252311 110382 252320
rect 108946 251288 109002 251297
rect 108946 251223 109002 251232
rect 108488 250844 108540 250850
rect 108488 250786 108540 250792
rect 107568 238740 107620 238746
rect 107568 238682 107620 238688
rect 108960 234598 108988 251223
rect 108948 234592 109000 234598
rect 108948 234534 109000 234540
rect 110340 233238 110368 252311
rect 110524 250782 110552 252447
rect 111706 252376 111762 252385
rect 111706 252311 111762 252320
rect 112994 252376 113050 252385
rect 112994 252311 113050 252320
rect 110512 250776 110564 250782
rect 110512 250718 110564 250724
rect 110328 233232 110380 233238
rect 110328 233174 110380 233180
rect 111720 231810 111748 252311
rect 113008 244186 113036 252311
rect 113100 250918 113128 252447
rect 114466 252376 114522 252385
rect 114466 252311 114522 252320
rect 114374 251968 114430 251977
rect 114374 251903 114430 251912
rect 113088 250912 113140 250918
rect 113088 250854 113140 250860
rect 114388 249694 114416 251903
rect 114376 249688 114428 249694
rect 114376 249630 114428 249636
rect 114480 248402 114508 252311
rect 114468 248396 114520 248402
rect 114468 248338 114520 248344
rect 112996 244180 113048 244186
rect 112996 244122 113048 244128
rect 115860 240106 115888 252447
rect 120920 251802 120948 252447
rect 126886 252376 126942 252385
rect 126886 252311 126942 252320
rect 129554 252376 129610 252385
rect 129554 252311 129610 252320
rect 132038 252376 132094 252385
rect 132038 252311 132094 252320
rect 133786 252376 133842 252385
rect 133786 252311 133842 252320
rect 120908 251796 120960 251802
rect 120908 251738 120960 251744
rect 121182 251696 121238 251705
rect 121182 251631 121238 251640
rect 117226 251288 117282 251297
rect 117226 251223 117282 251232
rect 118606 251288 118662 251297
rect 118606 251223 118662 251232
rect 119986 251288 120042 251297
rect 119986 251223 120042 251232
rect 115848 240100 115900 240106
rect 115848 240042 115900 240048
rect 117240 237386 117268 251223
rect 117228 237380 117280 237386
rect 117228 237322 117280 237328
rect 118620 235958 118648 251223
rect 120000 242826 120028 251223
rect 119988 242820 120040 242826
rect 119988 242762 120040 242768
rect 118608 235952 118660 235958
rect 118608 235894 118660 235900
rect 121196 234530 121224 251631
rect 121274 251288 121330 251297
rect 121274 251223 121330 251232
rect 122746 251288 122802 251297
rect 122746 251223 122802 251232
rect 124126 251288 124182 251297
rect 124126 251223 124182 251232
rect 125506 251288 125562 251297
rect 125506 251223 125562 251232
rect 121288 241398 121316 251223
rect 122760 245546 122788 251223
rect 124140 246974 124168 251223
rect 124128 246968 124180 246974
rect 124128 246910 124180 246916
rect 122748 245540 122800 245546
rect 122748 245482 122800 245488
rect 121276 241392 121328 241398
rect 121276 241334 121328 241340
rect 121184 234524 121236 234530
rect 121184 234466 121236 234472
rect 125520 233170 125548 251223
rect 126900 248266 126928 252311
rect 128266 251288 128322 251297
rect 128266 251223 128322 251232
rect 126888 248260 126940 248266
rect 126888 248202 126940 248208
rect 128280 238678 128308 251223
rect 129568 249762 129596 252311
rect 129646 251288 129702 251297
rect 129646 251223 129702 251232
rect 131026 251288 131082 251297
rect 131026 251223 131082 251232
rect 129556 249756 129608 249762
rect 129556 249698 129608 249704
rect 129660 240038 129688 251223
rect 129648 240032 129700 240038
rect 129648 239974 129700 239980
rect 128268 238672 128320 238678
rect 128268 238614 128320 238620
rect 131040 234462 131068 251223
rect 132052 248334 132080 252311
rect 132040 248328 132092 248334
rect 132040 248270 132092 248276
rect 131028 234456 131080 234462
rect 131028 234398 131080 234404
rect 125508 233164 125560 233170
rect 125508 233106 125560 233112
rect 111708 231804 111760 231810
rect 111708 231746 111760 231752
rect 50344 229084 50396 229090
rect 50344 229026 50396 229032
rect 35216 227760 35218 227769
rect 29840 140146 29868 227734
rect 35162 227695 35218 227704
rect 46754 227760 46810 227769
rect 46754 227695 46810 227704
rect 47582 227760 47638 227769
rect 133800 227730 133828 252311
rect 136008 251734 136036 252447
rect 135996 251728 136048 251734
rect 135996 251670 136048 251676
rect 136362 251696 136418 251705
rect 136362 251631 136418 251640
rect 135166 251288 135222 251297
rect 135166 251223 135222 251232
rect 135180 229090 135208 251223
rect 135168 229084 135220 229090
rect 135168 229026 135220 229032
rect 47582 227695 47638 227704
rect 133788 227724 133840 227730
rect 133788 227666 133840 227672
rect 136376 227594 136404 251631
rect 136468 229022 136496 253535
rect 143354 252512 143410 252521
rect 143354 252447 143410 252456
rect 148322 252512 148378 252521
rect 148322 252447 148378 252456
rect 151082 252512 151138 252521
rect 151082 252447 151138 252456
rect 138294 252376 138350 252385
rect 138294 252311 138350 252320
rect 137926 251288 137982 251297
rect 137926 251223 137982 251232
rect 136456 229016 136508 229022
rect 136456 228958 136508 228964
rect 137940 227662 137968 251223
rect 138308 250714 138336 252311
rect 142066 251968 142122 251977
rect 142066 251903 142122 251912
rect 139214 251288 139270 251297
rect 139214 251223 139270 251232
rect 140686 251288 140742 251297
rect 140686 251223 140742 251232
rect 138296 250708 138348 250714
rect 138296 250650 138348 250656
rect 139228 235890 139256 251223
rect 140700 246362 140728 251223
rect 140688 246356 140740 246362
rect 140688 246298 140740 246304
rect 142080 237318 142108 251903
rect 143368 249626 143396 252447
rect 143446 252376 143502 252385
rect 143446 252311 143502 252320
rect 143356 249620 143408 249626
rect 143356 249562 143408 249568
rect 143460 244118 143488 252311
rect 143448 244112 143500 244118
rect 143448 244054 143500 244060
rect 142068 237312 142120 237318
rect 142068 237254 142120 237260
rect 139216 235884 139268 235890
rect 139216 235826 139268 235832
rect 148336 231130 148364 252447
rect 151096 251666 151124 252447
rect 166736 251802 166764 254526
rect 167012 252770 167040 360590
rect 167196 354674 167224 361082
rect 167932 361078 167960 361490
rect 167920 361072 167972 361078
rect 167920 361014 167972 361020
rect 167644 359508 167696 359514
rect 167644 359450 167696 359456
rect 166920 252742 167040 252770
rect 167104 354646 167224 354674
rect 166920 252362 166948 252742
rect 166998 252648 167054 252657
rect 166998 252583 167054 252592
rect 167012 252482 167040 252583
rect 167000 252476 167052 252482
rect 167000 252418 167052 252424
rect 166920 252334 167040 252362
rect 167012 251802 167040 252334
rect 167104 252113 167132 354646
rect 167656 318782 167684 359450
rect 167828 356720 167880 356726
rect 167828 356662 167880 356668
rect 167736 352640 167788 352646
rect 167736 352582 167788 352588
rect 167644 318776 167696 318782
rect 167644 318718 167696 318724
rect 167748 314634 167776 352582
rect 167840 322930 167868 356662
rect 168300 347682 168328 457506
rect 168392 402937 168420 514927
rect 168470 511864 168526 511873
rect 168470 511799 168526 511808
rect 168378 402928 168434 402937
rect 168378 402863 168434 402872
rect 168392 401713 168420 402863
rect 168378 401704 168434 401713
rect 168378 401639 168434 401648
rect 168484 399809 168512 511799
rect 168576 506161 168604 618151
rect 168930 599992 168986 600001
rect 168930 599927 168986 599936
rect 168746 598088 168802 598097
rect 168746 598023 168802 598032
rect 168654 512000 168710 512009
rect 168654 511935 168710 511944
rect 168668 510785 168696 511935
rect 168654 510776 168710 510785
rect 168654 510711 168710 510720
rect 168562 506152 168618 506161
rect 168562 506087 168618 506096
rect 168562 456240 168618 456249
rect 168562 456175 168618 456184
rect 168576 455569 168604 456175
rect 168562 455560 168618 455569
rect 168562 455495 168618 455504
rect 168470 399800 168526 399809
rect 168470 399735 168526 399744
rect 168668 398857 168696 510711
rect 168760 499574 168788 598023
rect 168760 499546 168880 499574
rect 168852 486470 168880 499546
rect 168944 487937 168972 599927
rect 169036 539646 169064 626855
rect 169114 625968 169170 625977
rect 169114 625903 169170 625912
rect 169128 539714 169156 625903
rect 169206 623792 169262 623801
rect 169206 623727 169262 623736
rect 169220 539782 169248 623727
rect 169298 622840 169354 622849
rect 169298 622775 169354 622784
rect 169312 539850 169340 622775
rect 169482 621072 169538 621081
rect 169482 621007 169538 621016
rect 169390 619984 169446 619993
rect 169390 619919 169446 619928
rect 169300 539844 169352 539850
rect 169300 539786 169352 539792
rect 169208 539776 169260 539782
rect 169208 539718 169260 539724
rect 169116 539708 169168 539714
rect 169116 539650 169168 539656
rect 169024 539640 169076 539646
rect 169024 539582 169076 539588
rect 169036 515001 169064 539582
rect 169022 514992 169078 515001
rect 169022 514927 169078 514936
rect 169128 513913 169156 539650
rect 169114 513904 169170 513913
rect 169114 513839 169170 513848
rect 169220 511873 169248 539718
rect 169312 512009 169340 539786
rect 169298 512000 169354 512009
rect 169298 511935 169354 511944
rect 169206 511864 169262 511873
rect 169206 511799 169262 511808
rect 169404 509234 169432 619919
rect 169036 509206 169432 509234
rect 169036 507929 169064 509206
rect 169496 509017 169524 621007
rect 169666 598360 169722 598369
rect 169666 598295 169722 598304
rect 169574 513904 169630 513913
rect 169574 513839 169630 513848
rect 169482 509008 169538 509017
rect 169482 508943 169538 508952
rect 169022 507920 169078 507929
rect 169022 507855 169078 507864
rect 168930 487928 168986 487937
rect 168930 487863 168986 487872
rect 168944 487257 168972 487863
rect 168930 487248 168986 487257
rect 168930 487183 168986 487192
rect 168840 486464 168892 486470
rect 168840 486406 168892 486412
rect 168852 486169 168880 486406
rect 168838 486160 168894 486169
rect 168838 486095 168894 486104
rect 168748 456748 168800 456754
rect 168748 456690 168800 456696
rect 168760 455841 168788 456690
rect 168746 455832 168802 455841
rect 168746 455767 168802 455776
rect 168760 455462 168788 455767
rect 168748 455456 168800 455462
rect 168748 455398 168800 455404
rect 169036 449886 169064 507855
rect 169114 506152 169170 506161
rect 169114 506087 169170 506096
rect 169024 449880 169076 449886
rect 169024 449822 169076 449828
rect 168838 448624 168894 448633
rect 168838 448559 168894 448568
rect 168746 399800 168802 399809
rect 168746 399735 168802 399744
rect 168654 398848 168710 398857
rect 168654 398783 168710 398792
rect 168654 397080 168710 397089
rect 168654 397015 168710 397024
rect 168378 375320 168434 375329
rect 168378 375255 168434 375264
rect 168392 374377 168420 375255
rect 168378 374368 168434 374377
rect 168378 374303 168434 374312
rect 168288 347676 168340 347682
rect 168288 347618 168340 347624
rect 167920 344344 167972 344350
rect 167920 344286 167972 344292
rect 167828 322924 167880 322930
rect 167828 322866 167880 322872
rect 167932 317422 167960 344286
rect 168012 339040 168064 339046
rect 168012 338982 168064 338988
rect 168024 335306 168052 338982
rect 168012 335300 168064 335306
rect 168012 335242 168064 335248
rect 167920 317416 167972 317422
rect 167920 317358 167972 317364
rect 167736 314628 167788 314634
rect 167736 314570 167788 314576
rect 167644 296744 167696 296750
rect 167644 296686 167696 296692
rect 167656 253298 167684 296686
rect 167736 291236 167788 291242
rect 167736 291178 167788 291184
rect 167748 253434 167776 291178
rect 167920 287088 167972 287094
rect 167920 287030 167972 287036
rect 167828 280220 167880 280226
rect 167828 280162 167880 280168
rect 167840 253502 167868 280162
rect 167828 253496 167880 253502
rect 167828 253438 167880 253444
rect 167736 253428 167788 253434
rect 167736 253370 167788 253376
rect 167644 253292 167696 253298
rect 167644 253234 167696 253240
rect 167090 252104 167146 252113
rect 167932 252074 167960 287030
rect 168012 284368 168064 284374
rect 168012 284310 168064 284316
rect 167090 252039 167146 252048
rect 167920 252068 167972 252074
rect 166724 251796 166776 251802
rect 166724 251738 166776 251744
rect 167000 251796 167052 251802
rect 167000 251738 167052 251744
rect 167012 251666 167040 251738
rect 151084 251660 151136 251666
rect 151084 251602 151136 251608
rect 167000 251660 167052 251666
rect 167000 251602 167052 251608
rect 148324 231124 148376 231130
rect 148324 231066 148376 231072
rect 137928 227656 137980 227662
rect 137928 227598 137980 227604
rect 136364 227588 136416 227594
rect 136364 227530 136416 227536
rect 167104 142154 167132 252039
rect 167920 252010 167972 252016
rect 168024 252006 168052 284310
rect 168104 282940 168156 282946
rect 168104 282882 168156 282888
rect 168012 252000 168064 252006
rect 168012 251942 168064 251948
rect 168116 251938 168144 282882
rect 168196 278792 168248 278798
rect 168196 278734 168248 278740
rect 168104 251932 168156 251938
rect 168104 251874 168156 251880
rect 168208 251870 168236 278734
rect 168392 262313 168420 374303
rect 168562 374096 168618 374105
rect 168562 374031 168618 374040
rect 168378 262304 168434 262313
rect 168288 262268 168340 262274
rect 168378 262239 168434 262248
rect 168288 262210 168340 262216
rect 168196 251864 168248 251870
rect 168196 251806 168248 251812
rect 167828 251796 167880 251802
rect 167828 251738 167880 251744
rect 167644 246356 167696 246362
rect 167644 246298 167696 246304
rect 167656 245721 167684 246298
rect 167642 245712 167698 245721
rect 167642 245647 167698 245656
rect 167656 155242 167684 245647
rect 167736 155304 167788 155310
rect 167736 155246 167788 155252
rect 167644 155236 167696 155242
rect 167644 155178 167696 155184
rect 167012 142126 167132 142154
rect 122746 141808 122802 141817
rect 122746 141743 122802 141752
rect 133142 141808 133198 141817
rect 133142 141743 133198 141752
rect 108486 141672 108542 141681
rect 108486 141607 108542 141616
rect 112166 141672 112222 141681
rect 112166 141607 112222 141616
rect 108500 140826 108528 141607
rect 112180 140894 112208 141607
rect 112168 140888 112220 140894
rect 112168 140830 112220 140836
rect 108488 140820 108540 140826
rect 108488 140762 108540 140768
rect 109590 140720 109646 140729
rect 109590 140655 109646 140664
rect 113270 140720 113326 140729
rect 113270 140655 113326 140664
rect 116766 140720 116822 140729
rect 116766 140655 116822 140664
rect 118974 140720 119030 140729
rect 118974 140655 119030 140664
rect 43074 140176 43130 140185
rect 29828 140140 29880 140146
rect 29828 140082 29880 140088
rect 35900 140140 35952 140146
rect 43074 140111 43130 140120
rect 63222 140176 63278 140185
rect 63222 140111 63278 140120
rect 65798 140176 65854 140185
rect 65798 140111 65854 140120
rect 35900 140082 35952 140088
rect 35912 117298 35940 140082
rect 43088 138718 43116 140111
rect 43442 139360 43498 139369
rect 43442 139295 43498 139304
rect 60646 139360 60702 139369
rect 60646 139295 60702 139304
rect 43456 138854 43484 139295
rect 43444 138848 43496 138854
rect 43444 138790 43496 138796
rect 43076 138712 43128 138718
rect 43076 138654 43128 138660
rect 60660 138038 60688 139295
rect 60648 138032 60700 138038
rect 60648 137974 60700 137980
rect 63236 137902 63264 140111
rect 63224 137896 63276 137902
rect 63224 137838 63276 137844
rect 65812 136610 65840 140111
rect 109604 140078 109632 140655
rect 113284 140146 113312 140655
rect 116780 140214 116808 140655
rect 118988 140282 119016 140655
rect 118976 140276 119028 140282
rect 118976 140218 119028 140224
rect 116768 140208 116820 140214
rect 115478 140176 115534 140185
rect 113272 140140 113324 140146
rect 115478 140111 115534 140120
rect 115846 140176 115902 140185
rect 116768 140150 116820 140156
rect 115846 140111 115902 140120
rect 113272 140082 113324 140088
rect 109592 140072 109644 140078
rect 109592 140014 109644 140020
rect 107382 139360 107438 139369
rect 107382 139295 107438 139304
rect 110878 139360 110934 139369
rect 110878 139295 110934 139304
rect 114374 139360 114430 139369
rect 114374 139295 114430 139304
rect 107396 139126 107424 139295
rect 107384 139120 107436 139126
rect 107384 139062 107436 139068
rect 110892 138990 110920 139295
rect 114388 139058 114416 139295
rect 115492 139194 115520 140111
rect 115480 139188 115532 139194
rect 115480 139130 115532 139136
rect 114376 139052 114428 139058
rect 114376 138994 114428 139000
rect 110880 138984 110932 138990
rect 110880 138926 110932 138932
rect 68926 138680 68982 138689
rect 68926 138615 68982 138624
rect 65800 136604 65852 136610
rect 65800 136546 65852 136552
rect 68940 135250 68968 138615
rect 71042 138136 71098 138145
rect 71042 138071 71098 138080
rect 74446 138136 74502 138145
rect 74446 138071 74502 138080
rect 75826 138136 75882 138145
rect 75826 138071 75882 138080
rect 78586 138136 78642 138145
rect 78586 138071 78642 138080
rect 81346 138136 81402 138145
rect 81346 138071 81402 138080
rect 84106 138136 84162 138145
rect 84106 138071 84162 138080
rect 86866 138136 86922 138145
rect 86866 138071 86922 138080
rect 88246 138136 88302 138145
rect 88246 138071 88302 138080
rect 91006 138136 91062 138145
rect 91006 138071 91062 138080
rect 93766 138136 93822 138145
rect 93766 138071 93822 138080
rect 96526 138136 96582 138145
rect 96526 138071 96582 138080
rect 99286 138136 99342 138145
rect 99286 138071 99342 138080
rect 100666 138136 100722 138145
rect 100666 138071 100722 138080
rect 103426 138136 103482 138145
rect 103426 138071 103482 138080
rect 106186 138136 106242 138145
rect 106186 138071 106242 138080
rect 108946 138136 109002 138145
rect 108946 138071 109002 138080
rect 111706 138136 111762 138145
rect 111706 138071 111762 138080
rect 113086 138136 113142 138145
rect 113086 138071 113142 138080
rect 68928 135244 68980 135250
rect 68928 135186 68980 135192
rect 71056 133890 71084 138071
rect 71044 133884 71096 133890
rect 71044 133826 71096 133832
rect 74460 132462 74488 138071
rect 74448 132456 74500 132462
rect 74448 132398 74500 132404
rect 75840 132394 75868 138071
rect 75828 132388 75880 132394
rect 75828 132330 75880 132336
rect 78600 131102 78628 138071
rect 78588 131096 78640 131102
rect 78588 131038 78640 131044
rect 81360 129742 81388 138071
rect 81348 129736 81400 129742
rect 81348 129678 81400 129684
rect 84120 128314 84148 138071
rect 84108 128308 84160 128314
rect 84108 128250 84160 128256
rect 86880 126954 86908 138071
rect 86868 126948 86920 126954
rect 86868 126890 86920 126896
rect 88260 125594 88288 138071
rect 88248 125588 88300 125594
rect 88248 125530 88300 125536
rect 91020 124166 91048 138071
rect 91008 124160 91060 124166
rect 91008 124102 91060 124108
rect 93780 122806 93808 138071
rect 93768 122800 93820 122806
rect 93768 122742 93820 122748
rect 96540 121446 96568 138071
rect 96528 121440 96580 121446
rect 96528 121382 96580 121388
rect 99300 120086 99328 138071
rect 99288 120080 99340 120086
rect 99288 120022 99340 120028
rect 100680 120018 100708 138071
rect 100668 120012 100720 120018
rect 100668 119954 100720 119960
rect 103440 118658 103468 138071
rect 103428 118652 103480 118658
rect 103428 118594 103480 118600
rect 35900 117292 35952 117298
rect 35900 117234 35952 117240
rect 35806 117192 35862 117201
rect 35912 117178 35940 117234
rect 106200 117230 106228 138071
rect 35862 117150 35940 117178
rect 46940 117224 46992 117230
rect 46940 117166 46992 117172
rect 106188 117224 106240 117230
rect 106188 117166 106240 117172
rect 45836 117156 45888 117162
rect 35806 117127 35862 117136
rect 45836 117098 45888 117104
rect 45848 117065 45876 117098
rect 45834 117056 45890 117065
rect 45834 116991 45890 117000
rect 46952 116793 46980 117166
rect 46938 116784 46994 116793
rect 46938 116719 46994 116728
rect 108960 115938 108988 138071
rect 108948 115932 109000 115938
rect 108948 115874 109000 115880
rect 111720 114510 111748 138071
rect 113100 123486 113128 138071
rect 115860 126274 115888 140111
rect 120356 139392 120408 139398
rect 117870 139360 117926 139369
rect 117870 139295 117926 139304
rect 120354 139360 120356 139369
rect 120408 139360 120410 139369
rect 120354 139295 120410 139304
rect 121366 139360 121422 139369
rect 121366 139295 121422 139304
rect 122654 139360 122710 139369
rect 122654 139295 122710 139304
rect 117884 138786 117912 139295
rect 121380 139262 121408 139295
rect 121368 139256 121420 139262
rect 121368 139198 121420 139204
rect 122668 138922 122696 139295
rect 122656 138916 122708 138922
rect 122656 138858 122708 138864
rect 117872 138780 117924 138786
rect 117872 138722 117924 138728
rect 122760 138689 122788 141743
rect 123758 141672 123814 141681
rect 123758 141607 123814 141616
rect 128542 141672 128598 141681
rect 128542 141607 128598 141616
rect 123772 141030 123800 141607
rect 128556 141234 128584 141607
rect 133156 141370 133184 141743
rect 134246 141672 134302 141681
rect 134246 141607 134302 141616
rect 136546 141672 136602 141681
rect 136546 141607 136602 141616
rect 140042 141672 140098 141681
rect 140042 141607 140098 141616
rect 142342 141672 142398 141681
rect 142342 141607 142398 141616
rect 133144 141364 133196 141370
rect 133144 141306 133196 141312
rect 128544 141228 128596 141234
rect 128544 141170 128596 141176
rect 134260 141098 134288 141607
rect 134248 141092 134300 141098
rect 134248 141034 134300 141040
rect 123760 141024 123812 141030
rect 123760 140966 123812 140972
rect 136560 140962 136588 141607
rect 140056 141302 140084 141607
rect 140044 141296 140096 141302
rect 140044 141238 140096 141244
rect 142356 141166 142384 141607
rect 166172 141500 166224 141506
rect 166172 141442 166224 141448
rect 142344 141160 142396 141166
rect 142344 141102 142396 141108
rect 136548 140956 136600 140962
rect 136548 140898 136600 140904
rect 137928 140752 137980 140758
rect 125966 140720 126022 140729
rect 125966 140655 126022 140664
rect 132038 140720 132094 140729
rect 132038 140655 132094 140664
rect 135350 140720 135406 140729
rect 135350 140655 135352 140664
rect 125980 140350 126008 140655
rect 132052 140418 132080 140655
rect 135404 140655 135406 140664
rect 137926 140720 137928 140729
rect 137980 140720 137982 140729
rect 137926 140655 137982 140664
rect 139030 140720 139086 140729
rect 139030 140655 139086 140664
rect 141238 140720 141294 140729
rect 141238 140655 141294 140664
rect 143446 140720 143502 140729
rect 143446 140655 143502 140664
rect 149518 140720 149574 140729
rect 149518 140655 149574 140664
rect 135352 140626 135404 140632
rect 139044 140554 139072 140655
rect 141252 140622 141280 140655
rect 141240 140616 141292 140622
rect 141240 140558 141292 140564
rect 139032 140548 139084 140554
rect 139032 140490 139084 140496
rect 143460 140486 143488 140655
rect 143448 140480 143500 140486
rect 143448 140422 143500 140428
rect 132040 140412 132092 140418
rect 132040 140354 132092 140360
rect 125968 140344 126020 140350
rect 125968 140286 126020 140292
rect 129646 140176 129702 140185
rect 129646 140111 129702 140120
rect 125230 139360 125286 139369
rect 125230 139295 125286 139304
rect 127714 139360 127770 139369
rect 129660 139330 129688 140111
rect 149532 139466 149560 140655
rect 149520 139460 149572 139466
rect 149520 139402 149572 139408
rect 130750 139360 130806 139369
rect 127714 139295 127770 139304
rect 129648 139324 129700 139330
rect 122746 138680 122802 138689
rect 122746 138615 122802 138624
rect 124126 138680 124182 138689
rect 125244 138650 125272 139295
rect 127728 138718 127756 139295
rect 130750 139295 130806 139304
rect 148414 139360 148470 139369
rect 148414 139295 148470 139304
rect 151082 139360 151138 139369
rect 151082 139295 151138 139304
rect 129648 139266 129700 139272
rect 130764 138854 130792 139295
rect 136454 139088 136510 139097
rect 136454 139023 136510 139032
rect 130752 138848 130804 138854
rect 130752 138790 130804 138796
rect 127716 138712 127768 138718
rect 127716 138654 127768 138660
rect 124126 138615 124182 138624
rect 125232 138644 125284 138650
rect 118422 138136 118478 138145
rect 118422 138071 118478 138080
rect 121366 138136 121422 138145
rect 121366 138071 121422 138080
rect 117228 138032 117280 138038
rect 117228 137974 117280 137980
rect 117240 137834 117268 137974
rect 117228 137828 117280 137834
rect 117228 137770 117280 137776
rect 118436 133210 118464 138071
rect 118424 133204 118476 133210
rect 118424 133146 118476 133152
rect 121380 130422 121408 138071
rect 124140 134570 124168 138615
rect 125232 138586 125284 138592
rect 125414 138136 125470 138145
rect 125414 138071 125470 138080
rect 128266 138136 128322 138145
rect 128266 138071 128322 138080
rect 131026 138136 131082 138145
rect 131026 138071 131082 138080
rect 133786 138136 133842 138145
rect 133786 138071 133842 138080
rect 124128 134564 124180 134570
rect 124128 134506 124180 134512
rect 121368 130416 121420 130422
rect 121368 130358 121420 130364
rect 125428 129062 125456 138071
rect 125416 129056 125468 129062
rect 125416 128998 125468 129004
rect 128280 127634 128308 138071
rect 128268 127628 128320 127634
rect 128268 127570 128320 127576
rect 115848 126268 115900 126274
rect 115848 126210 115900 126216
rect 131040 124914 131068 138071
rect 133800 126342 133828 138071
rect 136468 135930 136496 139023
rect 148428 138582 148456 139295
rect 148416 138576 148468 138582
rect 148416 138518 148468 138524
rect 151096 138514 151124 139295
rect 166184 138582 166212 141442
rect 166264 141432 166316 141438
rect 166264 141374 166316 141380
rect 166276 139126 166304 141374
rect 167012 139942 167040 142126
rect 167000 139936 167052 139942
rect 167000 139878 167052 139884
rect 167012 139466 167040 139878
rect 167000 139460 167052 139466
rect 167000 139402 167052 139408
rect 166264 139120 166316 139126
rect 166264 139062 166316 139068
rect 166172 138576 166224 138582
rect 166172 138518 166224 138524
rect 151084 138508 151136 138514
rect 151084 138450 151136 138456
rect 139306 138136 139362 138145
rect 139306 138071 139362 138080
rect 136456 135924 136508 135930
rect 136456 135866 136508 135872
rect 133788 126336 133840 126342
rect 133788 126278 133840 126284
rect 131028 124908 131080 124914
rect 131028 124850 131080 124856
rect 139320 123554 139348 138071
rect 164884 136876 164936 136882
rect 164884 136818 164936 136824
rect 139308 123548 139360 123554
rect 139308 123490 139360 123496
rect 113088 123480 113140 123486
rect 113088 123422 113140 123428
rect 164896 117298 164924 136818
rect 164884 117292 164936 117298
rect 164884 117234 164936 117240
rect 111708 114504 111760 114510
rect 111708 114446 111760 114452
rect 28906 109304 28962 109313
rect 28906 109239 28962 109248
rect 143172 29912 143224 29918
rect 128358 29880 128414 29889
rect 143172 29854 143224 29860
rect 128358 29815 128414 29824
rect 135812 29844 135864 29850
rect 128372 29782 128400 29815
rect 135812 29786 135864 29792
rect 128360 29776 128412 29782
rect 128360 29718 128412 29724
rect 127624 29708 127676 29714
rect 127624 29650 127676 29656
rect 124036 29640 124088 29646
rect 75550 29608 75606 29617
rect 75550 29543 75606 29552
rect 88062 29608 88118 29617
rect 88062 29543 88118 29552
rect 90730 29608 90786 29617
rect 90730 29543 90786 29552
rect 122746 29608 122802 29617
rect 124036 29582 124088 29588
rect 122746 29543 122802 29552
rect 60646 28928 60702 28937
rect 60646 28863 60702 28872
rect 68190 28928 68246 28937
rect 68190 28863 68246 28872
rect 60660 28354 60688 28863
rect 60648 28348 60700 28354
rect 60648 28290 60700 28296
rect 68204 28286 68232 28863
rect 75564 28422 75592 29543
rect 78126 28928 78182 28937
rect 78126 28863 78182 28872
rect 80702 28928 80758 28937
rect 80702 28863 80758 28872
rect 83094 28928 83150 28937
rect 83094 28863 83150 28872
rect 78140 28490 78168 28863
rect 80716 28558 80744 28863
rect 83108 28626 83136 28863
rect 88076 28694 88104 29543
rect 90744 28762 90772 29543
rect 103150 28928 103206 28937
rect 103150 28863 103206 28872
rect 103164 28830 103192 28863
rect 103152 28824 103204 28830
rect 103152 28766 103204 28772
rect 90732 28756 90784 28762
rect 90732 28698 90784 28704
rect 88064 28688 88116 28694
rect 88064 28630 88116 28636
rect 83096 28620 83148 28626
rect 83096 28562 83148 28568
rect 80704 28552 80756 28558
rect 80704 28494 80756 28500
rect 78128 28484 78180 28490
rect 78128 28426 78180 28432
rect 75552 28416 75604 28422
rect 75552 28358 75604 28364
rect 68192 28280 68244 28286
rect 63222 28248 63278 28257
rect 68192 28222 68244 28228
rect 112166 28248 112222 28257
rect 63222 28183 63278 28192
rect 112166 28183 112222 28192
rect 115662 28248 115718 28257
rect 115662 28183 115718 28192
rect 42800 27600 42852 27606
rect 42798 27568 42800 27577
rect 42852 27568 42854 27577
rect 28816 27532 28868 27538
rect 42798 27503 42854 27512
rect 43626 27568 43682 27577
rect 43626 27503 43628 27512
rect 28816 27474 28868 27480
rect 43680 27503 43682 27512
rect 43628 27474 43680 27480
rect 63236 26722 63264 28183
rect 64878 27568 64934 27577
rect 64878 27503 64934 27512
rect 71594 27568 71650 27577
rect 71594 27503 71650 27512
rect 73986 27568 74042 27577
rect 73986 27503 74042 27512
rect 86590 27568 86646 27577
rect 86590 27503 86646 27512
rect 92754 27568 92810 27577
rect 92754 27503 92810 27512
rect 95238 27568 95294 27577
rect 95238 27503 95294 27512
rect 98274 27568 98330 27577
rect 98274 27503 98330 27512
rect 100206 27568 100262 27577
rect 100206 27503 100262 27512
rect 105542 27568 105598 27577
rect 105542 27503 105598 27512
rect 106278 27568 106334 27577
rect 106278 27503 106334 27512
rect 108026 27568 108082 27577
rect 108026 27503 108082 27512
rect 108762 27568 108818 27577
rect 108762 27503 108818 27512
rect 110326 27568 110382 27577
rect 110326 27503 110382 27512
rect 110970 27568 111026 27577
rect 110970 27503 111026 27512
rect 64892 26858 64920 27503
rect 64880 26852 64932 26858
rect 64880 26794 64932 26800
rect 63224 26716 63276 26722
rect 63224 26658 63276 26664
rect 71608 26654 71636 27503
rect 71596 26648 71648 26654
rect 71596 26590 71648 26596
rect 60740 25628 60792 25634
rect 60740 25570 60792 25576
rect 46940 24200 46992 24206
rect 46940 24142 46992 24148
rect 10324 24132 10376 24138
rect 10324 24074 10376 24080
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2792 16574 2820 22714
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 21626
rect 2792 16546 2912 16574
rect 4172 16546 5304 16574
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 4762
rect 2884 480 2912 16546
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 4080 480 4108 7550
rect 5276 480 5304 16546
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 354 6040 11766
rect 7668 480 7696 15846
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 480 8800 3470
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 11834
rect 10336 3534 10364 24074
rect 37280 22840 37332 22846
rect 37280 22782 37332 22788
rect 34520 21480 34572 21486
rect 34520 21422 34572 21428
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16592 16574 16620 21354
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22112 16574 22140 19926
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23492 16574 23520 18906
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 16592 16546 17080 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 12348 4888 12400 4894
rect 12348 4830 12400 4836
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11164 480 11192 3470
rect 12360 480 12388 4830
rect 13556 480 13584 8910
rect 14740 7676 14792 7682
rect 14740 7618 14792 7624
rect 14752 480 14780 7618
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15948 480 15976 4082
rect 17052 480 17080 16546
rect 18604 11960 18656 11966
rect 18604 11902 18656 11908
rect 17960 10328 18012 10334
rect 17960 10270 18012 10276
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 10270
rect 18616 4146 18644 11902
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19444 480 19472 3538
rect 20640 480 20668 3606
rect 21836 480 21864 6122
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25320 14476 25372 14482
rect 25320 14418 25372 14424
rect 25332 480 25360 14418
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 18566
rect 33140 17264 33192 17270
rect 33140 17206 33192 17212
rect 33152 16574 33180 17206
rect 33152 16546 33640 16574
rect 31944 12028 31996 12034
rect 31944 11970 31996 11976
rect 31300 9104 31352 9110
rect 31300 9046 31352 9052
rect 27712 9036 27764 9042
rect 27712 8978 27764 8984
rect 27724 480 27752 8978
rect 30104 6248 30156 6254
rect 30104 6190 30156 6196
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 28920 480 28948 3674
rect 30116 480 30144 6190
rect 31312 480 31340 9046
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 11970
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 21422
rect 37292 16574 37320 22782
rect 38660 20188 38712 20194
rect 38660 20130 38712 20136
rect 38672 16574 38700 20130
rect 44180 18692 44232 18698
rect 44180 18634 44232 18640
rect 44192 16574 44220 18634
rect 46952 16574 46980 24142
rect 53840 22908 53892 22914
rect 53840 22850 53892 22856
rect 51080 20120 51132 20126
rect 51080 20062 51132 20068
rect 48320 20052 48372 20058
rect 48320 19994 48372 20000
rect 48332 16574 48360 19994
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 44192 16546 45048 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 36728 10396 36780 10402
rect 36728 10338 36780 10344
rect 35992 3800 36044 3806
rect 35992 3742 36044 3748
rect 36004 480 36032 3742
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 10338
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 40224 15972 40276 15978
rect 40224 15914 40276 15920
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 15914
rect 41880 12096 41932 12102
rect 41880 12038 41932 12044
rect 41892 480 41920 12038
rect 44272 6316 44324 6322
rect 44272 6258 44324 6264
rect 43076 3868 43128 3874
rect 43076 3810 43128 3816
rect 43088 480 43116 3810
rect 44284 480 44312 6258
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46664 14544 46716 14550
rect 46664 14486 46716 14492
rect 46676 480 46704 14486
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50160 12164 50212 12170
rect 50160 12106 50212 12112
rect 50172 480 50200 12106
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 20062
rect 53852 16574 53880 22850
rect 57980 21548 58032 21554
rect 57980 21490 58032 21496
rect 57992 16574 58020 21490
rect 53852 16546 54984 16574
rect 57992 16546 58480 16574
rect 52552 9172 52604 9178
rect 52552 9114 52604 9120
rect 52564 480 52592 9114
rect 53748 4956 53800 4962
rect 53748 4898 53800 4904
rect 53760 480 53788 4898
rect 54956 480 54984 16546
rect 56784 12232 56836 12238
rect 56784 12174 56836 12180
rect 56048 9240 56100 9246
rect 56048 9182 56100 9188
rect 56060 480 56088 9182
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 12174
rect 58452 480 58480 16546
rect 59636 9308 59688 9314
rect 59636 9250 59688 9256
rect 59648 480 59676 9250
rect 60752 6914 60780 25570
rect 60832 25560 60884 25566
rect 60832 25502 60884 25508
rect 60844 16574 60872 25502
rect 74000 24002 74028 27503
rect 86604 24750 86632 27503
rect 86592 24744 86644 24750
rect 86592 24686 86644 24692
rect 92768 24682 92796 27503
rect 92756 24676 92808 24682
rect 92756 24618 92808 24624
rect 89720 24336 89772 24342
rect 89720 24278 89772 24284
rect 85580 24268 85632 24274
rect 85580 24210 85632 24216
rect 73988 23996 74040 24002
rect 73988 23938 74040 23944
rect 69020 22976 69072 22982
rect 69020 22918 69072 22924
rect 62120 21616 62172 21622
rect 62120 21558 62172 21564
rect 62132 16574 62160 21558
rect 67640 17400 67692 17406
rect 67640 17342 67692 17348
rect 60844 16546 61608 16574
rect 62132 16546 63264 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64328 10464 64380 10470
rect 64328 10406 64380 10412
rect 64340 480 64368 10406
rect 66720 9376 66772 9382
rect 66720 9318 66772 9324
rect 65524 5024 65576 5030
rect 65524 4966 65576 4972
rect 65536 480 65564 4966
rect 66732 480 66760 9318
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 17342
rect 69032 3398 69060 22918
rect 84200 18828 84252 18834
rect 84200 18770 84252 18776
rect 69112 18760 69164 18766
rect 69112 18702 69164 18708
rect 69020 3392 69072 3398
rect 69020 3334 69072 3340
rect 69124 480 69152 18702
rect 81624 13592 81676 13598
rect 81624 13534 81676 13540
rect 80888 13184 80940 13190
rect 80888 13126 80940 13132
rect 77392 13116 77444 13122
rect 77392 13058 77444 13064
rect 75000 10736 75052 10742
rect 75000 10678 75052 10684
rect 72608 7744 72660 7750
rect 72608 7686 72660 7692
rect 71504 6384 71556 6390
rect 71504 6326 71556 6332
rect 69940 3392 69992 3398
rect 69940 3334 69992 3340
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3334
rect 71516 480 71544 6326
rect 72620 480 72648 7686
rect 73804 5092 73856 5098
rect 73804 5034 73856 5040
rect 73816 480 73844 5034
rect 75012 480 75040 10678
rect 76196 6520 76248 6526
rect 76196 6462 76248 6468
rect 76208 480 76236 6462
rect 77404 480 77432 13058
rect 78588 9444 78640 9450
rect 78588 9386 78640 9392
rect 78600 480 78628 9386
rect 79692 6452 79744 6458
rect 79692 6394 79744 6400
rect 79704 480 79732 6394
rect 80900 480 80928 13126
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 13534
rect 83280 6588 83332 6594
rect 83280 6530 83332 6536
rect 83292 480 83320 6530
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 18770
rect 85592 16574 85620 24210
rect 88340 23384 88392 23390
rect 88340 23326 88392 23332
rect 88352 16574 88380 23326
rect 89732 16574 89760 24278
rect 95252 23934 95280 27503
rect 98288 26246 98316 27503
rect 98276 26240 98328 26246
rect 98276 26182 98328 26188
rect 100220 26178 100248 27503
rect 100208 26172 100260 26178
rect 100208 26114 100260 26120
rect 105556 26110 105584 27503
rect 105544 26104 105596 26110
rect 105544 26046 105596 26052
rect 104900 25696 104952 25702
rect 104900 25638 104952 25644
rect 95240 23928 95292 23934
rect 95240 23870 95292 23876
rect 96620 20256 96672 20262
rect 96620 20198 96672 20204
rect 93860 17332 93912 17338
rect 93860 17274 93912 17280
rect 93872 16574 93900 17274
rect 96632 16574 96660 20198
rect 104912 16574 104940 25638
rect 106292 23458 106320 27503
rect 108040 25362 108068 27503
rect 108028 25356 108080 25362
rect 108028 25298 108080 25304
rect 106280 23452 106332 23458
rect 106280 23394 106332 23400
rect 107660 23044 107712 23050
rect 107660 22986 107712 22992
rect 107672 16574 107700 22986
rect 108776 22098 108804 27503
rect 110340 26926 110368 27503
rect 110328 26920 110380 26926
rect 110328 26862 110380 26868
rect 110984 22642 111012 27503
rect 111522 27432 111578 27441
rect 111522 27367 111578 27376
rect 111536 25498 111564 27367
rect 112180 26994 112208 28183
rect 112902 27568 112958 27577
rect 112902 27503 112958 27512
rect 112168 26988 112220 26994
rect 112168 26930 112220 26936
rect 111524 25492 111576 25498
rect 111524 25434 111576 25440
rect 112916 25430 112944 27503
rect 115676 27402 115704 28183
rect 122760 27713 122788 29543
rect 122746 27704 122802 27713
rect 122746 27639 122802 27648
rect 120632 27600 120684 27606
rect 117134 27568 117190 27577
rect 117134 27503 117190 27512
rect 118238 27568 118294 27577
rect 118238 27503 118294 27512
rect 118422 27568 118478 27577
rect 120632 27542 120684 27548
rect 120814 27568 120870 27577
rect 118422 27503 118478 27512
rect 115664 27396 115716 27402
rect 115664 27338 115716 27344
rect 114560 25764 114612 25770
rect 114560 25706 114612 25712
rect 112904 25424 112956 25430
rect 112904 25366 112956 25372
rect 111800 24404 111852 24410
rect 111800 24346 111852 24352
rect 110972 22636 111024 22642
rect 110972 22578 111024 22584
rect 108764 22092 108816 22098
rect 108764 22034 108816 22040
rect 111812 16574 111840 24346
rect 114572 16574 114600 25706
rect 117148 21350 117176 27503
rect 118252 22710 118280 27503
rect 118436 27470 118464 27503
rect 118424 27464 118476 27470
rect 118424 27406 118476 27412
rect 120078 27432 120134 27441
rect 120078 27367 120134 27376
rect 118240 22704 118292 22710
rect 118240 22646 118292 22652
rect 120092 22030 120120 27367
rect 120644 27305 120672 27542
rect 120814 27503 120870 27512
rect 120630 27296 120686 27305
rect 120630 27231 120686 27240
rect 120828 22574 120856 27503
rect 124048 27402 124076 29582
rect 127636 27606 127664 29650
rect 130566 29608 130622 29617
rect 130566 29543 130622 29552
rect 130580 29102 130608 29543
rect 130568 29096 130620 29102
rect 130568 29038 130620 29044
rect 134248 28960 134300 28966
rect 128542 28928 128598 28937
rect 128542 28863 128598 28872
rect 134246 28928 134248 28937
rect 134300 28928 134302 28937
rect 134246 28863 134302 28872
rect 128556 28218 128584 28863
rect 129646 28248 129702 28257
rect 128544 28212 128596 28218
rect 129646 28183 129702 28192
rect 132038 28248 132094 28257
rect 132038 28183 132094 28192
rect 128544 28154 128596 28160
rect 127624 27600 127676 27606
rect 124126 27568 124182 27577
rect 124126 27503 124182 27512
rect 126334 27568 126390 27577
rect 127624 27542 127676 27548
rect 128174 27568 128230 27577
rect 126334 27503 126390 27512
rect 128174 27503 128230 27512
rect 124036 27396 124088 27402
rect 124036 27338 124088 27344
rect 124140 27334 124168 27503
rect 124128 27328 124180 27334
rect 124128 27270 124180 27276
rect 126348 27198 126376 27503
rect 126336 27192 126388 27198
rect 123758 27160 123814 27169
rect 126336 27134 126388 27140
rect 123758 27095 123760 27104
rect 123812 27095 123814 27104
rect 123760 27066 123812 27072
rect 128188 27062 128216 27503
rect 129660 27266 129688 28183
rect 132052 27470 132080 28183
rect 132776 27600 132828 27606
rect 132774 27568 132776 27577
rect 132828 27568 132830 27577
rect 132774 27503 132830 27512
rect 135350 27568 135406 27577
rect 135350 27503 135406 27512
rect 132040 27464 132092 27470
rect 132040 27406 132092 27412
rect 129648 27260 129700 27266
rect 129648 27202 129700 27208
rect 128176 27056 128228 27062
rect 128176 26998 128228 27004
rect 128360 25832 128412 25838
rect 128360 25774 128412 25780
rect 120816 22568 120868 22574
rect 120816 22510 120868 22516
rect 120080 22024 120132 22030
rect 120080 21966 120132 21972
rect 126980 21752 127032 21758
rect 126980 21694 127032 21700
rect 117136 21344 117188 21350
rect 117136 21286 117188 21292
rect 118700 17808 118752 17814
rect 118700 17750 118752 17756
rect 85592 16546 85712 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 93872 16546 93992 16574
rect 96632 16546 97488 16574
rect 104912 16546 105768 16574
rect 107672 16546 108160 16574
rect 111812 16546 112392 16574
rect 114572 16546 114784 16574
rect 85684 480 85712 16546
rect 86408 16040 86460 16046
rect 86408 15982 86460 15988
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 15982
rect 87512 13252 87564 13258
rect 87512 13194 87564 13200
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 13194
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 92480 14612 92532 14618
rect 92480 14554 92532 14560
rect 91560 13320 91612 13326
rect 91560 13262 91612 13268
rect 91572 480 91600 13262
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 14554
rect 93964 480 93992 16546
rect 94688 13388 94740 13394
rect 94688 13330 94740 13336
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 13330
rect 95792 10804 95844 10810
rect 95792 10746 95844 10752
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 10746
rect 97460 480 97488 16546
rect 102140 16176 102192 16182
rect 102140 16118 102192 16124
rect 99840 14680 99892 14686
rect 99840 14622 99892 14628
rect 98644 6656 98696 6662
rect 98644 6598 98696 6604
rect 98656 480 98684 6598
rect 99852 480 99880 14622
rect 101036 5160 101088 5166
rect 101036 5102 101088 5108
rect 101048 480 101076 5102
rect 102152 3398 102180 16118
rect 102232 13456 102284 13462
rect 102232 13398 102284 13404
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 102244 480 102272 13398
rect 104072 10532 104124 10538
rect 104072 10474 104124 10480
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103348 480 103376 3334
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 10474
rect 105740 480 105768 16546
rect 106464 14748 106516 14754
rect 106464 14690 106516 14696
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 14690
rect 108132 480 108160 16546
rect 110512 14816 110564 14822
rect 110512 14758 110564 14764
rect 109040 13524 109092 13530
rect 109040 13466 109092 13472
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 13466
rect 110524 480 110552 14758
rect 111616 10600 111668 10606
rect 111616 10542 111668 10548
rect 111628 480 111656 10542
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 113824 11756 113876 11762
rect 113824 11698 113876 11704
rect 113836 3466 113864 11698
rect 114008 3936 114060 3942
rect 114008 3878 114060 3884
rect 113824 3460 113876 3466
rect 113824 3402 113876 3408
rect 114020 480 114048 3878
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116400 16108 116452 16114
rect 116400 16050 116452 16056
rect 116412 480 116440 16050
rect 117320 14884 117372 14890
rect 117320 14826 117372 14832
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 14826
rect 118712 3466 118740 17750
rect 125600 16244 125652 16250
rect 125600 16186 125652 16192
rect 120632 14952 120684 14958
rect 120632 14894 120684 14900
rect 118792 5228 118844 5234
rect 118792 5170 118844 5176
rect 118700 3460 118752 3466
rect 118700 3402 118752 3408
rect 118804 480 118832 5170
rect 119896 3460 119948 3466
rect 119896 3402 119948 3408
rect 119908 480 119936 3402
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 14894
rect 123484 7880 123536 7886
rect 123484 7822 123536 7828
rect 122288 7812 122340 7818
rect 122288 7754 122340 7760
rect 122300 480 122328 7754
rect 123496 480 123524 7822
rect 124680 4004 124732 4010
rect 124680 3946 124732 3952
rect 124692 480 124720 3946
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 16186
rect 126992 480 127020 21694
rect 127072 18896 127124 18902
rect 127072 18838 127124 18844
rect 127084 16574 127112 18838
rect 128372 16574 128400 25774
rect 135364 24070 135392 27503
rect 135824 26858 135852 29786
rect 138938 29608 138994 29617
rect 138938 29543 138994 29552
rect 138952 29034 138980 29543
rect 138940 29028 138992 29034
rect 138940 28970 138992 28976
rect 135902 28928 135958 28937
rect 135902 28863 135958 28872
rect 138294 28928 138350 28937
rect 138294 28863 138350 28872
rect 135916 28150 135944 28863
rect 135904 28144 135956 28150
rect 135904 28086 135956 28092
rect 138308 28082 138336 28863
rect 138296 28076 138348 28082
rect 138296 28018 138348 28024
rect 137190 27568 137246 27577
rect 137190 27503 137246 27512
rect 140134 27568 140190 27577
rect 140134 27503 140190 27512
rect 141238 27568 141294 27577
rect 141238 27503 141294 27512
rect 135812 26852 135864 26858
rect 135812 26794 135864 26800
rect 137204 24857 137232 27503
rect 140148 26858 140176 27503
rect 140136 26852 140188 26858
rect 140136 26794 140188 26800
rect 141252 26790 141280 27503
rect 141240 26784 141292 26790
rect 141240 26726 141292 26732
rect 143184 26654 143212 29854
rect 166172 29572 166224 29578
rect 166172 29514 166224 29520
rect 143264 28892 143316 28898
rect 143264 28834 143316 28840
rect 143276 27606 143304 28834
rect 149058 28384 149114 28393
rect 149058 28319 149114 28328
rect 143446 28248 143502 28257
rect 143446 28183 143502 28192
rect 143354 28112 143410 28121
rect 143354 28047 143410 28056
rect 143264 27600 143316 27606
rect 143264 27542 143316 27548
rect 143368 26926 143396 28047
rect 143460 27538 143488 28183
rect 147678 27568 147734 27577
rect 143448 27532 143500 27538
rect 147678 27503 147734 27512
rect 143448 27474 143500 27480
rect 143356 26920 143408 26926
rect 143356 26862 143408 26868
rect 143448 26920 143500 26926
rect 143448 26862 143500 26868
rect 143172 26648 143224 26654
rect 143460 26625 143488 26862
rect 143172 26590 143224 26596
rect 143446 26616 143502 26625
rect 143446 26551 143502 26560
rect 142160 26036 142212 26042
rect 142160 25978 142212 25984
rect 137190 24848 137246 24857
rect 137190 24783 137246 24792
rect 140780 24472 140832 24478
rect 140780 24414 140832 24420
rect 135352 24064 135404 24070
rect 135352 24006 135404 24012
rect 139400 23112 139452 23118
rect 139400 23054 139452 23060
rect 132500 21820 132552 21826
rect 132500 21762 132552 21768
rect 131120 17468 131172 17474
rect 131120 17410 131172 17416
rect 131132 16574 131160 17410
rect 132512 16574 132540 21762
rect 138020 20528 138072 20534
rect 138020 20470 138072 20476
rect 135260 19032 135312 19038
rect 135260 18974 135312 18980
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130568 7948 130620 7954
rect 130568 7890 130620 7896
rect 130580 480 130608 7890
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 134156 8016 134208 8022
rect 134156 7958 134208 7964
rect 134168 480 134196 7958
rect 135272 4078 135300 18974
rect 136640 17536 136692 17542
rect 136640 17478 136692 17484
rect 136652 16574 136680 17478
rect 138032 16574 138060 20470
rect 139412 16574 139440 23054
rect 140792 16574 140820 24414
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 135352 16312 135404 16318
rect 135352 16254 135404 16260
rect 135260 4072 135312 4078
rect 135260 4014 135312 4020
rect 135364 3482 135392 16254
rect 136456 4072 136508 4078
rect 136456 4014 136508 4020
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 4014
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 25978
rect 147692 24818 147720 27503
rect 149072 26994 149100 28319
rect 150624 27600 150676 27606
rect 150070 27568 150126 27577
rect 150070 27503 150126 27512
rect 150622 27568 150624 27577
rect 150676 27568 150678 27577
rect 150622 27503 150678 27512
rect 150084 26994 150112 27503
rect 166184 27062 166212 29514
rect 166264 29504 166316 29510
rect 166264 29446 166316 29452
rect 166276 27130 166304 29446
rect 166356 29436 166408 29442
rect 166356 29378 166408 29384
rect 166264 27124 166316 27130
rect 166264 27066 166316 27072
rect 166172 27056 166224 27062
rect 166172 26998 166224 27004
rect 149060 26988 149112 26994
rect 149060 26930 149112 26936
rect 150072 26988 150124 26994
rect 150072 26930 150124 26936
rect 166368 26722 166396 29378
rect 167012 26994 167040 139402
rect 167092 138508 167144 138514
rect 167092 138450 167144 138456
rect 167104 138310 167132 138450
rect 167092 138304 167144 138310
rect 167092 138246 167144 138252
rect 167104 27606 167132 138246
rect 167092 27600 167144 27606
rect 167092 27542 167144 27548
rect 167000 26988 167052 26994
rect 167000 26930 167052 26936
rect 167656 26858 167684 155178
rect 167644 26852 167696 26858
rect 167644 26794 167696 26800
rect 167748 26790 167776 155246
rect 167840 140010 167868 251738
rect 168300 251734 168328 262210
rect 168392 258074 168420 262239
rect 168576 262041 168604 374031
rect 168668 285025 168696 397015
rect 168760 288425 168788 399735
rect 168852 398342 168880 448559
rect 168930 401704 168986 401713
rect 168930 401639 168986 401648
rect 168840 398336 168892 398342
rect 168840 398278 168892 398284
rect 168838 395992 168894 396001
rect 168838 395927 168894 395936
rect 168746 288416 168802 288425
rect 168746 288351 168802 288360
rect 168746 285696 168802 285705
rect 168746 285631 168802 285640
rect 168654 285016 168710 285025
rect 168654 284951 168710 284960
rect 168562 262032 168618 262041
rect 168562 261967 168618 261976
rect 168576 261526 168604 261967
rect 168564 261520 168616 261526
rect 168564 261462 168616 261468
rect 168392 258046 168512 258074
rect 168288 251728 168340 251734
rect 168288 251670 168340 251676
rect 168196 238740 168248 238746
rect 168196 238682 168248 238688
rect 168208 238649 168236 238682
rect 168194 238640 168250 238649
rect 168194 238575 168250 238584
rect 168208 237454 168236 238575
rect 168196 237448 168248 237454
rect 168196 237390 168248 237396
rect 167920 211812 167972 211818
rect 167920 211754 167972 211760
rect 167828 140004 167880 140010
rect 167828 139946 167880 139952
rect 167840 138310 167868 139946
rect 167932 138650 167960 211754
rect 168104 204264 168156 204270
rect 168104 204206 168156 204212
rect 168012 203584 168064 203590
rect 168012 203526 168064 203532
rect 168024 140418 168052 203526
rect 168116 141370 168144 204206
rect 168196 200796 168248 200802
rect 168196 200738 168248 200744
rect 168104 141364 168156 141370
rect 168104 141306 168156 141312
rect 168208 140690 168236 200738
rect 168288 198008 168340 198014
rect 168288 197950 168340 197956
rect 168300 140758 168328 197950
rect 168484 171134 168512 258046
rect 168564 229084 168616 229090
rect 168564 229026 168616 229032
rect 168576 228993 168604 229026
rect 168562 228984 168618 228993
rect 168562 228919 168618 228928
rect 168576 227798 168604 228919
rect 168564 227792 168616 227798
rect 168564 227734 168616 227740
rect 168668 174706 168696 284951
rect 168760 174842 168788 285631
rect 168852 283937 168880 395927
rect 168944 290873 168972 401639
rect 169036 396001 169064 449822
rect 169128 449206 169156 506087
rect 169496 489914 169524 508943
rect 169312 489886 169524 489914
rect 169206 455560 169262 455569
rect 169206 455495 169262 455504
rect 169116 449200 169168 449206
rect 169116 449142 169168 449148
rect 169022 395992 169078 396001
rect 169022 395927 169078 395936
rect 169116 392012 169168 392018
rect 169116 391954 169168 391960
rect 168930 290864 168986 290873
rect 168930 290799 168986 290808
rect 168838 283928 168894 283937
rect 168838 283863 168894 283872
rect 168852 174978 168880 283863
rect 168944 178945 168972 290799
rect 169022 288416 169078 288425
rect 169022 288351 169078 288360
rect 169036 287745 169064 288351
rect 169022 287736 169078 287745
rect 169022 287671 169078 287680
rect 168930 178936 168986 178945
rect 168930 178871 168986 178880
rect 168944 178702 168972 178871
rect 168932 178696 168984 178702
rect 168932 178638 168984 178644
rect 169036 177562 169064 287671
rect 169128 282169 169156 391954
rect 169220 379545 169248 455495
rect 169312 451110 169340 489886
rect 169390 487248 169446 487257
rect 169390 487183 169446 487192
rect 169300 451104 169352 451110
rect 169300 451046 169352 451052
rect 169312 450226 169340 451046
rect 169300 450220 169352 450226
rect 169300 450162 169352 450168
rect 169404 448458 169432 487183
rect 169484 450220 169536 450226
rect 169484 450162 169536 450168
rect 169392 448452 169444 448458
rect 169392 448394 169444 448400
rect 169300 448384 169352 448390
rect 169300 448326 169352 448332
rect 169206 379536 169262 379545
rect 169206 379471 169262 379480
rect 169312 375329 169340 448326
rect 169404 376009 169432 448394
rect 169496 397089 169524 450162
rect 169588 401985 169616 513839
rect 169680 487150 169708 598295
rect 173162 587480 173218 587489
rect 170864 587444 170916 587450
rect 173162 587415 173218 587424
rect 170864 587386 170916 587392
rect 169760 586968 169812 586974
rect 169760 586910 169812 586916
rect 169668 487144 169720 487150
rect 169668 487086 169720 487092
rect 169680 486305 169708 487086
rect 169666 486296 169722 486305
rect 169666 486231 169722 486240
rect 169680 448390 169708 486231
rect 169668 448384 169720 448390
rect 169668 448326 169720 448332
rect 169772 440162 169800 586910
rect 170772 586696 170824 586702
rect 170772 586638 170824 586644
rect 169852 464500 169904 464506
rect 169852 464442 169904 464448
rect 169864 463758 169892 464442
rect 169852 463752 169904 463758
rect 169852 463694 169904 463700
rect 170404 463752 170456 463758
rect 170404 463694 170456 463700
rect 169852 455388 169904 455394
rect 169852 455330 169904 455336
rect 169864 454986 169892 455330
rect 169852 454980 169904 454986
rect 169852 454922 169904 454928
rect 169850 454744 169906 454753
rect 169850 454679 169906 454688
rect 169864 454073 169892 454679
rect 169850 454064 169906 454073
rect 169850 453999 169906 454008
rect 169852 453756 169904 453762
rect 169852 453698 169904 453704
rect 169864 452742 169892 453698
rect 169852 452736 169904 452742
rect 169852 452678 169904 452684
rect 169944 452260 169996 452266
rect 169944 452202 169996 452208
rect 169956 451314 169984 452202
rect 169944 451308 169996 451314
rect 169944 451250 169996 451256
rect 169760 440156 169812 440162
rect 169760 440098 169812 440104
rect 169772 438938 169800 440098
rect 169760 438932 169812 438938
rect 169760 438874 169812 438880
rect 169956 431954 169984 451250
rect 170312 451240 170364 451246
rect 170310 451208 170312 451217
rect 170364 451208 170366 451217
rect 170310 451143 170366 451152
rect 169864 431926 169984 431954
rect 169574 401976 169630 401985
rect 169574 401911 169630 401920
rect 169482 397080 169538 397089
rect 169482 397015 169538 397024
rect 169482 394224 169538 394233
rect 169482 394159 169538 394168
rect 169496 393310 169524 394159
rect 169484 393304 169536 393310
rect 169484 393246 169536 393252
rect 169496 392018 169524 393246
rect 169484 392012 169536 392018
rect 169484 391954 169536 391960
rect 169390 376000 169446 376009
rect 169390 375935 169446 375944
rect 169298 375320 169354 375329
rect 169298 375255 169354 375264
rect 169404 354674 169432 375935
rect 169220 354646 169432 354674
rect 169114 282160 169170 282169
rect 169114 282095 169170 282104
rect 168944 177534 169064 177562
rect 168944 176050 168972 177534
rect 168932 176044 168984 176050
rect 168932 175986 168984 175992
rect 168944 175817 168972 175986
rect 168930 175808 168986 175817
rect 168930 175743 168986 175752
rect 168852 174950 168972 174978
rect 168838 174856 168894 174865
rect 168760 174814 168838 174842
rect 168838 174791 168894 174800
rect 168668 174678 168788 174706
rect 168760 173194 168788 174678
rect 168852 174622 168880 174791
rect 168840 174616 168892 174622
rect 168840 174558 168892 174564
rect 168748 173188 168800 173194
rect 168748 173130 168800 173136
rect 168760 173097 168788 173130
rect 168746 173088 168802 173097
rect 168746 173023 168802 173032
rect 168944 172009 168972 174950
rect 168930 172000 168986 172009
rect 168930 171935 168986 171944
rect 168944 171834 168972 171935
rect 168932 171828 168984 171834
rect 168932 171770 168984 171776
rect 168484 171106 168604 171134
rect 168378 153096 168434 153105
rect 168378 153031 168434 153040
rect 168392 152017 168420 153031
rect 168378 152008 168434 152017
rect 168378 151943 168434 151952
rect 168288 140752 168340 140758
rect 168288 140694 168340 140700
rect 168196 140684 168248 140690
rect 168196 140626 168248 140632
rect 168012 140412 168064 140418
rect 168012 140354 168064 140360
rect 167920 138644 167972 138650
rect 167920 138586 167972 138592
rect 167828 138304 167880 138310
rect 167828 138246 167880 138252
rect 167828 126336 167880 126342
rect 167828 126278 167880 126284
rect 167840 103494 167868 126278
rect 167828 103488 167880 103494
rect 167828 103430 167880 103436
rect 167828 98048 167880 98054
rect 167828 97990 167880 97996
rect 167840 28354 167868 97990
rect 167920 92540 167972 92546
rect 167920 92482 167972 92488
rect 167828 28348 167880 28354
rect 167828 28290 167880 28296
rect 167736 26784 167788 26790
rect 167736 26726 167788 26732
rect 166356 26716 166408 26722
rect 166356 26658 166408 26664
rect 157340 25968 157392 25974
rect 157340 25910 157392 25916
rect 154580 25900 154632 25906
rect 154580 25842 154632 25848
rect 147680 24812 147732 24818
rect 147680 24754 147732 24760
rect 146300 24540 146352 24546
rect 146300 24482 146352 24488
rect 143540 17604 143592 17610
rect 143540 17546 143592 17552
rect 143552 480 143580 17546
rect 146312 16574 146340 24482
rect 149060 21956 149112 21962
rect 149060 21898 149112 21904
rect 147680 20324 147732 20330
rect 147680 20266 147732 20272
rect 147692 16574 147720 20266
rect 149072 16574 149100 21898
rect 150440 20392 150492 20398
rect 150440 20334 150492 20340
rect 150452 16574 150480 20334
rect 151820 19168 151872 19174
rect 151820 19110 151872 19116
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144736 16380 144788 16386
rect 144736 16322 144788 16328
rect 144748 480 144776 16322
rect 145932 8084 145984 8090
rect 145932 8026 145984 8032
rect 145944 480 145972 8026
rect 147140 480 147168 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 4078 151860 19110
rect 154592 16574 154620 25842
rect 157352 16574 157380 25910
rect 162860 24608 162912 24614
rect 162860 24550 162912 24556
rect 158720 21888 158772 21894
rect 158720 21830 158772 21836
rect 158732 16574 158760 21830
rect 161480 19100 161532 19106
rect 161480 19042 161532 19048
rect 160192 17740 160244 17746
rect 160192 17682 160244 17688
rect 160100 17672 160152 17678
rect 160100 17614 160152 17620
rect 154592 16546 155448 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153752 16448 153804 16454
rect 153752 16390 153804 16396
rect 151912 8152 151964 8158
rect 151912 8094 151964 8100
rect 151820 4072 151872 4078
rect 151820 4014 151872 4020
rect 151924 3482 151952 8094
rect 153016 4072 153068 4078
rect 153016 4014 153068 4020
rect 151832 3454 151952 3482
rect 151832 480 151860 3454
rect 153028 480 153056 4014
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16390
rect 155420 480 155448 16546
rect 156604 5296 156656 5302
rect 156604 5238 156656 5244
rect 156616 480 156644 5238
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11694 160140 17614
rect 160100 11688 160152 11694
rect 160100 11630 160152 11636
rect 160204 6914 160232 17682
rect 161492 16574 161520 19042
rect 162872 16574 162900 24550
rect 167932 24002 167960 92482
rect 168012 82884 168064 82890
rect 168012 82826 168064 82832
rect 168024 28762 168052 82826
rect 168196 77308 168248 77314
rect 168196 77250 168248 77256
rect 168104 74588 168156 74594
rect 168104 74530 168156 74536
rect 168012 28756 168064 28762
rect 168012 28698 168064 28704
rect 168116 25362 168144 74530
rect 168208 28830 168236 77250
rect 168392 39953 168420 151943
rect 168576 150414 168604 171106
rect 169128 170542 169156 282095
rect 169220 264246 169248 354646
rect 169588 289921 169616 401911
rect 169666 398848 169722 398857
rect 169666 398783 169722 398792
rect 169574 289912 169630 289921
rect 169574 289847 169630 289856
rect 169588 277394 169616 289847
rect 169680 286793 169708 398783
rect 169864 362982 169892 431926
rect 170312 429004 170364 429010
rect 170312 428946 170364 428952
rect 170128 423632 170180 423638
rect 170126 423600 170128 423609
rect 170180 423600 170182 423609
rect 170126 423535 170182 423544
rect 170220 408468 170272 408474
rect 170220 408410 170272 408416
rect 169944 398336 169996 398342
rect 169944 398278 169996 398284
rect 169852 362976 169904 362982
rect 169852 362918 169904 362924
rect 169760 361548 169812 361554
rect 169760 361490 169812 361496
rect 169666 286784 169722 286793
rect 169666 286719 169722 286728
rect 169680 285705 169708 286719
rect 169666 285696 169722 285705
rect 169666 285631 169722 285640
rect 169312 277366 169616 277394
rect 169208 264240 169260 264246
rect 169208 264182 169260 264188
rect 169220 264081 169248 264182
rect 169206 264072 169262 264081
rect 169206 264007 169262 264016
rect 169312 177993 169340 277366
rect 169772 204270 169800 361490
rect 169852 356040 169904 356046
rect 169852 355982 169904 355988
rect 169864 355570 169892 355982
rect 169852 355564 169904 355570
rect 169852 355506 169904 355512
rect 169956 354674 169984 398278
rect 170232 356046 170260 408410
rect 170324 363526 170352 428946
rect 170312 363520 170364 363526
rect 170312 363462 170364 363468
rect 170220 356040 170272 356046
rect 170220 355982 170272 355988
rect 169864 354646 169984 354674
rect 169864 347750 169892 354646
rect 169852 347744 169904 347750
rect 169852 347686 169904 347692
rect 169864 347274 169892 347686
rect 169852 347268 169904 347274
rect 169852 347210 169904 347216
rect 169852 258120 169904 258126
rect 169852 258062 169904 258068
rect 169864 251433 169892 258062
rect 169850 251424 169906 251433
rect 169850 251359 169906 251368
rect 169852 245540 169904 245546
rect 169852 245482 169904 245488
rect 169864 244934 169892 245482
rect 169852 244928 169904 244934
rect 169852 244870 169904 244876
rect 169852 234592 169904 234598
rect 169852 234534 169904 234540
rect 169864 233918 169892 234534
rect 169852 233912 169904 233918
rect 169852 233854 169904 233860
rect 170416 229094 170444 463694
rect 170586 454064 170642 454073
rect 170586 453999 170642 454008
rect 170496 452124 170548 452130
rect 170496 452066 170548 452072
rect 170508 451382 170536 452066
rect 170496 451376 170548 451382
rect 170496 451318 170548 451324
rect 170232 229066 170444 229094
rect 170232 227594 170260 229066
rect 170508 229022 170536 451318
rect 170600 233918 170628 453999
rect 170680 452736 170732 452742
rect 170680 452678 170732 452684
rect 170692 244934 170720 452678
rect 170784 398818 170812 586638
rect 170876 400178 170904 587386
rect 171600 587376 171652 587382
rect 171600 587318 171652 587324
rect 171416 587036 171468 587042
rect 171416 586978 171468 586984
rect 171232 584724 171284 584730
rect 171232 584666 171284 584672
rect 171138 584624 171194 584633
rect 171138 584559 171194 584568
rect 170956 563780 171008 563786
rect 170956 563722 171008 563728
rect 170968 409834 170996 563722
rect 171048 455388 171100 455394
rect 171048 455330 171100 455336
rect 171060 449818 171088 455330
rect 171048 449812 171100 449818
rect 171048 449754 171100 449760
rect 170956 409828 171008 409834
rect 170956 409770 171008 409776
rect 170864 400172 170916 400178
rect 170864 400114 170916 400120
rect 170772 398812 170824 398818
rect 170772 398754 170824 398760
rect 170956 363588 171008 363594
rect 170956 363530 171008 363536
rect 170772 362364 170824 362370
rect 170772 362306 170824 362312
rect 170784 361729 170812 362306
rect 170770 361720 170826 361729
rect 170770 361655 170826 361664
rect 170680 244928 170732 244934
rect 170680 244870 170732 244876
rect 170588 233912 170640 233918
rect 170588 233854 170640 233860
rect 170496 229016 170548 229022
rect 170496 228958 170548 228964
rect 170508 228614 170536 228958
rect 170496 228608 170548 228614
rect 170496 228550 170548 228556
rect 170220 227588 170272 227594
rect 170220 227530 170272 227536
rect 170232 227186 170260 227530
rect 170220 227180 170272 227186
rect 170220 227122 170272 227128
rect 170784 213246 170812 361655
rect 170968 361010 170996 363530
rect 171060 361146 171088 449754
rect 171048 361140 171100 361146
rect 171048 361082 171100 361088
rect 170956 361004 171008 361010
rect 170956 360946 171008 360952
rect 170864 351416 170916 351422
rect 170864 351358 170916 351364
rect 170772 213240 170824 213246
rect 170772 213182 170824 213188
rect 170772 210452 170824 210458
rect 170772 210394 170824 210400
rect 169760 204264 169812 204270
rect 169760 204206 169812 204212
rect 170496 182844 170548 182850
rect 170496 182786 170548 182792
rect 170404 181484 170456 181490
rect 170404 181426 170456 181432
rect 169298 177984 169354 177993
rect 169298 177919 169354 177928
rect 169312 177410 169340 177919
rect 169300 177404 169352 177410
rect 169300 177346 169352 177352
rect 169208 175976 169260 175982
rect 169208 175918 169260 175924
rect 169116 170536 169168 170542
rect 169116 170478 169168 170484
rect 169024 170400 169076 170406
rect 169024 170342 169076 170348
rect 168748 151088 168800 151094
rect 168748 151030 168800 151036
rect 168564 150408 168616 150414
rect 168562 150376 168564 150385
rect 168616 150376 168618 150385
rect 168562 150311 168618 150320
rect 168470 150104 168526 150113
rect 168470 150039 168526 150048
rect 168378 39944 168434 39953
rect 168378 39879 168434 39888
rect 168484 38185 168512 150039
rect 168576 136882 168604 150311
rect 168760 150113 168788 151030
rect 168746 150104 168802 150113
rect 168746 150039 168802 150048
rect 169036 138990 169064 170342
rect 169128 170241 169156 170478
rect 169114 170232 169170 170241
rect 169114 170167 169170 170176
rect 169116 164892 169168 164898
rect 169116 164834 169168 164840
rect 169128 153105 169156 164834
rect 169114 153096 169170 153105
rect 169114 153031 169170 153040
rect 169024 138984 169076 138990
rect 169024 138926 169076 138932
rect 169220 138786 169248 175918
rect 169208 138780 169260 138786
rect 169208 138722 169260 138728
rect 168564 136876 168616 136882
rect 168564 136818 168616 136824
rect 168564 117292 168616 117298
rect 168564 117234 168616 117240
rect 168576 38457 168604 117234
rect 169024 84244 169076 84250
rect 169024 84186 169076 84192
rect 168840 69692 168892 69698
rect 168840 69634 168892 69640
rect 168852 67017 168880 69634
rect 168838 67008 168894 67017
rect 168838 66943 168894 66952
rect 168840 66224 168892 66230
rect 168840 66166 168892 66172
rect 168852 66065 168880 66166
rect 168838 66056 168894 66065
rect 168838 65991 168894 66000
rect 168840 64864 168892 64870
rect 168840 64806 168892 64812
rect 168852 63889 168880 64806
rect 168932 64184 168984 64190
rect 168932 64126 168984 64132
rect 168838 63880 168894 63889
rect 168838 63815 168894 63824
rect 168840 61396 168892 61402
rect 168840 61338 168892 61344
rect 168852 60081 168880 61338
rect 168944 61169 168972 64126
rect 168930 61160 168986 61169
rect 168930 61095 168986 61104
rect 168838 60072 168894 60081
rect 168838 60007 168894 60016
rect 168840 59356 168892 59362
rect 168840 59298 168892 59304
rect 168852 58313 168880 59298
rect 168838 58304 168894 58313
rect 168838 58239 168894 58248
rect 168562 38448 168618 38457
rect 168562 38383 168618 38392
rect 168470 38176 168526 38185
rect 168470 38111 168526 38120
rect 168380 31068 168432 31074
rect 168380 31010 168432 31016
rect 168196 28824 168248 28830
rect 168196 28766 168248 28772
rect 168104 25356 168156 25362
rect 168104 25298 168156 25304
rect 167920 23996 167972 24002
rect 167920 23938 167972 23944
rect 165620 23316 165672 23322
rect 165620 23258 165672 23264
rect 164240 23180 164292 23186
rect 164240 23122 164292 23128
rect 164252 16574 164280 23122
rect 165632 16574 165660 23258
rect 167000 23248 167052 23254
rect 167000 23190 167052 23196
rect 167012 16574 167040 23190
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11688 161348 11694
rect 161296 11630 161348 11636
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11630
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 3466 168420 31010
rect 169036 28694 169064 84186
rect 169116 78736 169168 78742
rect 169116 78678 169168 78684
rect 169024 28688 169076 28694
rect 169024 28630 169076 28636
rect 169128 26178 169156 78678
rect 169208 73228 169260 73234
rect 169208 73170 169260 73176
rect 169116 26172 169168 26178
rect 169116 26114 169168 26120
rect 169220 25498 169248 73170
rect 169392 63504 169444 63510
rect 169392 63446 169444 63452
rect 169404 62937 169432 63446
rect 169390 62928 169446 62937
rect 169390 62863 169446 62872
rect 169300 59424 169352 59430
rect 169300 59366 169352 59372
rect 169312 28082 169340 59366
rect 169392 31272 169444 31278
rect 169392 31214 169444 31220
rect 169300 28076 169352 28082
rect 169300 28018 169352 28024
rect 169208 25492 169260 25498
rect 169208 25434 169260 25440
rect 169404 4010 169432 31214
rect 170416 26217 170444 181426
rect 170508 27305 170536 182786
rect 170680 174548 170732 174554
rect 170680 174490 170732 174496
rect 170588 160744 170640 160750
rect 170588 160686 170640 160692
rect 170600 28801 170628 160686
rect 170586 28792 170642 28801
rect 170586 28727 170642 28736
rect 170494 27296 170550 27305
rect 170494 27231 170550 27240
rect 170692 26897 170720 174490
rect 170784 140350 170812 210394
rect 170876 204950 170904 351358
rect 170968 215966 170996 360946
rect 171152 340882 171180 584559
rect 171244 354686 171272 584666
rect 171324 584588 171376 584594
rect 171324 584530 171376 584536
rect 171336 408474 171364 584530
rect 171428 423570 171456 586978
rect 171508 584248 171560 584254
rect 171508 584190 171560 584196
rect 171520 429010 171548 584190
rect 171612 455394 171640 587318
rect 172150 587208 172206 587217
rect 172150 587143 172206 587152
rect 171784 474972 171836 474978
rect 171784 474914 171836 474920
rect 171600 455388 171652 455394
rect 171600 455330 171652 455336
rect 171508 429004 171560 429010
rect 171508 428946 171560 428952
rect 171416 423564 171468 423570
rect 171416 423506 171468 423512
rect 171428 422346 171456 423506
rect 171416 422340 171468 422346
rect 171416 422282 171468 422288
rect 171324 408468 171376 408474
rect 171324 408410 171376 408416
rect 171232 354680 171284 354686
rect 171232 354622 171284 354628
rect 171140 340876 171192 340882
rect 171140 340818 171192 340824
rect 171692 340876 171744 340882
rect 171692 340818 171744 340824
rect 171704 340474 171732 340818
rect 171692 340468 171744 340474
rect 171692 340410 171744 340416
rect 171048 271924 171100 271930
rect 171048 271866 171100 271872
rect 171060 253774 171088 271866
rect 171692 263628 171744 263634
rect 171692 263570 171744 263576
rect 171048 253768 171100 253774
rect 171048 253710 171100 253716
rect 171704 253094 171732 263570
rect 171692 253088 171744 253094
rect 171692 253030 171744 253036
rect 171796 233238 171824 474914
rect 171876 455524 171928 455530
rect 171876 455466 171928 455472
rect 171784 233232 171836 233238
rect 171784 233174 171836 233180
rect 171140 231124 171192 231130
rect 171140 231066 171192 231072
rect 171048 217320 171100 217326
rect 171048 217262 171100 217268
rect 170956 215960 171008 215966
rect 170956 215902 171008 215908
rect 170956 206304 171008 206310
rect 170956 206246 171008 206252
rect 170864 204944 170916 204950
rect 170864 204886 170916 204892
rect 170772 140344 170824 140350
rect 170772 140286 170824 140292
rect 170968 138718 170996 206246
rect 171060 140282 171088 217262
rect 171048 140276 171100 140282
rect 171048 140218 171100 140224
rect 170956 138712 171008 138718
rect 170956 138654 171008 138660
rect 170956 63572 171008 63578
rect 170956 63514 171008 63520
rect 170772 57452 170824 57458
rect 170772 57394 170824 57400
rect 170678 26888 170734 26897
rect 170678 26823 170734 26832
rect 170402 26208 170458 26217
rect 170402 26143 170458 26152
rect 170784 10742 170812 57394
rect 170864 57248 170916 57254
rect 170864 57190 170916 57196
rect 170876 23390 170904 57190
rect 170968 29102 170996 63514
rect 170956 29096 171008 29102
rect 170956 29038 171008 29044
rect 171152 24818 171180 231066
rect 171888 227662 171916 455466
rect 172060 454096 172112 454102
rect 172060 454038 172112 454044
rect 171968 452192 172020 452198
rect 171968 452134 172020 452140
rect 171980 451450 172008 452134
rect 171968 451444 172020 451450
rect 171968 451386 172020 451392
rect 171980 235890 172008 451386
rect 172072 244186 172100 454038
rect 172164 427650 172192 587143
rect 172796 586832 172848 586838
rect 172796 586774 172848 586780
rect 172520 584792 172572 584798
rect 172520 584734 172572 584740
rect 172426 475280 172482 475289
rect 172426 475215 172482 475224
rect 172440 474978 172468 475215
rect 172428 474972 172480 474978
rect 172428 474914 172480 474920
rect 172428 456136 172480 456142
rect 172428 456078 172480 456084
rect 172440 455530 172468 456078
rect 172428 455524 172480 455530
rect 172428 455466 172480 455472
rect 172428 454844 172480 454850
rect 172428 454786 172480 454792
rect 172440 454102 172468 454786
rect 172428 454096 172480 454102
rect 172428 454038 172480 454044
rect 172152 427644 172204 427650
rect 172152 427586 172204 427592
rect 172336 426420 172388 426426
rect 172336 426362 172388 426368
rect 172152 421116 172204 421122
rect 172152 421058 172204 421064
rect 172060 244180 172112 244186
rect 172060 244122 172112 244128
rect 171968 235884 172020 235890
rect 171968 235826 172020 235832
rect 171876 227656 171928 227662
rect 171876 227598 171928 227604
rect 172164 227050 172192 421058
rect 172244 421048 172296 421054
rect 172244 420990 172296 420996
rect 172256 338910 172284 420990
rect 172348 364002 172376 426362
rect 172336 363996 172388 364002
rect 172336 363938 172388 363944
rect 172428 354680 172480 354686
rect 172428 354622 172480 354628
rect 172440 354210 172468 354622
rect 172428 354204 172480 354210
rect 172428 354146 172480 354152
rect 172336 351348 172388 351354
rect 172336 351290 172388 351296
rect 172244 338904 172296 338910
rect 172244 338846 172296 338852
rect 172348 309126 172376 351290
rect 172532 346322 172560 584734
rect 172612 584656 172664 584662
rect 172612 584598 172664 584604
rect 172624 358698 172652 584598
rect 172704 453892 172756 453898
rect 172704 453834 172756 453840
rect 172716 452878 172744 453834
rect 172704 452872 172756 452878
rect 172704 452814 172756 452820
rect 172612 358692 172664 358698
rect 172612 358634 172664 358640
rect 172520 346316 172572 346322
rect 172520 346258 172572 346264
rect 172428 345704 172480 345710
rect 172428 345646 172480 345652
rect 172440 328438 172468 345646
rect 172428 328432 172480 328438
rect 172428 328374 172480 328380
rect 172336 309120 172388 309126
rect 172336 309062 172388 309068
rect 172244 294024 172296 294030
rect 172244 293966 172296 293972
rect 172256 253366 172284 293966
rect 172336 285728 172388 285734
rect 172336 285670 172388 285676
rect 172244 253360 172296 253366
rect 172244 253302 172296 253308
rect 172348 251122 172376 285670
rect 172428 274712 172480 274718
rect 172428 274654 172480 274660
rect 172336 251116 172388 251122
rect 172336 251058 172388 251064
rect 172440 250782 172468 274654
rect 172428 250776 172480 250782
rect 172428 250718 172480 250724
rect 172428 235884 172480 235890
rect 172428 235826 172480 235832
rect 172440 235346 172468 235826
rect 172428 235340 172480 235346
rect 172428 235282 172480 235288
rect 172716 234530 172744 452814
rect 172808 427689 172836 586774
rect 172888 585132 172940 585138
rect 172888 585074 172940 585080
rect 172794 427680 172850 427689
rect 172794 427615 172850 427624
rect 172900 426426 172928 585074
rect 173070 455696 173126 455705
rect 173070 455631 173126 455640
rect 172888 426420 172940 426426
rect 172888 426362 172940 426368
rect 172704 234524 172756 234530
rect 172704 234466 172756 234472
rect 172428 233232 172480 233238
rect 172428 233174 172480 233180
rect 172440 232626 172468 233174
rect 172428 232620 172480 232626
rect 172428 232562 172480 232568
rect 173084 231810 173112 455631
rect 173176 426358 173204 587415
rect 173532 586764 173584 586770
rect 173532 586706 173584 586712
rect 173256 584384 173308 584390
rect 173256 584326 173308 584332
rect 173268 438870 173296 584326
rect 173544 460934 173572 586706
rect 174636 586628 174688 586634
rect 174636 586570 174688 586576
rect 173990 584352 174046 584361
rect 173990 584287 174046 584296
rect 173900 475312 173952 475318
rect 173900 475254 173952 475260
rect 173544 460906 173848 460934
rect 173440 453824 173492 453830
rect 173440 453766 173492 453772
rect 173452 452810 173480 453766
rect 173440 452804 173492 452810
rect 173440 452746 173492 452752
rect 173256 438864 173308 438870
rect 173256 438806 173308 438812
rect 173164 426352 173216 426358
rect 173164 426294 173216 426300
rect 173164 421252 173216 421258
rect 173164 421194 173216 421200
rect 173072 231804 173124 231810
rect 173072 231746 173124 231752
rect 172428 227656 172480 227662
rect 172428 227598 172480 227604
rect 172440 227118 172468 227598
rect 172428 227112 172480 227118
rect 172428 227054 172480 227060
rect 172152 227044 172204 227050
rect 172152 226986 172204 226992
rect 171784 225616 171836 225622
rect 171784 225558 171836 225564
rect 171796 140894 171824 225558
rect 171876 222896 171928 222902
rect 171876 222838 171928 222844
rect 171784 140888 171836 140894
rect 171784 140830 171836 140836
rect 171888 139058 171916 222838
rect 171876 139052 171928 139058
rect 171876 138994 171928 139000
rect 171784 123480 171836 123486
rect 171784 123422 171836 123428
rect 171796 113150 171824 123422
rect 173176 113898 173204 421194
rect 173256 421184 173308 421190
rect 173256 421126 173308 421132
rect 173268 115394 173296 421126
rect 173452 241398 173480 452746
rect 173820 451178 173848 460906
rect 173808 451172 173860 451178
rect 173808 451114 173860 451120
rect 173624 427848 173676 427854
rect 173624 427790 173676 427796
rect 173532 420980 173584 420986
rect 173532 420922 173584 420928
rect 173544 338842 173572 420922
rect 173636 363934 173664 427790
rect 173716 427780 173768 427786
rect 173716 427722 173768 427728
rect 173728 427689 173756 427722
rect 173714 427680 173770 427689
rect 173714 427615 173770 427624
rect 173624 363928 173676 363934
rect 173624 363870 173676 363876
rect 173820 360126 173848 451114
rect 173808 360120 173860 360126
rect 173808 360062 173860 360068
rect 173808 358692 173860 358698
rect 173808 358634 173860 358640
rect 173820 358086 173848 358634
rect 173808 358080 173860 358086
rect 173808 358022 173860 358028
rect 173716 354000 173768 354006
rect 173716 353942 173768 353948
rect 173624 344480 173676 344486
rect 173624 344422 173676 344428
rect 173532 338836 173584 338842
rect 173532 338778 173584 338784
rect 173636 310486 173664 344422
rect 173728 325650 173756 353942
rect 173808 346316 173860 346322
rect 173808 346258 173860 346264
rect 173820 345710 173848 346258
rect 173808 345704 173860 345710
rect 173808 345646 173860 345652
rect 173716 325644 173768 325650
rect 173716 325586 173768 325592
rect 173624 310480 173676 310486
rect 173624 310422 173676 310428
rect 173532 299532 173584 299538
rect 173532 299474 173584 299480
rect 173544 253230 173572 299474
rect 173624 292596 173676 292602
rect 173624 292538 173676 292544
rect 173532 253224 173584 253230
rect 173532 253166 173584 253172
rect 173636 252278 173664 292538
rect 173716 276072 173768 276078
rect 173716 276014 173768 276020
rect 173624 252272 173676 252278
rect 173624 252214 173676 252220
rect 173728 250986 173756 276014
rect 173716 250980 173768 250986
rect 173716 250922 173768 250928
rect 173440 241392 173492 241398
rect 173440 241334 173492 241340
rect 173808 241392 173860 241398
rect 173808 241334 173860 241340
rect 173820 240786 173848 241334
rect 173808 240780 173860 240786
rect 173808 240722 173860 240728
rect 173912 240038 173940 475254
rect 174004 350538 174032 584287
rect 174084 453620 174136 453626
rect 174084 453562 174136 453568
rect 174096 453014 174124 453562
rect 174544 453484 174596 453490
rect 174544 453426 174596 453432
rect 174556 453150 174584 453426
rect 174544 453144 174596 453150
rect 174544 453086 174596 453092
rect 174084 453008 174136 453014
rect 174084 452950 174136 452956
rect 173992 350532 174044 350538
rect 173992 350474 174044 350480
rect 173900 240032 173952 240038
rect 173900 239974 173952 239980
rect 173912 239290 173940 239974
rect 173900 239284 173952 239290
rect 173900 239226 173952 239232
rect 174096 237386 174124 452950
rect 174176 449200 174228 449206
rect 174176 449142 174228 449148
rect 174188 393310 174216 449142
rect 174176 393304 174228 393310
rect 174176 393246 174228 393252
rect 174556 249694 174584 453086
rect 174648 398750 174676 586570
rect 174728 585812 174780 585818
rect 174728 585754 174780 585760
rect 174636 398744 174688 398750
rect 174636 398686 174688 398692
rect 174740 397458 174768 585754
rect 175372 584996 175424 585002
rect 175372 584938 175424 584944
rect 174912 475312 174964 475318
rect 174912 475254 174964 475260
rect 174924 474774 174952 475254
rect 175292 475046 175320 475077
rect 175280 475040 175332 475046
rect 175278 475008 175280 475017
rect 175332 475008 175334 475017
rect 175278 474943 175334 474952
rect 174912 474768 174964 474774
rect 174912 474710 174964 474716
rect 174820 470008 174872 470014
rect 174820 469950 174872 469956
rect 174728 397452 174780 397458
rect 174728 397394 174780 397400
rect 174728 359576 174780 359582
rect 174728 359518 174780 359524
rect 174636 355564 174688 355570
rect 174636 355506 174688 355512
rect 174544 249688 174596 249694
rect 174544 249630 174596 249636
rect 174084 237380 174136 237386
rect 174084 237322 174136 237328
rect 174096 236026 174124 237322
rect 174084 236020 174136 236026
rect 174084 235962 174136 235968
rect 174544 236020 174596 236026
rect 174544 235962 174596 235968
rect 173348 234524 173400 234530
rect 173348 234466 173400 234472
rect 173360 177342 173388 234466
rect 173440 196648 173492 196654
rect 173440 196590 173492 196596
rect 173348 177336 173400 177342
rect 173348 177278 173400 177284
rect 173256 115388 173308 115394
rect 173256 115330 173308 115336
rect 173164 113892 173216 113898
rect 173164 113834 173216 113840
rect 171784 113144 171836 113150
rect 171784 113086 171836 113092
rect 173164 85604 173216 85610
rect 173164 85546 173216 85552
rect 171784 75948 171836 75954
rect 171784 75890 171836 75896
rect 171232 55888 171284 55894
rect 171232 55830 171284 55836
rect 171140 24812 171192 24818
rect 171140 24754 171192 24760
rect 170864 23384 170916 23390
rect 170864 23326 170916 23332
rect 171244 16574 171272 55830
rect 171796 26110 171824 75890
rect 172060 60784 172112 60790
rect 172060 60726 172112 60732
rect 171968 57724 172020 57730
rect 171968 57666 172020 57672
rect 171876 57588 171928 57594
rect 171876 57530 171928 57536
rect 171784 26104 171836 26110
rect 171784 26046 171836 26052
rect 171888 18970 171916 57530
rect 171980 21690 172008 57666
rect 172072 28150 172100 60726
rect 172520 44872 172572 44878
rect 172520 44814 172572 44820
rect 172152 33856 172204 33862
rect 172152 33798 172204 33804
rect 172060 28144 172112 28150
rect 172060 28086 172112 28092
rect 171968 21684 172020 21690
rect 171968 21626 172020 21632
rect 171876 18964 171928 18970
rect 171876 18906 171928 18912
rect 171244 16546 172008 16574
rect 170772 10736 170824 10742
rect 170772 10678 170824 10684
rect 170312 10668 170364 10674
rect 170312 10610 170364 10616
rect 169392 4004 169444 4010
rect 169392 3946 169444 3952
rect 168380 3460 168432 3466
rect 168380 3402 168432 3408
rect 169576 3460 169628 3466
rect 169576 3402 169628 3408
rect 168380 3324 168432 3330
rect 168380 3266 168432 3272
rect 168392 480 168420 3266
rect 169588 480 169616 3402
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 10610
rect 171980 480 172008 16546
rect 172164 3670 172192 33798
rect 172532 16574 172560 44814
rect 173176 24750 173204 85546
rect 173256 81456 173308 81462
rect 173256 81398 173308 81404
rect 173164 24744 173216 24750
rect 173164 24686 173216 24692
rect 173268 23934 173296 81398
rect 173256 23928 173308 23934
rect 173256 23870 173308 23876
rect 173360 22574 173388 177278
rect 173452 140554 173480 196590
rect 174556 180130 174584 235962
rect 174648 228478 174676 355506
rect 174740 302190 174768 359518
rect 174832 349110 174860 469950
rect 174912 460216 174964 460222
rect 174912 460158 174964 460164
rect 174924 365634 174952 460158
rect 175004 451988 175056 451994
rect 175004 451930 175056 451936
rect 175016 376718 175044 451930
rect 175188 449404 175240 449410
rect 175188 449346 175240 449352
rect 175200 449206 175228 449346
rect 175188 449200 175240 449206
rect 175188 449142 175240 449148
rect 175004 376712 175056 376718
rect 175004 376654 175056 376660
rect 174912 365628 174964 365634
rect 174912 365570 174964 365576
rect 174912 352572 174964 352578
rect 174912 352514 174964 352520
rect 174820 349104 174872 349110
rect 174820 349046 174872 349052
rect 174820 347132 174872 347138
rect 174820 347074 174872 347080
rect 174832 311846 174860 347074
rect 174924 332586 174952 352514
rect 175188 350532 175240 350538
rect 175188 350474 175240 350480
rect 175200 350062 175228 350474
rect 175188 350056 175240 350062
rect 175188 349998 175240 350004
rect 174912 332580 174964 332586
rect 174912 332522 174964 332528
rect 174820 311840 174872 311846
rect 174820 311782 174872 311788
rect 174728 302184 174780 302190
rect 174728 302126 174780 302132
rect 174728 298172 174780 298178
rect 174728 298114 174780 298120
rect 174740 251598 174768 298114
rect 174820 288448 174872 288454
rect 174820 288390 174872 288396
rect 174728 251592 174780 251598
rect 174728 251534 174780 251540
rect 174832 251190 174860 288390
rect 174912 276140 174964 276146
rect 174912 276082 174964 276088
rect 174820 251184 174872 251190
rect 174820 251126 174872 251132
rect 174924 250850 174952 276082
rect 175004 251864 175056 251870
rect 175004 251806 175056 251812
rect 174912 250844 174964 250850
rect 174912 250786 174964 250792
rect 174728 239284 174780 239290
rect 174728 239226 174780 239232
rect 174636 228472 174688 228478
rect 174636 228414 174688 228420
rect 174544 180124 174596 180130
rect 174544 180066 174596 180072
rect 173440 140548 173492 140554
rect 173440 140490 173492 140496
rect 173440 71800 173492 71806
rect 173440 71742 173492 71748
rect 173452 25430 173480 71742
rect 173532 49020 173584 49026
rect 173532 48962 173584 48968
rect 173440 25424 173492 25430
rect 173440 25366 173492 25372
rect 173348 22568 173400 22574
rect 173348 22510 173400 22516
rect 172532 16546 172744 16574
rect 172152 3664 172204 3670
rect 172152 3606 172204 3612
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173544 3874 173572 48962
rect 174556 21350 174584 180066
rect 174636 172508 174688 172514
rect 174636 172450 174688 172456
rect 174648 27033 174676 172450
rect 174740 167686 174768 239226
rect 175016 238066 175044 251806
rect 175188 249688 175240 249694
rect 175188 249630 175240 249636
rect 175200 249082 175228 249630
rect 175188 249076 175240 249082
rect 175188 249018 175240 249024
rect 175292 240106 175320 474943
rect 175384 429146 175412 584938
rect 176200 567860 176252 567866
rect 176200 567802 176252 567808
rect 175924 475380 175976 475386
rect 175924 475322 175976 475328
rect 175936 474842 175964 475322
rect 175924 474836 175976 474842
rect 175924 474778 175976 474784
rect 175372 429140 175424 429146
rect 175372 429082 175424 429088
rect 175384 427854 175412 429082
rect 175372 427848 175424 427854
rect 175372 427790 175424 427796
rect 175280 240100 175332 240106
rect 175280 240042 175332 240048
rect 175004 238060 175056 238066
rect 175004 238002 175056 238008
rect 174820 218748 174872 218754
rect 174820 218690 174872 218696
rect 174728 167680 174780 167686
rect 174728 167622 174780 167628
rect 174740 28218 174768 167622
rect 174832 139194 174860 218690
rect 174912 193860 174964 193866
rect 174912 193802 174964 193808
rect 174924 140622 174952 193802
rect 175292 182170 175320 240042
rect 175936 237318 175964 474778
rect 176108 454776 176160 454782
rect 176108 454718 176160 454724
rect 176120 454170 176148 454718
rect 176108 454164 176160 454170
rect 176108 454106 176160 454112
rect 176016 453960 176068 453966
rect 176016 453902 176068 453908
rect 176028 452674 176056 453902
rect 176016 452668 176068 452674
rect 176016 452610 176068 452616
rect 176028 244118 176056 452610
rect 176120 248402 176148 454106
rect 176212 396030 176240 567802
rect 176660 475244 176712 475250
rect 176660 475186 176712 475192
rect 176672 475153 176700 475186
rect 176658 475144 176714 475153
rect 176658 475079 176714 475088
rect 176292 467288 176344 467294
rect 176292 467230 176344 467236
rect 176200 396024 176252 396030
rect 176200 395966 176252 395972
rect 176304 351898 176332 467230
rect 176476 463752 176528 463758
rect 176476 463694 176528 463700
rect 176384 458856 176436 458862
rect 176384 458798 176436 458804
rect 176396 364342 176424 458798
rect 176488 452606 176516 463694
rect 176476 452600 176528 452606
rect 176476 452542 176528 452548
rect 176384 364336 176436 364342
rect 176384 364278 176436 364284
rect 176384 360868 176436 360874
rect 176384 360810 176436 360816
rect 176292 351892 176344 351898
rect 176292 351834 176344 351840
rect 176292 349920 176344 349926
rect 176292 349862 176344 349868
rect 176200 341556 176252 341562
rect 176200 341498 176252 341504
rect 176108 248396 176160 248402
rect 176108 248338 176160 248344
rect 176120 247110 176148 248338
rect 176108 247104 176160 247110
rect 176108 247046 176160 247052
rect 176016 244112 176068 244118
rect 176016 244054 176068 244060
rect 176028 243574 176056 244054
rect 176016 243568 176068 243574
rect 176016 243510 176068 243516
rect 175924 237312 175976 237318
rect 175924 237254 175976 237260
rect 175936 236774 175964 237254
rect 175924 236768 175976 236774
rect 175924 236710 175976 236716
rect 176108 228540 176160 228546
rect 176108 228482 176160 228488
rect 175280 182164 175332 182170
rect 175280 182106 175332 182112
rect 175740 182164 175792 182170
rect 175740 182106 175792 182112
rect 175752 181490 175780 182106
rect 175740 181484 175792 181490
rect 175740 181426 175792 181432
rect 175004 174616 175056 174622
rect 175004 174558 175056 174564
rect 175016 146266 175044 174558
rect 175924 153876 175976 153882
rect 175924 153818 175976 153824
rect 175004 146260 175056 146266
rect 175004 146202 175056 146208
rect 174912 140616 174964 140622
rect 174912 140558 174964 140564
rect 174820 139188 174872 139194
rect 174820 139130 174872 139136
rect 174820 129056 174872 129062
rect 174820 128998 174872 129004
rect 174832 107642 174860 128998
rect 174912 124908 174964 124914
rect 174912 124850 174964 124856
rect 174820 107636 174872 107642
rect 174820 107578 174872 107584
rect 174924 104854 174952 124850
rect 174912 104848 174964 104854
rect 174912 104790 174964 104796
rect 174820 87032 174872 87038
rect 174820 86974 174872 86980
rect 174832 28626 174860 86974
rect 174912 81524 174964 81530
rect 174912 81466 174964 81472
rect 174820 28620 174872 28626
rect 174820 28562 174872 28568
rect 174728 28212 174780 28218
rect 174728 28154 174780 28160
rect 174634 27024 174690 27033
rect 174634 26959 174690 26968
rect 174924 24682 174952 81466
rect 175004 80096 175056 80102
rect 175004 80038 175056 80044
rect 175016 26246 175044 80038
rect 175096 57656 175148 57662
rect 175096 57598 175148 57604
rect 175004 26240 175056 26246
rect 175004 26182 175056 26188
rect 174912 24676 174964 24682
rect 174912 24618 174964 24624
rect 174544 21344 174596 21350
rect 174544 21286 174596 21292
rect 173900 10736 173952 10742
rect 173900 10678 173952 10684
rect 173532 3868 173584 3874
rect 173532 3810 173584 3816
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 10678
rect 175108 3738 175136 57598
rect 175188 57316 175240 57322
rect 175188 57258 175240 57264
rect 175200 10810 175228 57258
rect 175936 26926 175964 153818
rect 176016 152516 176068 152522
rect 176016 152458 176068 152464
rect 176028 27538 176056 152458
rect 176120 140826 176148 228482
rect 176212 213994 176240 341498
rect 176304 313274 176332 349862
rect 176396 333946 176424 360810
rect 176384 333940 176436 333946
rect 176384 333882 176436 333888
rect 176292 313268 176344 313274
rect 176292 313210 176344 313216
rect 176292 287156 176344 287162
rect 176292 287098 176344 287104
rect 176304 252210 176332 287098
rect 176384 263696 176436 263702
rect 176384 263638 176436 263644
rect 176396 253162 176424 263638
rect 176384 253156 176436 253162
rect 176384 253098 176436 253104
rect 176292 252204 176344 252210
rect 176292 252146 176344 252152
rect 176672 248266 176700 475079
rect 177316 442338 177344 700470
rect 184204 700460 184256 700466
rect 184204 700402 184256 700408
rect 178776 683188 178828 683194
rect 178776 683130 178828 683136
rect 178040 584860 178092 584866
rect 178040 584802 178092 584808
rect 177488 576224 177540 576230
rect 177488 576166 177540 576172
rect 177396 472796 177448 472802
rect 177396 472738 177448 472744
rect 177408 472054 177436 472738
rect 177396 472048 177448 472054
rect 177396 471990 177448 471996
rect 177304 442332 177356 442338
rect 177304 442274 177356 442280
rect 177304 427848 177356 427854
rect 177304 427790 177356 427796
rect 177316 363798 177344 427790
rect 177304 363792 177356 363798
rect 177304 363734 177356 363740
rect 177304 362228 177356 362234
rect 177304 362170 177356 362176
rect 176752 360120 176804 360126
rect 176752 360062 176804 360068
rect 176660 248260 176712 248266
rect 176660 248202 176712 248208
rect 176672 247178 176700 248202
rect 176660 247172 176712 247178
rect 176660 247114 176712 247120
rect 176764 219434 176792 360062
rect 176844 340332 176896 340338
rect 176844 340274 176896 340280
rect 176856 336734 176884 340274
rect 176844 336728 176896 336734
rect 176844 336670 176896 336676
rect 177316 315994 177344 362170
rect 177304 315988 177356 315994
rect 177304 315930 177356 315936
rect 177304 295384 177356 295390
rect 177304 295326 177356 295332
rect 177316 252414 177344 295326
rect 177304 252408 177356 252414
rect 177304 252350 177356 252356
rect 176844 249620 176896 249626
rect 176844 249562 176896 249568
rect 176856 249150 176884 249562
rect 177408 249150 177436 471990
rect 177500 393310 177528 576166
rect 177580 573436 177632 573442
rect 177580 573378 177632 573384
rect 177592 415410 177620 573378
rect 177764 465724 177816 465730
rect 177764 465666 177816 465672
rect 177672 464432 177724 464438
rect 177672 464374 177724 464380
rect 177580 415404 177632 415410
rect 177580 415346 177632 415352
rect 177488 393304 177540 393310
rect 177488 393246 177540 393252
rect 177684 360126 177712 464374
rect 177776 372570 177804 465666
rect 178052 429078 178080 584802
rect 178684 486464 178736 486470
rect 178684 486406 178736 486412
rect 178040 429072 178092 429078
rect 178040 429014 178092 429020
rect 177856 428528 177908 428534
rect 177856 428470 177908 428476
rect 177764 372564 177816 372570
rect 177764 372506 177816 372512
rect 177868 363594 177896 428470
rect 178052 427854 178080 429014
rect 178040 427848 178092 427854
rect 178040 427790 178092 427796
rect 177856 363588 177908 363594
rect 177856 363530 177908 363536
rect 177672 360120 177724 360126
rect 177672 360062 177724 360068
rect 177488 342984 177540 342990
rect 177488 342926 177540 342932
rect 177500 304978 177528 342926
rect 177488 304972 177540 304978
rect 177488 304914 177540 304920
rect 177488 277432 177540 277438
rect 177488 277374 177540 277380
rect 177500 251054 177528 277374
rect 177488 251048 177540 251054
rect 177488 250990 177540 250996
rect 176844 249144 176896 249150
rect 176844 249086 176896 249092
rect 177396 249144 177448 249150
rect 177396 249086 177448 249092
rect 177396 247172 177448 247178
rect 177396 247114 177448 247120
rect 177304 247104 177356 247110
rect 177304 247046 177356 247052
rect 176672 219406 176792 219434
rect 176200 213988 176252 213994
rect 176200 213930 176252 213936
rect 176672 211138 176700 219406
rect 176660 211132 176712 211138
rect 176660 211074 176712 211080
rect 176672 210458 176700 211074
rect 176660 210452 176712 210458
rect 176660 210394 176712 210400
rect 176200 208344 176252 208350
rect 176200 208286 176252 208292
rect 176212 141234 176240 208286
rect 177316 184210 177344 247046
rect 177304 184204 177356 184210
rect 177304 184146 177356 184152
rect 176200 141228 176252 141234
rect 176200 141170 176252 141176
rect 176108 140820 176160 140826
rect 176108 140762 176160 140768
rect 176108 91112 176160 91118
rect 176108 91054 176160 91060
rect 176120 28422 176148 91054
rect 176200 88392 176252 88398
rect 176200 88334 176252 88340
rect 176212 28558 176240 88334
rect 176292 70440 176344 70446
rect 176292 70382 176344 70388
rect 176200 28552 176252 28558
rect 176200 28494 176252 28500
rect 176108 28416 176160 28422
rect 176108 28358 176160 28364
rect 176016 27532 176068 27538
rect 176016 27474 176068 27480
rect 176304 27402 176332 70382
rect 176660 42084 176712 42090
rect 176660 42026 176712 42032
rect 176292 27396 176344 27402
rect 176292 27338 176344 27344
rect 175924 26920 175976 26926
rect 175924 26862 175976 26868
rect 175280 18964 175332 18970
rect 175280 18906 175332 18912
rect 175292 16574 175320 18906
rect 175292 16546 175504 16574
rect 175188 10804 175240 10810
rect 175188 10746 175240 10752
rect 175096 3732 175148 3738
rect 175096 3674 175148 3680
rect 175476 480 175504 16546
rect 176672 480 176700 42026
rect 177316 27441 177344 184146
rect 177408 170474 177436 247114
rect 178696 238066 178724 486406
rect 178788 443698 178816 683130
rect 181536 585880 181588 585886
rect 181536 585822 181588 585828
rect 180800 584928 180852 584934
rect 180800 584870 180852 584876
rect 178960 583024 179012 583030
rect 178960 582966 179012 582972
rect 178866 453248 178922 453257
rect 178866 453183 178922 453192
rect 178776 443692 178828 443698
rect 178776 443634 178828 443640
rect 178776 428460 178828 428466
rect 178776 428402 178828 428408
rect 178788 364206 178816 428402
rect 178776 364200 178828 364206
rect 178776 364142 178828 364148
rect 178776 355496 178828 355502
rect 178776 355438 178828 355444
rect 178684 238060 178736 238066
rect 178684 238002 178736 238008
rect 178040 233232 178092 233238
rect 178040 233174 178092 233180
rect 177580 228608 177632 228614
rect 177580 228550 177632 228556
rect 177396 170468 177448 170474
rect 177396 170410 177448 170416
rect 177302 27432 177358 27441
rect 177302 27367 177358 27376
rect 177408 27198 177436 170410
rect 177488 166320 177540 166326
rect 177488 166262 177540 166268
rect 177396 27192 177448 27198
rect 177396 27134 177448 27140
rect 177500 26761 177528 166262
rect 177592 159390 177620 228550
rect 177764 192500 177816 192506
rect 177764 192442 177816 192448
rect 177580 159384 177632 159390
rect 177580 159326 177632 159332
rect 177486 26752 177542 26761
rect 177486 26687 177542 26696
rect 177592 24070 177620 159326
rect 177672 147620 177724 147626
rect 177672 147562 177724 147568
rect 177684 64870 177712 147562
rect 177776 140486 177804 192442
rect 178052 172514 178080 233174
rect 178132 213240 178184 213246
rect 178132 213182 178184 213188
rect 178144 212566 178172 213182
rect 178132 212560 178184 212566
rect 178132 212502 178184 212508
rect 178040 172508 178092 172514
rect 178040 172450 178092 172456
rect 177856 171828 177908 171834
rect 177856 171770 177908 171776
rect 177868 144226 177896 171770
rect 178040 146260 178092 146266
rect 178040 146202 178092 146208
rect 178052 144974 178080 146202
rect 178040 144968 178092 144974
rect 178040 144910 178092 144916
rect 177856 144220 177908 144226
rect 177856 144162 177908 144168
rect 177764 140480 177816 140486
rect 177764 140422 177816 140428
rect 177764 127628 177816 127634
rect 177764 127570 177816 127576
rect 177776 106282 177804 127570
rect 177764 106276 177816 106282
rect 177764 106218 177816 106224
rect 177764 89752 177816 89758
rect 177764 89694 177816 89700
rect 177672 64864 177724 64870
rect 177672 64806 177724 64812
rect 177672 57520 177724 57526
rect 177672 57462 177724 57468
rect 177580 24064 177632 24070
rect 177580 24006 177632 24012
rect 177580 10804 177632 10810
rect 177580 10746 177632 10752
rect 177592 3482 177620 10746
rect 177684 3806 177712 57462
rect 177776 28490 177804 89694
rect 178052 63510 178080 144910
rect 178144 141030 178172 212502
rect 178788 209098 178816 355438
rect 178880 233238 178908 453183
rect 178972 383654 179000 582966
rect 180064 581732 180116 581738
rect 180064 581674 180116 581680
rect 179052 562352 179104 562358
rect 179052 562294 179104 562300
rect 179064 419490 179092 562294
rect 179144 474020 179196 474026
rect 179144 473962 179196 473968
rect 179052 419484 179104 419490
rect 179052 419426 179104 419432
rect 178960 383648 179012 383654
rect 178960 383590 179012 383596
rect 179156 361554 179184 473962
rect 179420 453688 179472 453694
rect 179420 453630 179472 453636
rect 179432 452946 179460 453630
rect 179420 452940 179472 452946
rect 179420 452882 179472 452888
rect 179236 450764 179288 450770
rect 179236 450706 179288 450712
rect 179144 361548 179196 361554
rect 179144 361490 179196 361496
rect 178960 348560 179012 348566
rect 178960 348502 179012 348508
rect 178868 233232 178920 233238
rect 178868 233174 178920 233180
rect 178972 232558 179000 348502
rect 179052 348492 179104 348498
rect 179052 348434 179104 348440
rect 179064 313206 179092 348434
rect 179248 345030 179276 450706
rect 179236 345024 179288 345030
rect 179236 344966 179288 344972
rect 179248 344350 179276 344966
rect 179236 344344 179288 344350
rect 179236 344286 179288 344292
rect 179052 313200 179104 313206
rect 179052 313142 179104 313148
rect 179052 264988 179104 264994
rect 179052 264930 179104 264936
rect 179064 253842 179092 264930
rect 179052 253836 179104 253842
rect 179052 253778 179104 253784
rect 179432 246974 179460 452882
rect 180076 387802 180104 581674
rect 180156 472660 180208 472666
rect 180156 472602 180208 472608
rect 180064 387796 180116 387802
rect 180064 387738 180116 387744
rect 180168 362914 180196 472602
rect 180248 471368 180300 471374
rect 180248 471310 180300 471316
rect 180156 362908 180208 362914
rect 180156 362850 180208 362856
rect 180064 354136 180116 354142
rect 180064 354078 180116 354084
rect 179420 246968 179472 246974
rect 179420 246910 179472 246916
rect 179432 245682 179460 246910
rect 179420 245676 179472 245682
rect 179420 245618 179472 245624
rect 179144 244180 179196 244186
rect 179144 244122 179196 244128
rect 179052 233300 179104 233306
rect 179052 233242 179104 233248
rect 178960 232552 179012 232558
rect 178960 232494 179012 232500
rect 178776 209092 178828 209098
rect 178776 209034 178828 209040
rect 178684 185632 178736 185638
rect 178684 185574 178736 185580
rect 178224 176044 178276 176050
rect 178224 175986 178276 175992
rect 178236 147626 178264 175986
rect 178224 147620 178276 147626
rect 178224 147562 178276 147568
rect 178132 141024 178184 141030
rect 178132 140966 178184 140972
rect 178040 63504 178092 63510
rect 178040 63446 178092 63452
rect 178040 54528 178092 54534
rect 178040 54470 178092 54476
rect 177764 28484 177816 28490
rect 177764 28426 177816 28432
rect 178052 16574 178080 54470
rect 178696 28393 178724 185574
rect 178960 170536 179012 170542
rect 178960 170478 179012 170484
rect 178776 169040 178828 169046
rect 178776 168982 178828 168988
rect 178682 28384 178738 28393
rect 178682 28319 178738 28328
rect 178788 27169 178816 168982
rect 178868 164960 178920 164966
rect 178868 164902 178920 164908
rect 178880 27470 178908 164902
rect 178972 142866 179000 170478
rect 179064 151094 179092 233242
rect 179156 185638 179184 244122
rect 179420 213988 179472 213994
rect 179420 213930 179472 213936
rect 179144 185632 179196 185638
rect 179144 185574 179196 185580
rect 179052 151088 179104 151094
rect 179052 151030 179104 151036
rect 178960 142860 179012 142866
rect 178960 142802 179012 142808
rect 179432 138922 179460 213930
rect 180076 206378 180104 354078
rect 180260 353258 180288 471310
rect 180812 427718 180840 584870
rect 181444 579692 181496 579698
rect 181444 579634 181496 579640
rect 181456 444961 181484 579634
rect 181442 444952 181498 444961
rect 181442 444887 181498 444896
rect 180340 427712 180392 427718
rect 180340 427654 180392 427660
rect 180800 427712 180852 427718
rect 180800 427654 180852 427660
rect 180352 363866 180380 427654
rect 181444 419756 181496 419762
rect 181444 419698 181496 419704
rect 180340 363860 180392 363866
rect 180340 363802 180392 363808
rect 180340 362432 180392 362438
rect 180340 362374 180392 362380
rect 180248 353252 180300 353258
rect 180248 353194 180300 353200
rect 180154 352608 180210 352617
rect 180154 352543 180210 352552
rect 180168 229770 180196 352543
rect 180248 347064 180300 347070
rect 180248 347006 180300 347012
rect 180260 320142 180288 347006
rect 180248 320136 180300 320142
rect 180248 320078 180300 320084
rect 180352 300830 180380 362374
rect 180340 300824 180392 300830
rect 180340 300766 180392 300772
rect 180248 289876 180300 289882
rect 180248 289818 180300 289824
rect 180260 252346 180288 289818
rect 180340 273284 180392 273290
rect 180340 273226 180392 273232
rect 180248 252340 180300 252346
rect 180248 252282 180300 252288
rect 180352 250918 180380 273226
rect 180340 250912 180392 250918
rect 180340 250854 180392 250860
rect 180248 245676 180300 245682
rect 180248 245618 180300 245624
rect 180156 229764 180208 229770
rect 180156 229706 180208 229712
rect 180064 206372 180116 206378
rect 180064 206314 180116 206320
rect 180064 186992 180116 186998
rect 180064 186934 180116 186940
rect 179420 138916 179472 138922
rect 179420 138858 179472 138864
rect 178960 134564 179012 134570
rect 178960 134506 179012 134512
rect 178972 109002 179000 134506
rect 178960 108996 179012 109002
rect 178960 108938 179012 108944
rect 178960 93900 179012 93906
rect 178960 93842 179012 93848
rect 178972 28286 179000 93842
rect 179420 46232 179472 46238
rect 179420 46174 179472 46180
rect 178960 28280 179012 28286
rect 178960 28222 179012 28228
rect 178868 27464 178920 27470
rect 178868 27406 178920 27412
rect 178774 27160 178830 27169
rect 178774 27095 178830 27104
rect 179432 16574 179460 46174
rect 180076 22642 180104 186934
rect 180260 173262 180288 245618
rect 180800 244928 180852 244934
rect 180800 244870 180852 244876
rect 180340 231804 180392 231810
rect 180340 231746 180392 231752
rect 180352 186998 180380 231746
rect 180340 186992 180392 186998
rect 180340 186934 180392 186940
rect 180340 177404 180392 177410
rect 180340 177346 180392 177352
rect 180248 173256 180300 173262
rect 180248 173198 180300 173204
rect 180260 161474 180288 173198
rect 180168 161446 180288 161474
rect 180168 27334 180196 161446
rect 180352 149054 180380 177346
rect 180812 174554 180840 244870
rect 180892 227180 180944 227186
rect 180892 227122 180944 227128
rect 180800 174548 180852 174554
rect 180800 174490 180852 174496
rect 180904 171134 180932 227122
rect 180984 209092 181036 209098
rect 180984 209034 181036 209040
rect 180996 206310 181024 209034
rect 180984 206304 181036 206310
rect 180984 206246 181036 206252
rect 180812 171106 180932 171134
rect 180812 161430 180840 171106
rect 180800 161424 180852 161430
rect 180800 161366 180852 161372
rect 180812 160750 180840 161366
rect 180800 160744 180852 160750
rect 180800 160686 180852 160692
rect 180340 149048 180392 149054
rect 180340 148990 180392 148996
rect 180800 147688 180852 147694
rect 180800 147630 180852 147636
rect 180248 133204 180300 133210
rect 180248 133146 180300 133152
rect 180260 110430 180288 133146
rect 180340 123548 180392 123554
rect 180340 123490 180392 123496
rect 180248 110424 180300 110430
rect 180248 110366 180300 110372
rect 180352 100706 180380 123490
rect 180340 100700 180392 100706
rect 180340 100642 180392 100648
rect 180812 66230 180840 147630
rect 181456 137970 181484 419698
rect 181548 380866 181576 585822
rect 182916 572008 182968 572014
rect 182916 571950 182968 571956
rect 181628 570648 181680 570654
rect 181628 570590 181680 570596
rect 181640 405686 181668 570590
rect 181904 475176 181956 475182
rect 181904 475118 181956 475124
rect 181720 474156 181772 474162
rect 181720 474098 181772 474104
rect 181628 405680 181680 405686
rect 181628 405622 181680 405628
rect 181536 380860 181588 380866
rect 181536 380802 181588 380808
rect 181732 340882 181760 474098
rect 181916 460934 181944 475118
rect 181916 460906 182128 460934
rect 181812 457496 181864 457502
rect 181812 457438 181864 457444
rect 181824 361486 181852 457438
rect 182100 449750 182128 460906
rect 182088 449744 182140 449750
rect 182088 449686 182140 449692
rect 181812 361480 181864 361486
rect 181812 361422 181864 361428
rect 181812 356924 181864 356930
rect 181812 356866 181864 356872
rect 181720 340876 181772 340882
rect 181720 340818 181772 340824
rect 181628 340468 181680 340474
rect 181628 340410 181680 340416
rect 181536 340400 181588 340406
rect 181536 340342 181588 340348
rect 181548 202842 181576 340342
rect 181640 224262 181668 340410
rect 181824 303618 181852 356866
rect 181904 351212 181956 351218
rect 181904 351154 181956 351160
rect 181916 321570 181944 351154
rect 181904 321564 181956 321570
rect 181904 321506 181956 321512
rect 181812 303612 181864 303618
rect 181812 303554 181864 303560
rect 181720 281580 181772 281586
rect 181720 281522 181772 281528
rect 181732 252142 181760 281522
rect 181812 266416 181864 266422
rect 181812 266358 181864 266364
rect 181824 253706 181852 266358
rect 181812 253700 181864 253706
rect 181812 253642 181864 253648
rect 181720 252136 181772 252142
rect 181720 252078 181772 252084
rect 182100 234462 182128 449686
rect 182928 413982 182956 571950
rect 183100 471300 183152 471306
rect 183100 471242 183152 471248
rect 183008 460284 183060 460290
rect 183008 460226 183060 460232
rect 182916 413976 182968 413982
rect 182916 413918 182968 413924
rect 182916 349852 182968 349858
rect 182916 349794 182968 349800
rect 182180 347200 182232 347206
rect 182180 347142 182232 347148
rect 182088 234456 182140 234462
rect 182088 234398 182140 234404
rect 181720 232620 181772 232626
rect 181720 232562 181772 232568
rect 181628 224256 181680 224262
rect 181628 224198 181680 224204
rect 181536 202836 181588 202842
rect 181536 202778 181588 202784
rect 181628 195288 181680 195294
rect 181628 195230 181680 195236
rect 181536 187740 181588 187746
rect 181536 187682 181588 187688
rect 181444 137964 181496 137970
rect 181444 137906 181496 137912
rect 181444 130416 181496 130422
rect 181444 130358 181496 130364
rect 181456 108934 181484 130358
rect 181444 108928 181496 108934
rect 181444 108870 181496 108876
rect 180800 66224 180852 66230
rect 180800 66166 180852 66172
rect 181444 57792 181496 57798
rect 181444 57734 181496 57740
rect 180156 27328 180208 27334
rect 180156 27270 180208 27276
rect 180064 22636 180116 22642
rect 180064 22578 180116 22584
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 177672 3800 177724 3806
rect 177672 3742 177724 3748
rect 177592 3454 177896 3482
rect 177868 480 177896 3454
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 180984 10872 181036 10878
rect 180984 10814 181036 10820
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 10814
rect 181456 3602 181484 57734
rect 181548 28257 181576 187682
rect 181640 141302 181668 195230
rect 181732 188358 181760 232562
rect 182192 208350 182220 347142
rect 182928 324290 182956 349794
rect 183020 346322 183048 460226
rect 183112 367062 183140 471242
rect 183468 454912 183520 454918
rect 183468 454854 183520 454860
rect 183480 454238 183508 454854
rect 183192 454232 183244 454238
rect 183192 454174 183244 454180
rect 183468 454232 183520 454238
rect 183468 454174 183520 454180
rect 183100 367056 183152 367062
rect 183100 366998 183152 367004
rect 183008 346316 183060 346322
rect 183008 346258 183060 346264
rect 182916 324284 182968 324290
rect 182916 324226 182968 324232
rect 183008 267776 183060 267782
rect 183008 267718 183060 267724
rect 182916 264240 182968 264246
rect 182916 264182 182968 264188
rect 182928 239426 182956 264182
rect 183020 253638 183048 267718
rect 183008 253632 183060 253638
rect 183008 253574 183060 253580
rect 182916 239420 182968 239426
rect 182916 239362 182968 239368
rect 182824 233912 182876 233918
rect 182824 233854 182876 233860
rect 182180 208344 182232 208350
rect 182180 208286 182232 208292
rect 182836 189786 182864 233854
rect 183204 231810 183232 454174
rect 184216 446418 184244 700402
rect 186964 700392 187016 700398
rect 186964 700334 187016 700340
rect 185676 581664 185728 581670
rect 185676 581606 185728 581612
rect 184296 577584 184348 577590
rect 184296 577526 184348 577532
rect 184204 446412 184256 446418
rect 184204 446354 184256 446360
rect 184204 426488 184256 426494
rect 184204 426430 184256 426436
rect 183560 350056 183612 350062
rect 183560 349998 183612 350004
rect 183008 231804 183060 231810
rect 183008 231746 183060 231752
rect 183192 231804 183244 231810
rect 183192 231746 183244 231752
rect 183020 231130 183048 231746
rect 183008 231124 183060 231130
rect 183008 231066 183060 231072
rect 183572 226302 183600 349998
rect 183652 243568 183704 243574
rect 183652 243510 183704 243516
rect 183560 226296 183612 226302
rect 183560 226238 183612 226244
rect 183572 225622 183600 226238
rect 183560 225616 183612 225622
rect 183560 225558 183612 225564
rect 182916 209228 182968 209234
rect 182916 209170 182968 209176
rect 182824 189780 182876 189786
rect 182824 189722 182876 189728
rect 181720 188352 181772 188358
rect 181720 188294 181772 188300
rect 181732 187746 181760 188294
rect 181720 187740 181772 187746
rect 181720 187682 181772 187688
rect 181720 178696 181772 178702
rect 181720 178638 181772 178644
rect 181732 149122 181760 178638
rect 182088 175228 182140 175234
rect 182088 175170 182140 175176
rect 182100 174554 182128 175170
rect 182088 174548 182140 174554
rect 182088 174490 182140 174496
rect 181720 149116 181772 149122
rect 181720 149058 181772 149064
rect 181904 149048 181956 149054
rect 181904 148990 181956 148996
rect 181916 147694 181944 148990
rect 181904 147688 181956 147694
rect 181904 147630 181956 147636
rect 181628 141296 181680 141302
rect 181628 141238 181680 141244
rect 181534 28248 181590 28257
rect 181534 28183 181590 28192
rect 182836 22098 182864 189722
rect 182928 139262 182956 209170
rect 183664 153882 183692 243510
rect 183744 234456 183796 234462
rect 183744 234398 183796 234404
rect 183756 166326 183784 234398
rect 183744 166320 183796 166326
rect 183744 166262 183796 166268
rect 183652 153876 183704 153882
rect 183652 153818 183704 153824
rect 182916 139256 182968 139262
rect 182916 139198 182968 139204
rect 183560 40724 183612 40730
rect 183560 40666 183612 40672
rect 182824 22092 182876 22098
rect 182824 22034 182876 22040
rect 182180 20460 182232 20466
rect 182180 20402 182232 20408
rect 181444 3596 181496 3602
rect 181444 3538 181496 3544
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 20402
rect 183572 16574 183600 40666
rect 184216 20670 184244 426430
rect 184308 391950 184336 577526
rect 184480 566500 184532 566506
rect 184480 566442 184532 566448
rect 184388 419620 184440 419626
rect 184388 419562 184440 419568
rect 184296 391944 184348 391950
rect 184296 391886 184348 391892
rect 184296 362296 184348 362302
rect 184296 362238 184348 362244
rect 184308 199442 184336 362238
rect 184400 241466 184428 419562
rect 184492 412622 184520 566442
rect 184664 467220 184716 467226
rect 184664 467162 184716 467168
rect 184572 450696 184624 450702
rect 184572 450638 184624 450644
rect 184480 412616 184532 412622
rect 184480 412558 184532 412564
rect 184480 342916 184532 342922
rect 184480 342858 184532 342864
rect 184492 324222 184520 342858
rect 184584 339386 184612 450638
rect 184676 357406 184704 467162
rect 184756 454708 184808 454714
rect 184756 454650 184808 454656
rect 184768 373998 184796 454650
rect 185688 401606 185716 581606
rect 185860 469872 185912 469878
rect 185860 469814 185912 469820
rect 185768 458924 185820 458930
rect 185768 458866 185820 458872
rect 185676 401600 185728 401606
rect 185676 401542 185728 401548
rect 184756 373992 184808 373998
rect 184756 373934 184808 373940
rect 184940 362976 184992 362982
rect 184940 362918 184992 362924
rect 184952 358154 184980 362918
rect 184940 358148 184992 358154
rect 184940 358090 184992 358096
rect 184664 357400 184716 357406
rect 184664 357342 184716 357348
rect 184572 339380 184624 339386
rect 184572 339322 184624 339328
rect 184848 339380 184900 339386
rect 184848 339322 184900 339328
rect 184860 338842 184888 339322
rect 184848 338836 184900 338842
rect 184848 338778 184900 338784
rect 184480 324216 184532 324222
rect 184480 324158 184532 324164
rect 184388 241460 184440 241466
rect 184388 241402 184440 241408
rect 184388 220108 184440 220114
rect 184388 220050 184440 220056
rect 184296 199436 184348 199442
rect 184296 199378 184348 199384
rect 184296 167748 184348 167754
rect 184296 167690 184348 167696
rect 184308 27266 184336 167690
rect 184400 140214 184428 220050
rect 184952 204202 184980 358090
rect 185676 355360 185728 355366
rect 185676 355302 185728 355308
rect 185032 347268 185084 347274
rect 185032 347210 185084 347216
rect 185044 229090 185072 347210
rect 185688 327078 185716 355302
rect 185780 350538 185808 458866
rect 185872 368490 185900 469814
rect 185952 453416 186004 453422
rect 185952 453358 186004 453364
rect 185860 368484 185912 368490
rect 185860 368426 185912 368432
rect 185768 350532 185820 350538
rect 185768 350474 185820 350480
rect 185676 327072 185728 327078
rect 185676 327014 185728 327020
rect 185584 237448 185636 237454
rect 185584 237390 185636 237396
rect 185032 229084 185084 229090
rect 185032 229026 185084 229032
rect 185044 228546 185072 229026
rect 185032 228540 185084 228546
rect 185032 228482 185084 228488
rect 185032 224256 185084 224262
rect 185032 224198 185084 224204
rect 184940 204196 184992 204202
rect 184940 204138 184992 204144
rect 184848 167000 184900 167006
rect 184848 166942 184900 166948
rect 184860 166326 184888 166942
rect 184848 166320 184900 166326
rect 184848 166262 184900 166268
rect 184848 154556 184900 154562
rect 184848 154498 184900 154504
rect 184860 153882 184888 154498
rect 184848 153876 184900 153882
rect 184848 153818 184900 153824
rect 184388 140208 184440 140214
rect 184388 140150 184440 140156
rect 185044 140146 185072 224198
rect 185400 204196 185452 204202
rect 185400 204138 185452 204144
rect 185412 203590 185440 204138
rect 185400 203584 185452 203590
rect 185400 203526 185452 203532
rect 185596 191146 185624 237390
rect 185964 235958 185992 453358
rect 186976 440910 187004 700334
rect 202800 700330 202828 703520
rect 218992 700398 219020 703520
rect 235184 700466 235212 703520
rect 267660 700534 267688 703520
rect 283852 700670 283880 703520
rect 300136 700738 300164 703520
rect 300124 700732 300176 700738
rect 300124 700674 300176 700680
rect 283840 700664 283892 700670
rect 283840 700606 283892 700612
rect 332520 700602 332548 703520
rect 348804 700670 348832 703520
rect 356704 700732 356756 700738
rect 356704 700674 356756 700680
rect 344284 700664 344336 700670
rect 344284 700606 344336 700612
rect 348792 700664 348844 700670
rect 348792 700606 348844 700612
rect 332508 700596 332560 700602
rect 332508 700538 332560 700544
rect 267648 700528 267700 700534
rect 267648 700470 267700 700476
rect 235172 700460 235224 700466
rect 235172 700402 235224 700408
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 188344 700324 188396 700330
rect 188344 700266 188396 700272
rect 202788 700324 202840 700330
rect 202788 700266 202840 700272
rect 187148 584520 187200 584526
rect 187148 584462 187200 584468
rect 187056 539980 187108 539986
rect 187056 539922 187108 539928
rect 187068 487150 187096 539922
rect 187056 487144 187108 487150
rect 187056 487086 187108 487092
rect 187056 452056 187108 452062
rect 187056 451998 187108 452004
rect 187068 451518 187096 451998
rect 187056 451512 187108 451518
rect 187056 451454 187108 451460
rect 186964 440904 187016 440910
rect 186964 440846 187016 440852
rect 186964 438184 187016 438190
rect 186964 438126 187016 438132
rect 186976 360942 187004 438126
rect 186964 360936 187016 360942
rect 186964 360878 187016 360884
rect 186320 344412 186372 344418
rect 186320 344354 186372 344360
rect 185952 235952 186004 235958
rect 185952 235894 186004 235900
rect 185964 235414 185992 235894
rect 185952 235408 186004 235414
rect 185952 235350 186004 235356
rect 186332 212498 186360 344354
rect 186964 344344 187016 344350
rect 186964 344286 187016 344292
rect 186412 249144 186464 249150
rect 186412 249086 186464 249092
rect 186320 212492 186372 212498
rect 186320 212434 186372 212440
rect 186332 211818 186360 212434
rect 186320 211812 186372 211818
rect 186320 211754 186372 211760
rect 186320 204944 186372 204950
rect 186320 204886 186372 204892
rect 186332 204338 186360 204886
rect 186320 204332 186372 204338
rect 186320 204274 186372 204280
rect 185584 191140 185636 191146
rect 185584 191082 185636 191088
rect 185032 140140 185084 140146
rect 185032 140082 185084 140088
rect 184388 126268 184440 126274
rect 184388 126210 184440 126216
rect 184400 111790 184428 126210
rect 184388 111784 184440 111790
rect 184388 111726 184440 111732
rect 184940 51740 184992 51746
rect 184940 51682 184992 51688
rect 184296 27260 184348 27266
rect 184296 27202 184348 27208
rect 184204 20664 184256 20670
rect 184204 20606 184256 20612
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 480 184980 51682
rect 185596 23458 185624 191082
rect 186424 161474 186452 249086
rect 186504 204332 186556 204338
rect 186504 204274 186556 204280
rect 186332 161446 186452 161474
rect 186332 153202 186360 161446
rect 186320 153196 186372 153202
rect 186320 153138 186372 153144
rect 186332 152522 186360 153138
rect 186320 152516 186372 152522
rect 186320 152458 186372 152464
rect 186320 142860 186372 142866
rect 186320 142802 186372 142808
rect 186332 142186 186360 142802
rect 186320 142180 186372 142186
rect 186320 142122 186372 142128
rect 186332 59362 186360 142122
rect 186516 138854 186544 204274
rect 186976 191894 187004 344286
rect 187068 227730 187096 451454
rect 187160 394670 187188 584462
rect 187700 475108 187752 475114
rect 187700 475050 187752 475056
rect 187712 474881 187740 475050
rect 187698 474872 187754 474881
rect 187698 474807 187754 474816
rect 187240 468580 187292 468586
rect 187240 468522 187292 468528
rect 187148 394664 187200 394670
rect 187148 394606 187200 394612
rect 187252 356046 187280 468522
rect 187424 464364 187476 464370
rect 187424 464306 187476 464312
rect 187332 450832 187384 450838
rect 187332 450774 187384 450780
rect 187240 356040 187292 356046
rect 187240 355982 187292 355988
rect 187148 355428 187200 355434
rect 187148 355370 187200 355376
rect 187160 306338 187188 355370
rect 187344 342242 187372 450774
rect 187436 375358 187464 464306
rect 187516 419552 187568 419558
rect 187516 419494 187568 419500
rect 187424 375352 187476 375358
rect 187424 375294 187476 375300
rect 187528 346390 187556 419494
rect 187516 346384 187568 346390
rect 187516 346326 187568 346332
rect 187332 342236 187384 342242
rect 187332 342178 187384 342184
rect 187344 340950 187372 342178
rect 187332 340944 187384 340950
rect 187332 340886 187384 340892
rect 187240 338972 187292 338978
rect 187240 338914 187292 338920
rect 187252 329798 187280 338914
rect 187240 329792 187292 329798
rect 187240 329734 187292 329740
rect 187148 306332 187200 306338
rect 187148 306274 187200 306280
rect 187148 270564 187200 270570
rect 187148 270506 187200 270512
rect 187160 253570 187188 270506
rect 187240 260908 187292 260914
rect 187240 260850 187292 260856
rect 187148 253564 187200 253570
rect 187148 253506 187200 253512
rect 187252 250714 187280 260850
rect 187240 250708 187292 250714
rect 187240 250650 187292 250656
rect 187712 238678 187740 474807
rect 187792 439680 187844 439686
rect 187792 439622 187844 439628
rect 187804 438870 187832 439622
rect 188356 439550 188384 700266
rect 340144 660340 340196 660346
rect 340144 660282 340196 660288
rect 246304 659728 246356 659734
rect 246302 659696 246304 659705
rect 337108 659728 337160 659734
rect 246356 659696 246358 659705
rect 340156 659705 340184 660282
rect 337108 659670 337160 659676
rect 340142 659696 340198 659705
rect 246302 659631 246358 659640
rect 237286 654528 237342 654537
rect 237286 654463 237342 654472
rect 237194 591696 237250 591705
rect 237194 591631 237250 591640
rect 196900 584452 196952 584458
rect 196900 584394 196952 584400
rect 189816 580304 189868 580310
rect 189816 580246 189868 580252
rect 188436 574864 188488 574870
rect 188436 574806 188488 574812
rect 188344 439544 188396 439550
rect 188344 439486 188396 439492
rect 187792 438864 187844 438870
rect 187792 438806 187844 438812
rect 187804 362982 187832 438806
rect 188448 390522 188476 574806
rect 188528 565208 188580 565214
rect 188528 565150 188580 565156
rect 188540 411262 188568 565150
rect 188620 461712 188672 461718
rect 188620 461654 188672 461660
rect 188528 411256 188580 411262
rect 188528 411198 188580 411204
rect 188436 390516 188488 390522
rect 188436 390458 188488 390464
rect 187792 362976 187844 362982
rect 187792 362918 187844 362924
rect 188632 358698 188660 461654
rect 188712 456068 188764 456074
rect 188712 456010 188764 456016
rect 188724 378146 188752 456010
rect 189724 453348 189776 453354
rect 189724 453290 189776 453296
rect 188712 378140 188764 378146
rect 188712 378082 188764 378088
rect 188620 358692 188672 358698
rect 188620 358634 188672 358640
rect 187884 358080 187936 358086
rect 187884 358022 187936 358028
rect 187792 340944 187844 340950
rect 187792 340886 187844 340892
rect 187700 238672 187752 238678
rect 187700 238614 187752 238620
rect 187148 227792 187200 227798
rect 187148 227734 187200 227740
rect 187056 227724 187108 227730
rect 187056 227666 187108 227672
rect 187068 226370 187096 227666
rect 187056 226364 187108 226370
rect 187056 226306 187108 226312
rect 186964 191888 187016 191894
rect 186964 191830 187016 191836
rect 187160 162178 187188 227734
rect 187712 169726 187740 238614
rect 187804 194546 187832 340886
rect 187896 223582 187924 358022
rect 189172 356788 189224 356794
rect 189172 356730 189224 356736
rect 188344 348424 188396 348430
rect 188344 348366 188396 348372
rect 188356 331226 188384 348366
rect 189080 345772 189132 345778
rect 189080 345714 189132 345720
rect 188344 331220 188396 331226
rect 188344 331162 188396 331168
rect 188436 235340 188488 235346
rect 188436 235282 188488 235288
rect 187884 223576 187936 223582
rect 187884 223518 187936 223524
rect 187896 222902 187924 223518
rect 187884 222896 187936 222902
rect 187884 222838 187936 222844
rect 187884 202836 187936 202842
rect 187884 202778 187936 202784
rect 187896 201550 187924 202778
rect 187884 201544 187936 201550
rect 187884 201486 187936 201492
rect 187792 194540 187844 194546
rect 187792 194482 187844 194488
rect 187804 193866 187832 194482
rect 187792 193860 187844 193866
rect 187792 193802 187844 193808
rect 187700 169720 187752 169726
rect 187700 169662 187752 169668
rect 187712 169046 187740 169662
rect 187700 169040 187752 169046
rect 187700 168982 187752 168988
rect 187148 162172 187200 162178
rect 187148 162114 187200 162120
rect 187160 161474 187188 162114
rect 186976 161446 187188 161474
rect 186504 138848 186556 138854
rect 186504 138790 186556 138796
rect 186320 59356 186372 59362
rect 186320 59298 186372 59304
rect 186320 39364 186372 39370
rect 186320 39306 186372 39312
rect 185584 23452 185636 23458
rect 185584 23394 185636 23400
rect 185032 21684 185084 21690
rect 185032 21626 185084 21632
rect 185044 16574 185072 21626
rect 186332 16574 186360 39306
rect 186976 28966 187004 161446
rect 187700 149116 187752 149122
rect 187700 149058 187752 149064
rect 187712 69698 187740 149058
rect 187896 141098 187924 201486
rect 188344 164212 188396 164218
rect 188344 164154 188396 164160
rect 187884 141092 187936 141098
rect 187884 141034 187936 141040
rect 187700 69692 187752 69698
rect 187700 69634 187752 69640
rect 186964 28960 187016 28966
rect 188356 28937 188384 164154
rect 188448 156670 188476 235282
rect 189092 197334 189120 345714
rect 189184 218006 189212 356730
rect 189264 252408 189316 252414
rect 189264 252350 189316 252356
rect 189276 251870 189304 252350
rect 189264 251864 189316 251870
rect 189264 251806 189316 251812
rect 189736 242826 189764 453290
rect 189828 416770 189856 580246
rect 191196 579012 191248 579018
rect 191196 578954 191248 578960
rect 190368 539912 190420 539918
rect 190368 539854 190420 539860
rect 189908 471436 189960 471442
rect 189908 471378 189960 471384
rect 189816 416764 189868 416770
rect 189816 416706 189868 416712
rect 189920 345030 189948 471378
rect 190000 461644 190052 461650
rect 190000 461586 190052 461592
rect 190012 369850 190040 461586
rect 190000 369844 190052 369850
rect 190000 369786 190052 369792
rect 189908 345024 189960 345030
rect 189908 344966 189960 344972
rect 190380 252414 190408 539854
rect 191104 453552 191156 453558
rect 191104 453494 191156 453500
rect 190460 426352 190512 426358
rect 190460 426294 190512 426300
rect 190472 363662 190500 426294
rect 190460 363656 190512 363662
rect 190460 363598 190512 363604
rect 190460 349988 190512 349994
rect 190460 349930 190512 349936
rect 190368 252408 190420 252414
rect 190368 252350 190420 252356
rect 189724 242820 189776 242826
rect 189724 242762 189776 242768
rect 190000 242820 190052 242826
rect 190000 242762 190052 242768
rect 190012 242214 190040 242762
rect 190000 242208 190052 242214
rect 190000 242150 190052 242156
rect 189264 236768 189316 236774
rect 189264 236710 189316 236716
rect 189172 218000 189224 218006
rect 189172 217942 189224 217948
rect 189184 217326 189212 217942
rect 189172 217320 189224 217326
rect 189172 217262 189224 217268
rect 189080 197328 189132 197334
rect 189080 197270 189132 197276
rect 189092 196654 189120 197270
rect 189080 196648 189132 196654
rect 189080 196590 189132 196596
rect 188436 156664 188488 156670
rect 188436 156606 188488 156612
rect 188448 29034 188476 156606
rect 189276 155922 189304 236710
rect 189356 226364 189408 226370
rect 189356 226306 189408 226312
rect 189368 164218 189396 226306
rect 190472 198014 190500 349930
rect 191116 248334 191144 453494
rect 191208 389162 191236 578954
rect 194048 578944 194100 578950
rect 194048 578886 194100 578892
rect 191288 574796 191340 574802
rect 191288 574738 191340 574744
rect 191300 409766 191328 574738
rect 191748 573436 191800 573442
rect 191748 573378 191800 573384
rect 191656 569356 191708 569362
rect 191656 569298 191708 569304
rect 191380 472728 191432 472734
rect 191380 472670 191432 472676
rect 191288 409760 191340 409766
rect 191288 409702 191340 409708
rect 191196 389156 191248 389162
rect 191196 389098 191248 389104
rect 191196 354204 191248 354210
rect 191196 354146 191248 354152
rect 191104 248328 191156 248334
rect 191104 248270 191156 248276
rect 191116 247110 191144 248270
rect 191104 247104 191156 247110
rect 191104 247046 191156 247052
rect 191104 240780 191156 240786
rect 191104 240722 191156 240728
rect 190460 198008 190512 198014
rect 190460 197950 190512 197956
rect 190460 191888 190512 191894
rect 190460 191830 190512 191836
rect 189356 164212 189408 164218
rect 189356 164154 189408 164160
rect 189080 155916 189132 155922
rect 189080 155858 189132 155864
rect 189264 155916 189316 155922
rect 189264 155858 189316 155864
rect 189092 155310 189120 155858
rect 189080 155304 189132 155310
rect 189080 155246 189132 155252
rect 190472 141166 190500 191830
rect 191116 175710 191144 240722
rect 191208 229022 191236 354146
rect 191392 343602 191420 472670
rect 191472 469940 191524 469946
rect 191472 469882 191524 469888
rect 191484 354414 191512 469882
rect 191564 462392 191616 462398
rect 191564 462334 191616 462340
rect 191576 434110 191604 462334
rect 191668 445058 191696 569298
rect 191656 445052 191708 445058
rect 191656 444994 191708 445000
rect 191760 442406 191788 573378
rect 193036 572484 193088 572490
rect 193036 572426 193088 572432
rect 192944 572280 192996 572286
rect 192944 572222 192996 572228
rect 192760 572076 192812 572082
rect 192760 572018 192812 572024
rect 192484 569220 192536 569226
rect 192484 569162 192536 569168
rect 191748 442400 191800 442406
rect 191748 442342 191800 442348
rect 191564 434104 191616 434110
rect 191564 434046 191616 434052
rect 191748 427100 191800 427106
rect 191748 427042 191800 427048
rect 191760 426358 191788 427042
rect 191748 426352 191800 426358
rect 191748 426294 191800 426300
rect 192496 404326 192524 569162
rect 192576 474088 192628 474094
rect 192576 474030 192628 474036
rect 192484 404320 192536 404326
rect 192484 404262 192536 404268
rect 191840 356856 191892 356862
rect 191840 356798 191892 356804
rect 191472 354408 191524 354414
rect 191472 354350 191524 354356
rect 191380 343596 191432 343602
rect 191380 343538 191432 343544
rect 191196 229016 191248 229022
rect 191196 228958 191248 228964
rect 191288 202836 191340 202842
rect 191288 202778 191340 202784
rect 191104 175704 191156 175710
rect 191104 175646 191156 175652
rect 190460 141160 190512 141166
rect 190460 141102 190512 141108
rect 188528 57384 188580 57390
rect 188528 57326 188580 57332
rect 188436 29028 188488 29034
rect 188436 28970 188488 28976
rect 186964 28902 187016 28908
rect 188342 28928 188398 28937
rect 188342 28863 188398 28872
rect 188540 16574 188568 57326
rect 190460 35216 190512 35222
rect 190460 35158 190512 35164
rect 189080 31136 189132 31142
rect 189080 31078 189132 31084
rect 189092 16574 189120 31078
rect 185044 16546 186176 16574
rect 186332 16546 186912 16574
rect 188540 16546 188660 16574
rect 189092 16546 189304 16574
rect 186148 480 186176 16546
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188528 10940 188580 10946
rect 188528 10882 188580 10888
rect 188540 480 188568 10882
rect 188632 3942 188660 16546
rect 188620 3936 188672 3942
rect 188620 3878 188672 3884
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 35158
rect 191116 22030 191144 175646
rect 191196 144764 191248 144770
rect 191196 144706 191248 144712
rect 191208 64190 191236 144706
rect 191300 139398 191328 202778
rect 191852 200802 191880 356798
rect 192482 342952 192538 342961
rect 192482 342887 192538 342896
rect 192024 249076 192076 249082
rect 192024 249018 192076 249024
rect 191932 228472 191984 228478
rect 191932 228414 191984 228420
rect 191840 200796 191892 200802
rect 191840 200738 191892 200744
rect 191944 140078 191972 228414
rect 192036 182850 192064 249018
rect 192496 227730 192524 342887
rect 192588 342242 192616 474030
rect 192668 468648 192720 468654
rect 192668 468590 192720 468596
rect 192680 349042 192708 468590
rect 192772 447710 192800 572018
rect 192852 569288 192904 569294
rect 192852 569230 192904 569236
rect 192760 447704 192812 447710
rect 192760 447646 192812 447652
rect 192864 445194 192892 569230
rect 192852 445188 192904 445194
rect 192852 445130 192904 445136
rect 192956 445097 192984 572222
rect 192942 445088 192998 445097
rect 192942 445023 192998 445032
rect 193048 444922 193076 572426
rect 193128 572144 193180 572150
rect 193128 572086 193180 572092
rect 193140 445369 193168 572086
rect 193956 570716 194008 570722
rect 193956 570658 194008 570664
rect 193864 474904 193916 474910
rect 193864 474846 193916 474852
rect 193772 468512 193824 468518
rect 193772 468454 193824 468460
rect 193588 454028 193640 454034
rect 193588 453970 193640 453976
rect 193600 453218 193628 453970
rect 193588 453212 193640 453218
rect 193588 453154 193640 453160
rect 193126 445360 193182 445369
rect 193126 445295 193182 445304
rect 193036 444916 193088 444922
rect 193036 444858 193088 444864
rect 193220 360936 193272 360942
rect 193220 360878 193272 360884
rect 192668 349036 192720 349042
rect 192668 348978 192720 348984
rect 192576 342236 192628 342242
rect 192576 342178 192628 342184
rect 192484 227724 192536 227730
rect 192484 227666 192536 227672
rect 193232 192506 193260 360878
rect 193600 249762 193628 453154
rect 193680 450900 193732 450906
rect 193680 450842 193732 450848
rect 193692 360194 193720 450842
rect 193784 372502 193812 468454
rect 193876 454034 193904 474846
rect 193864 454028 193916 454034
rect 193864 453970 193916 453976
rect 193864 421660 193916 421666
rect 193864 421602 193916 421608
rect 193772 372496 193824 372502
rect 193772 372438 193824 372444
rect 193680 360188 193732 360194
rect 193680 360130 193732 360136
rect 193588 249756 193640 249762
rect 193588 249698 193640 249704
rect 193600 249218 193628 249698
rect 193588 249212 193640 249218
rect 193588 249154 193640 249160
rect 193404 247104 193456 247110
rect 193404 247046 193456 247052
rect 193312 199436 193364 199442
rect 193312 199378 193364 199384
rect 193220 192500 193272 192506
rect 193220 192442 193272 192448
rect 192024 182844 192076 182850
rect 192024 182786 192076 182792
rect 193324 140962 193352 199378
rect 193416 164966 193444 247046
rect 193496 220856 193548 220862
rect 193496 220798 193548 220804
rect 193508 218754 193536 220798
rect 193496 218748 193548 218754
rect 193496 218690 193548 218696
rect 193404 164960 193456 164966
rect 193404 164902 193456 164908
rect 193312 140956 193364 140962
rect 193312 140898 193364 140904
rect 191932 140072 191984 140078
rect 191932 140014 191984 140020
rect 191288 139392 191340 139398
rect 191288 139334 191340 139340
rect 193876 115326 193904 421602
rect 193968 386306 193996 570658
rect 194060 408474 194088 578886
rect 195428 577516 195480 577522
rect 195428 577458 195480 577464
rect 194416 572416 194468 572422
rect 194416 572358 194468 572364
rect 194324 572348 194376 572354
rect 194324 572290 194376 572296
rect 194140 572008 194192 572014
rect 194140 571950 194192 571956
rect 194152 450974 194180 571950
rect 194232 569424 194284 569430
rect 194232 569366 194284 569372
rect 194140 450968 194192 450974
rect 194140 450910 194192 450916
rect 194244 445126 194272 569366
rect 194336 445233 194364 572290
rect 194322 445224 194378 445233
rect 194322 445159 194378 445168
rect 194232 445120 194284 445126
rect 194232 445062 194284 445068
rect 194428 444854 194456 572358
rect 194508 572212 194560 572218
rect 194508 572154 194560 572160
rect 194520 447642 194548 572154
rect 195336 569492 195388 569498
rect 195336 569434 195388 569440
rect 195244 472048 195296 472054
rect 195244 471990 195296 471996
rect 195152 467152 195204 467158
rect 195152 467094 195204 467100
rect 195060 457768 195112 457774
rect 195060 457710 195112 457716
rect 195072 451654 195100 457710
rect 195060 451648 195112 451654
rect 195060 451590 195112 451596
rect 194508 447636 194560 447642
rect 194508 447578 194560 447584
rect 194416 444848 194468 444854
rect 194416 444790 194468 444796
rect 194048 408468 194100 408474
rect 194048 408410 194100 408416
rect 193956 386300 194008 386306
rect 193956 386242 194008 386248
rect 195164 371210 195192 467094
rect 195256 457638 195284 471990
rect 195244 457632 195296 457638
rect 195244 457574 195296 457580
rect 195244 455524 195296 455530
rect 195244 455466 195296 455472
rect 195256 452402 195284 455466
rect 195244 452396 195296 452402
rect 195244 452338 195296 452344
rect 195244 421524 195296 421530
rect 195244 421466 195296 421472
rect 195152 371204 195204 371210
rect 195152 371146 195204 371152
rect 194600 360188 194652 360194
rect 194600 360130 194652 360136
rect 193956 227112 194008 227118
rect 193956 227054 194008 227060
rect 193968 158370 193996 227054
rect 194612 195974 194640 360130
rect 194876 340264 194928 340270
rect 194876 340206 194928 340212
rect 194888 336666 194916 340206
rect 194876 336660 194928 336666
rect 194876 336602 194928 336608
rect 194692 249212 194744 249218
rect 194692 249154 194744 249160
rect 194600 195968 194652 195974
rect 194600 195910 194652 195916
rect 194612 195294 194640 195910
rect 194600 195288 194652 195294
rect 194600 195230 194652 195236
rect 194600 173188 194652 173194
rect 194600 173130 194652 173136
rect 193956 158364 194008 158370
rect 193956 158306 194008 158312
rect 193864 115320 193916 115326
rect 193864 115262 193916 115268
rect 191196 64184 191248 64190
rect 191196 64126 191248 64132
rect 191840 44940 191892 44946
rect 191840 44882 191892 44888
rect 191104 22024 191156 22030
rect 191104 21966 191156 21972
rect 191852 16574 191880 44882
rect 193220 43444 193272 43450
rect 193220 43386 193272 43392
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 3602 193260 43386
rect 193312 26920 193364 26926
rect 193312 26862 193364 26868
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 193324 3482 193352 26862
rect 193968 24857 193996 158306
rect 194612 144770 194640 173130
rect 194704 168366 194732 249154
rect 195256 228410 195284 421466
rect 195348 386374 195376 569434
rect 195440 407114 195468 577458
rect 196808 576156 196860 576162
rect 196808 576098 196860 576104
rect 195704 575136 195756 575142
rect 195704 575078 195756 575084
rect 195612 574728 195664 574734
rect 195612 574670 195664 574676
rect 195520 574116 195572 574122
rect 195520 574058 195572 574064
rect 195532 457774 195560 574058
rect 195520 457768 195572 457774
rect 195520 457710 195572 457716
rect 195520 457632 195572 457638
rect 195520 457574 195572 457580
rect 195532 452538 195560 457574
rect 195520 452532 195572 452538
rect 195520 452474 195572 452480
rect 195624 447846 195652 574670
rect 195716 448050 195744 575078
rect 195888 574932 195940 574938
rect 195888 574874 195940 574880
rect 195796 574592 195848 574598
rect 195796 574534 195848 574540
rect 195704 448044 195756 448050
rect 195704 447986 195756 447992
rect 195808 447982 195836 574534
rect 195796 447976 195848 447982
rect 195796 447918 195848 447924
rect 195612 447840 195664 447846
rect 195612 447782 195664 447788
rect 195900 445602 195928 574874
rect 196716 574252 196768 574258
rect 196716 574194 196768 574200
rect 196624 572552 196676 572558
rect 196624 572494 196676 572500
rect 196072 455456 196124 455462
rect 196072 455398 196124 455404
rect 195980 454096 196032 454102
rect 195980 454038 196032 454044
rect 195992 452266 196020 454038
rect 196084 452334 196112 455398
rect 196164 453416 196216 453422
rect 196164 453358 196216 453364
rect 196176 453257 196204 453358
rect 196162 453248 196218 453257
rect 196162 453183 196218 453192
rect 196072 452328 196124 452334
rect 196072 452270 196124 452276
rect 195980 452260 196032 452266
rect 195980 452202 196032 452208
rect 195888 445596 195940 445602
rect 195888 445538 195940 445544
rect 196636 445398 196664 572494
rect 196728 448118 196756 574194
rect 196716 448112 196768 448118
rect 196716 448054 196768 448060
rect 196624 445392 196676 445398
rect 196624 445334 196676 445340
rect 196624 421728 196676 421734
rect 196624 421670 196676 421676
rect 195520 419688 195572 419694
rect 195520 419630 195572 419636
rect 195428 407108 195480 407114
rect 195428 407050 195480 407056
rect 195336 386368 195388 386374
rect 195336 386310 195388 386316
rect 195532 358766 195560 419630
rect 195520 358760 195572 358766
rect 195520 358702 195572 358708
rect 195428 354068 195480 354074
rect 195428 354010 195480 354016
rect 195336 351280 195388 351286
rect 195336 351222 195388 351228
rect 195244 228404 195296 228410
rect 195244 228346 195296 228352
rect 195348 218822 195376 351222
rect 195440 307766 195468 354010
rect 195428 307760 195480 307766
rect 195428 307702 195480 307708
rect 195428 261520 195480 261526
rect 195428 261462 195480 261468
rect 195440 235958 195468 261462
rect 195980 239420 196032 239426
rect 195980 239362 196032 239368
rect 195992 238950 196020 239362
rect 195980 238944 196032 238950
rect 195980 238886 196032 238892
rect 195428 235952 195480 235958
rect 195428 235894 195480 235900
rect 195428 235408 195480 235414
rect 195428 235350 195480 235356
rect 195336 218816 195388 218822
rect 195336 218758 195388 218764
rect 195440 180794 195468 235350
rect 195256 180766 195468 180794
rect 195256 179518 195284 180766
rect 195244 179512 195296 179518
rect 195244 179454 195296 179460
rect 194692 168360 194744 168366
rect 194692 168302 194744 168308
rect 194704 167754 194732 168302
rect 194692 167748 194744 167754
rect 194692 167690 194744 167696
rect 194600 144764 194652 144770
rect 194600 144706 194652 144712
rect 194600 144220 194652 144226
rect 194600 144162 194652 144168
rect 194612 143614 194640 144162
rect 194600 143608 194652 143614
rect 194600 143550 194652 143556
rect 194048 135924 194100 135930
rect 194048 135866 194100 135872
rect 194060 102134 194088 135866
rect 194048 102128 194100 102134
rect 194048 102070 194100 102076
rect 194612 61402 194640 143550
rect 194600 61396 194652 61402
rect 194600 61338 194652 61344
rect 194600 42152 194652 42158
rect 194600 42094 194652 42100
rect 193954 24848 194010 24857
rect 193954 24783 194010 24792
rect 194612 16574 194640 42094
rect 195256 22710 195284 179454
rect 195992 164898 196020 238886
rect 196072 206372 196124 206378
rect 196072 206314 196124 206320
rect 195980 164892 196032 164898
rect 195980 164834 196032 164840
rect 196084 139330 196112 206314
rect 196072 139324 196124 139330
rect 196072 139266 196124 139272
rect 196636 113830 196664 421670
rect 196714 421424 196770 421433
rect 196714 421359 196770 421368
rect 196728 115258 196756 421359
rect 196820 402393 196848 576098
rect 196912 417217 196940 584394
rect 199384 575204 199436 575210
rect 199384 575146 199436 575152
rect 198648 575068 198700 575074
rect 198648 575010 198700 575016
rect 197084 574864 197136 574870
rect 197084 574806 197136 574812
rect 196992 574184 197044 574190
rect 196992 574126 197044 574132
rect 197004 447914 197032 574126
rect 197096 456210 197124 574806
rect 197176 574796 197228 574802
rect 197176 574738 197228 574744
rect 197084 456204 197136 456210
rect 197084 456146 197136 456152
rect 197188 456090 197216 574738
rect 198370 574696 198426 574705
rect 198370 574631 198426 574640
rect 197358 533216 197414 533225
rect 197096 456062 197216 456090
rect 197280 533174 197358 533202
rect 196992 447908 197044 447914
rect 196992 447850 197044 447856
rect 197096 444990 197124 456062
rect 197176 456000 197228 456006
rect 197176 455942 197228 455948
rect 197188 445670 197216 455942
rect 197176 445664 197228 445670
rect 197176 445606 197228 445612
rect 197084 444984 197136 444990
rect 197084 444926 197136 444932
rect 196992 421456 197044 421462
rect 196992 421398 197044 421404
rect 196898 417208 196954 417217
rect 196898 417143 196954 417152
rect 196806 402384 196862 402393
rect 196806 402319 196862 402328
rect 196808 338836 196860 338842
rect 196808 338778 196860 338784
rect 196820 215422 196848 338778
rect 197004 338774 197032 421398
rect 197084 421388 197136 421394
rect 197084 421330 197136 421336
rect 197096 340202 197124 421330
rect 197176 421320 197228 421326
rect 197176 421262 197228 421268
rect 197188 365702 197216 421262
rect 197176 365696 197228 365702
rect 197176 365638 197228 365644
rect 197084 340196 197136 340202
rect 197084 340138 197136 340144
rect 196992 338768 197044 338774
rect 196992 338710 197044 338716
rect 197280 248849 197308 533174
rect 197358 533151 197414 533160
rect 198278 473376 198334 473385
rect 198278 473311 198334 473320
rect 198186 471744 198242 471753
rect 198186 471679 198242 471688
rect 198094 470384 198150 470393
rect 198094 470319 198150 470328
rect 198002 468888 198058 468897
rect 198002 468823 198058 468832
rect 197818 467664 197874 467673
rect 197818 467599 197874 467608
rect 197832 460934 197860 467599
rect 197832 460906 197952 460934
rect 197360 454232 197412 454238
rect 197360 454174 197412 454180
rect 197372 452470 197400 454174
rect 197360 452464 197412 452470
rect 197360 452406 197412 452412
rect 197924 448526 197952 460906
rect 197912 448520 197964 448526
rect 198016 448497 198044 468823
rect 197912 448462 197964 448468
rect 198002 448488 198058 448497
rect 197818 421696 197874 421705
rect 197818 421631 197874 421640
rect 197360 419484 197412 419490
rect 197360 419426 197412 419432
rect 197372 419121 197400 419426
rect 197358 419112 197414 419121
rect 197358 419047 197414 419056
rect 197360 416764 197412 416770
rect 197360 416706 197412 416712
rect 197372 416673 197400 416706
rect 197358 416664 197414 416673
rect 197358 416599 197414 416608
rect 197360 415404 197412 415410
rect 197360 415346 197412 415352
rect 197372 415041 197400 415346
rect 197358 415032 197414 415041
rect 197358 414967 197414 414976
rect 197360 413976 197412 413982
rect 197360 413918 197412 413924
rect 197372 413545 197400 413918
rect 197358 413536 197414 413545
rect 197358 413471 197414 413480
rect 197360 412616 197412 412622
rect 197360 412558 197412 412564
rect 197372 412321 197400 412558
rect 197358 412312 197414 412321
rect 197358 412247 197414 412256
rect 197360 411256 197412 411262
rect 197360 411198 197412 411204
rect 197372 411097 197400 411198
rect 197358 411088 197414 411097
rect 197358 411023 197414 411032
rect 197358 409864 197414 409873
rect 197358 409799 197360 409808
rect 197412 409799 197414 409808
rect 197360 409770 197412 409776
rect 197452 409760 197504 409766
rect 197452 409702 197504 409708
rect 197464 408649 197492 409702
rect 197450 408640 197506 408649
rect 197450 408575 197506 408584
rect 197360 408468 197412 408474
rect 197360 408410 197412 408416
rect 197372 407969 197400 408410
rect 197358 407960 197414 407969
rect 197358 407895 197414 407904
rect 197728 407108 197780 407114
rect 197728 407050 197780 407056
rect 197740 406065 197768 407050
rect 197726 406056 197782 406065
rect 197726 405991 197782 406000
rect 197360 405680 197412 405686
rect 197360 405622 197412 405628
rect 197372 404841 197400 405622
rect 197358 404832 197414 404841
rect 197358 404767 197414 404776
rect 197360 404320 197412 404326
rect 197360 404262 197412 404268
rect 197372 403617 197400 404262
rect 197358 403608 197414 403617
rect 197358 403543 197414 403552
rect 197360 401600 197412 401606
rect 197360 401542 197412 401548
rect 197372 401169 197400 401542
rect 197358 401160 197414 401169
rect 197358 401095 197414 401104
rect 197360 400172 197412 400178
rect 197360 400114 197412 400120
rect 197372 399945 197400 400114
rect 197358 399936 197414 399945
rect 197358 399871 197414 399880
rect 197360 398812 197412 398818
rect 197360 398754 197412 398760
rect 197372 398721 197400 398754
rect 197452 398744 197504 398750
rect 197358 398712 197414 398721
rect 197452 398686 197504 398692
rect 197358 398647 197414 398656
rect 197464 397497 197492 398686
rect 197450 397488 197506 397497
rect 197360 397452 197412 397458
rect 197450 397423 197506 397432
rect 197360 397394 197412 397400
rect 197372 396137 197400 397394
rect 197358 396128 197414 396137
rect 197358 396063 197414 396072
rect 197360 396024 197412 396030
rect 197360 395966 197412 395972
rect 197372 394913 197400 395966
rect 197358 394904 197414 394913
rect 197358 394839 197414 394848
rect 197360 394664 197412 394670
rect 197360 394606 197412 394612
rect 197372 393689 197400 394606
rect 197358 393680 197414 393689
rect 197358 393615 197414 393624
rect 197360 393304 197412 393310
rect 197360 393246 197412 393252
rect 197372 392465 197400 393246
rect 197358 392456 197414 392465
rect 197358 392391 197414 392400
rect 197360 391944 197412 391950
rect 197360 391886 197412 391892
rect 197372 391241 197400 391886
rect 197358 391232 197414 391241
rect 197358 391167 197414 391176
rect 197360 390516 197412 390522
rect 197360 390458 197412 390464
rect 197372 390017 197400 390458
rect 197358 390008 197414 390017
rect 197358 389943 197414 389952
rect 197360 389156 197412 389162
rect 197360 389098 197412 389104
rect 197372 388793 197400 389098
rect 197358 388784 197414 388793
rect 197358 388719 197414 388728
rect 197360 387796 197412 387802
rect 197360 387738 197412 387744
rect 197372 387569 197400 387738
rect 197358 387560 197414 387569
rect 197358 387495 197414 387504
rect 197728 386368 197780 386374
rect 197358 386336 197414 386345
rect 197728 386310 197780 386316
rect 197358 386271 197360 386280
rect 197412 386271 197414 386280
rect 197360 386242 197412 386248
rect 197740 385121 197768 386310
rect 197726 385112 197782 385121
rect 197726 385047 197782 385056
rect 197360 385008 197412 385014
rect 197360 384950 197412 384956
rect 197372 384441 197400 384950
rect 197358 384432 197414 384441
rect 197358 384367 197414 384376
rect 197360 383648 197412 383654
rect 197360 383590 197412 383596
rect 197372 383217 197400 383590
rect 197358 383208 197414 383217
rect 197358 383143 197414 383152
rect 197360 382220 197412 382226
rect 197360 382162 197412 382168
rect 197372 381313 197400 382162
rect 197358 381304 197414 381313
rect 197358 381239 197414 381248
rect 197360 380860 197412 380866
rect 197360 380802 197412 380808
rect 197372 380089 197400 380802
rect 197358 380080 197414 380089
rect 197358 380015 197414 380024
rect 197360 379500 197412 379506
rect 197360 379442 197412 379448
rect 197372 378865 197400 379442
rect 197358 378856 197414 378865
rect 197358 378791 197414 378800
rect 197360 378140 197412 378146
rect 197360 378082 197412 378088
rect 197372 377641 197400 378082
rect 197358 377632 197414 377641
rect 197358 377567 197414 377576
rect 197360 376712 197412 376718
rect 197360 376654 197412 376660
rect 197372 376417 197400 376654
rect 197358 376408 197414 376417
rect 197358 376343 197414 376352
rect 197360 375352 197412 375358
rect 197360 375294 197412 375300
rect 197372 375193 197400 375294
rect 197358 375184 197414 375193
rect 197358 375119 197414 375128
rect 197360 373992 197412 373998
rect 197358 373960 197360 373969
rect 197412 373960 197414 373969
rect 197358 373895 197414 373904
rect 197358 372600 197414 372609
rect 197358 372535 197360 372544
rect 197412 372535 197414 372544
rect 197360 372506 197412 372512
rect 197452 372496 197504 372502
rect 197452 372438 197504 372444
rect 197464 371385 197492 372438
rect 197450 371376 197506 371385
rect 197450 371311 197506 371320
rect 197360 371204 197412 371210
rect 197360 371146 197412 371152
rect 197372 370161 197400 371146
rect 197358 370152 197414 370161
rect 197358 370087 197414 370096
rect 197360 369844 197412 369850
rect 197360 369786 197412 369792
rect 197372 368937 197400 369786
rect 197358 368928 197414 368937
rect 197358 368863 197414 368872
rect 197360 368484 197412 368490
rect 197360 368426 197412 368432
rect 197372 368393 197400 368426
rect 197358 368384 197414 368393
rect 197358 368319 197414 368328
rect 197360 367056 197412 367062
rect 197358 367024 197360 367033
rect 197412 367024 197414 367033
rect 197358 366959 197414 366968
rect 197360 365628 197412 365634
rect 197360 365570 197412 365576
rect 197372 365265 197400 365570
rect 197358 365256 197414 365265
rect 197358 365191 197414 365200
rect 197832 365158 197860 421631
rect 197820 365152 197872 365158
rect 197820 365094 197872 365100
rect 197360 364336 197412 364342
rect 197360 364278 197412 364284
rect 197372 364041 197400 364278
rect 197358 364032 197414 364041
rect 197358 363967 197414 363976
rect 197360 362908 197412 362914
rect 197360 362850 197412 362856
rect 197372 362817 197400 362850
rect 197358 362808 197414 362817
rect 197358 362743 197414 362752
rect 197360 361548 197412 361554
rect 197360 361490 197412 361496
rect 197372 361457 197400 361490
rect 197452 361480 197504 361486
rect 197358 361448 197414 361457
rect 197452 361422 197504 361428
rect 197358 361383 197414 361392
rect 197464 360233 197492 361422
rect 197450 360224 197506 360233
rect 197450 360159 197506 360168
rect 197360 360120 197412 360126
rect 197360 360062 197412 360068
rect 197372 359689 197400 360062
rect 197358 359680 197414 359689
rect 197358 359615 197414 359624
rect 197360 358692 197412 358698
rect 197360 358634 197412 358640
rect 197372 357785 197400 358634
rect 197358 357776 197414 357785
rect 197358 357711 197414 357720
rect 197360 357400 197412 357406
rect 197360 357342 197412 357348
rect 197372 356561 197400 357342
rect 197358 356552 197414 356561
rect 197358 356487 197414 356496
rect 197360 356040 197412 356046
rect 197360 355982 197412 355988
rect 197372 355337 197400 355982
rect 197358 355328 197414 355337
rect 197358 355263 197414 355272
rect 197360 354408 197412 354414
rect 197360 354350 197412 354356
rect 197372 354113 197400 354350
rect 197358 354104 197414 354113
rect 197358 354039 197414 354048
rect 197360 353252 197412 353258
rect 197360 353194 197412 353200
rect 197372 352889 197400 353194
rect 197358 352880 197414 352889
rect 197358 352815 197414 352824
rect 197360 351892 197412 351898
rect 197360 351834 197412 351840
rect 197372 351665 197400 351834
rect 197358 351656 197414 351665
rect 197358 351591 197414 351600
rect 197360 350532 197412 350538
rect 197360 350474 197412 350480
rect 197372 350441 197400 350474
rect 197358 350432 197414 350441
rect 197358 350367 197414 350376
rect 197360 349104 197412 349110
rect 197360 349046 197412 349052
rect 197450 349072 197506 349081
rect 197372 347857 197400 349046
rect 197450 349007 197452 349016
rect 197504 349007 197506 349016
rect 197452 348978 197504 348984
rect 197358 347848 197414 347857
rect 197358 347783 197414 347792
rect 197360 347676 197412 347682
rect 197360 347618 197412 347624
rect 197372 346633 197400 347618
rect 197358 346624 197414 346633
rect 197358 346559 197414 346568
rect 197360 346316 197412 346322
rect 197360 346258 197412 346264
rect 197372 345409 197400 346258
rect 197358 345400 197414 345409
rect 197358 345335 197414 345344
rect 197360 345024 197412 345030
rect 197360 344966 197412 344972
rect 197372 344865 197400 344966
rect 197358 344856 197414 344865
rect 197358 344791 197414 344800
rect 197360 343596 197412 343602
rect 197360 343538 197412 343544
rect 197372 343505 197400 343538
rect 197358 343496 197414 343505
rect 197358 343431 197414 343440
rect 197360 342236 197412 342242
rect 197360 342178 197412 342184
rect 197372 341737 197400 342178
rect 197358 341728 197414 341737
rect 197358 341663 197414 341672
rect 197360 340876 197412 340882
rect 197360 340818 197412 340824
rect 197372 340513 197400 340818
rect 197358 340504 197414 340513
rect 197358 340439 197414 340448
rect 197360 339448 197412 339454
rect 197360 339390 197412 339396
rect 197372 339289 197400 339390
rect 197358 339280 197414 339289
rect 197358 339215 197414 339224
rect 197360 338088 197412 338094
rect 197360 338030 197412 338036
rect 197372 337929 197400 338030
rect 197358 337920 197414 337929
rect 197358 337855 197414 337864
rect 197360 336728 197412 336734
rect 197360 336670 197412 336676
rect 197450 336696 197506 336705
rect 197372 336161 197400 336670
rect 197450 336631 197452 336640
rect 197504 336631 197506 336640
rect 197452 336602 197504 336608
rect 197358 336152 197414 336161
rect 197358 336087 197414 336096
rect 197360 335300 197412 335306
rect 197360 335242 197412 335248
rect 197372 334257 197400 335242
rect 197358 334248 197414 334257
rect 197358 334183 197414 334192
rect 197360 333940 197412 333946
rect 197360 333882 197412 333888
rect 197372 333033 197400 333882
rect 197358 333024 197414 333033
rect 197358 332959 197414 332968
rect 197360 332580 197412 332586
rect 197360 332522 197412 332528
rect 197372 331809 197400 332522
rect 197358 331800 197414 331809
rect 197358 331735 197414 331744
rect 197360 331220 197412 331226
rect 197360 331162 197412 331168
rect 197372 330585 197400 331162
rect 197358 330576 197414 330585
rect 197358 330511 197414 330520
rect 197360 329792 197412 329798
rect 197360 329734 197412 329740
rect 197372 329361 197400 329734
rect 197358 329352 197414 329361
rect 197358 329287 197414 329296
rect 197360 328432 197412 328438
rect 197358 328400 197360 328409
rect 197412 328400 197414 328409
rect 197358 328335 197414 328344
rect 197360 327072 197412 327078
rect 197358 327040 197360 327049
rect 197412 327040 197414 327049
rect 197358 326975 197414 326984
rect 197360 325644 197412 325650
rect 197360 325586 197412 325592
rect 197372 325553 197400 325586
rect 197358 325544 197414 325553
rect 197358 325479 197414 325488
rect 197358 324320 197414 324329
rect 197358 324255 197414 324264
rect 197452 324284 197504 324290
rect 197372 324222 197400 324255
rect 197452 324226 197504 324232
rect 197360 324216 197412 324222
rect 197360 324158 197412 324164
rect 197464 323105 197492 324226
rect 197450 323096 197506 323105
rect 197450 323031 197506 323040
rect 197360 322924 197412 322930
rect 197360 322866 197412 322872
rect 197372 321881 197400 322866
rect 197358 321872 197414 321881
rect 197358 321807 197414 321816
rect 197360 321564 197412 321570
rect 197360 321506 197412 321512
rect 197372 320657 197400 321506
rect 197358 320648 197414 320657
rect 197358 320583 197414 320592
rect 197360 320136 197412 320142
rect 197360 320078 197412 320084
rect 197372 319433 197400 320078
rect 197358 319424 197414 319433
rect 197358 319359 197414 319368
rect 197360 318776 197412 318782
rect 197360 318718 197412 318724
rect 197372 318209 197400 318718
rect 197358 318200 197414 318209
rect 197358 318135 197414 318144
rect 197360 317416 197412 317422
rect 197360 317358 197412 317364
rect 197372 316985 197400 317358
rect 197358 316976 197414 316985
rect 197358 316911 197414 316920
rect 197360 315988 197412 315994
rect 197360 315930 197412 315936
rect 197372 315761 197400 315930
rect 197358 315752 197414 315761
rect 197358 315687 197414 315696
rect 197360 314628 197412 314634
rect 197360 314570 197412 314576
rect 197372 314401 197400 314570
rect 197358 314392 197414 314401
rect 197358 314327 197414 314336
rect 197452 313268 197504 313274
rect 197452 313210 197504 313216
rect 197360 313200 197412 313206
rect 197358 313168 197360 313177
rect 197412 313168 197414 313177
rect 197358 313103 197414 313112
rect 197464 312633 197492 313210
rect 197450 312624 197506 312633
rect 197450 312559 197506 312568
rect 197360 311840 197412 311846
rect 197360 311782 197412 311788
rect 197372 311409 197400 311782
rect 197358 311400 197414 311409
rect 197358 311335 197414 311344
rect 197360 310480 197412 310486
rect 197360 310422 197412 310428
rect 197372 309505 197400 310422
rect 197358 309496 197414 309505
rect 197358 309431 197414 309440
rect 197360 309120 197412 309126
rect 197360 309062 197412 309068
rect 197372 308281 197400 309062
rect 197358 308272 197414 308281
rect 197358 308207 197414 308216
rect 197728 307760 197780 307766
rect 197728 307702 197780 307708
rect 197740 307057 197768 307702
rect 197726 307048 197782 307057
rect 197726 306983 197782 306992
rect 197360 306332 197412 306338
rect 197360 306274 197412 306280
rect 197372 305833 197400 306274
rect 197358 305824 197414 305833
rect 197358 305759 197414 305768
rect 197360 304972 197412 304978
rect 197360 304914 197412 304920
rect 197372 304609 197400 304914
rect 197358 304600 197414 304609
rect 197358 304535 197414 304544
rect 197360 303612 197412 303618
rect 197360 303554 197412 303560
rect 197372 303521 197400 303554
rect 197358 303512 197414 303521
rect 197358 303447 197414 303456
rect 197360 302184 197412 302190
rect 197360 302126 197412 302132
rect 197372 302025 197400 302126
rect 197358 302016 197414 302025
rect 197358 301951 197414 301960
rect 197360 300824 197412 300830
rect 197358 300792 197360 300801
rect 197412 300792 197414 300801
rect 197358 300727 197414 300736
rect 197358 299568 197414 299577
rect 197358 299503 197360 299512
rect 197412 299503 197414 299512
rect 197360 299474 197412 299480
rect 197358 298344 197414 298353
rect 197358 298279 197414 298288
rect 197372 298178 197400 298279
rect 197360 298172 197412 298178
rect 197360 298114 197412 298120
rect 197358 297120 197414 297129
rect 197358 297055 197414 297064
rect 197372 296750 197400 297055
rect 197360 296744 197412 296750
rect 197360 296686 197412 296692
rect 197358 295488 197414 295497
rect 197358 295423 197414 295432
rect 197372 295390 197400 295423
rect 197360 295384 197412 295390
rect 197360 295326 197412 295332
rect 197358 294400 197414 294409
rect 197358 294335 197414 294344
rect 197372 294030 197400 294335
rect 197360 294024 197412 294030
rect 197360 293966 197412 293972
rect 197358 293448 197414 293457
rect 197358 293383 197414 293392
rect 197372 292602 197400 293383
rect 197360 292596 197412 292602
rect 197360 292538 197412 292544
rect 197358 292088 197414 292097
rect 197358 292023 197414 292032
rect 197372 291242 197400 292023
rect 197360 291236 197412 291242
rect 197360 291178 197412 291184
rect 197358 290864 197414 290873
rect 197358 290799 197414 290808
rect 197372 289882 197400 290799
rect 197360 289876 197412 289882
rect 197360 289818 197412 289824
rect 197358 289640 197414 289649
rect 197358 289575 197414 289584
rect 197372 288454 197400 289575
rect 197360 288448 197412 288454
rect 197360 288390 197412 288396
rect 197450 288416 197506 288425
rect 197450 288351 197506 288360
rect 197358 287192 197414 287201
rect 197464 287162 197492 288351
rect 197358 287127 197414 287136
rect 197452 287156 197504 287162
rect 197372 287094 197400 287127
rect 197452 287098 197504 287104
rect 197360 287088 197412 287094
rect 197360 287030 197412 287036
rect 197358 285968 197414 285977
rect 197358 285903 197414 285912
rect 197372 285734 197400 285903
rect 197360 285728 197412 285734
rect 197360 285670 197412 285676
rect 197358 284744 197414 284753
rect 197358 284679 197414 284688
rect 197372 284374 197400 284679
rect 197360 284368 197412 284374
rect 197360 284310 197412 284316
rect 197358 283520 197414 283529
rect 197358 283455 197414 283464
rect 197372 282946 197400 283455
rect 197360 282940 197412 282946
rect 197360 282882 197412 282888
rect 197358 282296 197414 282305
rect 197358 282231 197414 282240
rect 197372 281586 197400 282231
rect 197360 281580 197412 281586
rect 197360 281522 197412 281528
rect 197358 281072 197414 281081
rect 197358 281007 197414 281016
rect 197372 280226 197400 281007
rect 197360 280220 197412 280226
rect 197360 280162 197412 280168
rect 197358 279168 197414 279177
rect 197358 279103 197414 279112
rect 197372 278798 197400 279103
rect 197360 278792 197412 278798
rect 197360 278734 197412 278740
rect 197358 278488 197414 278497
rect 197358 278423 197414 278432
rect 197372 277438 197400 278423
rect 197360 277432 197412 277438
rect 197360 277374 197412 277380
rect 197450 277264 197506 277273
rect 197450 277199 197506 277208
rect 197360 276140 197412 276146
rect 197360 276082 197412 276088
rect 197372 276049 197400 276082
rect 197464 276078 197492 277199
rect 197452 276072 197504 276078
rect 197358 276040 197414 276049
rect 197452 276014 197504 276020
rect 197358 275975 197414 275984
rect 197358 274816 197414 274825
rect 197358 274751 197414 274760
rect 197372 274718 197400 274751
rect 197360 274712 197412 274718
rect 197360 274654 197412 274660
rect 197358 273592 197414 273601
rect 197358 273527 197414 273536
rect 197372 273290 197400 273527
rect 197360 273284 197412 273290
rect 197360 273226 197412 273232
rect 197358 272368 197414 272377
rect 197358 272303 197414 272312
rect 197372 271930 197400 272303
rect 197360 271924 197412 271930
rect 197360 271866 197412 271872
rect 197358 270600 197414 270609
rect 197358 270535 197360 270544
rect 197412 270535 197414 270544
rect 197360 270506 197412 270512
rect 197818 269920 197874 269929
rect 197818 269855 197874 269864
rect 197358 268560 197414 268569
rect 197358 268495 197414 268504
rect 197372 267782 197400 268495
rect 197360 267776 197412 267782
rect 197360 267718 197412 267724
rect 197358 267336 197414 267345
rect 197358 267271 197414 267280
rect 197372 266422 197400 267271
rect 197360 266416 197412 266422
rect 197360 266358 197412 266364
rect 197358 266112 197414 266121
rect 197358 266047 197414 266056
rect 197372 264994 197400 266047
rect 197360 264988 197412 264994
rect 197360 264930 197412 264936
rect 197450 264888 197506 264897
rect 197450 264823 197506 264832
rect 197464 263702 197492 264823
rect 197452 263696 197504 263702
rect 197358 263664 197414 263673
rect 197452 263638 197504 263644
rect 197358 263599 197360 263608
rect 197412 263599 197414 263608
rect 197360 263570 197412 263576
rect 197358 262440 197414 262449
rect 197358 262375 197414 262384
rect 197372 262274 197400 262375
rect 197360 262268 197412 262274
rect 197360 262210 197412 262216
rect 197358 261216 197414 261225
rect 197358 261151 197414 261160
rect 197372 260914 197400 261151
rect 197360 260908 197412 260914
rect 197360 260850 197412 260856
rect 197358 258768 197414 258777
rect 197358 258703 197414 258712
rect 197372 258126 197400 258703
rect 197360 258120 197412 258126
rect 197360 258062 197412 258068
rect 197542 254824 197598 254833
rect 197542 254759 197598 254768
rect 197450 252512 197506 252521
rect 197450 252447 197452 252456
rect 197504 252447 197506 252456
rect 197452 252418 197504 252424
rect 197360 252408 197412 252414
rect 197360 252350 197412 252356
rect 197372 251297 197400 252350
rect 197556 251569 197584 254759
rect 197832 254590 197860 269855
rect 197924 257417 197952 448462
rect 198002 448423 198058 448432
rect 197910 257408 197966 257417
rect 197910 257343 197966 257352
rect 197820 254584 197872 254590
rect 197820 254526 197872 254532
rect 197924 253910 197952 257343
rect 198016 256193 198044 448423
rect 198108 448361 198136 470319
rect 198094 448352 198150 448361
rect 198094 448287 198150 448296
rect 198002 256184 198058 256193
rect 198002 256119 198058 256128
rect 197912 253904 197964 253910
rect 197912 253846 197964 253852
rect 198016 252550 198044 256119
rect 198108 254833 198136 448287
rect 198200 448225 198228 471679
rect 198186 448216 198242 448225
rect 198186 448151 198242 448160
rect 198094 254824 198150 254833
rect 198094 254759 198150 254768
rect 198200 253881 198228 448151
rect 198292 448089 198320 473311
rect 198384 451586 198412 574631
rect 198556 574456 198608 574462
rect 198556 574398 198608 574404
rect 198464 572620 198516 572626
rect 198464 572562 198516 572568
rect 198372 451580 198424 451586
rect 198372 451522 198424 451528
rect 198278 448080 198334 448089
rect 198278 448015 198334 448024
rect 198186 253872 198242 253881
rect 198186 253807 198242 253816
rect 198004 252544 198056 252550
rect 198292 252521 198320 448015
rect 198476 445534 198504 572562
rect 198568 448186 198596 574398
rect 198556 448180 198608 448186
rect 198556 448122 198608 448128
rect 198660 447778 198688 575010
rect 199200 474836 199252 474842
rect 199200 474778 199252 474784
rect 198740 454164 198792 454170
rect 198740 454106 198792 454112
rect 198752 452198 198780 454106
rect 199212 453082 199240 474778
rect 199292 474768 199344 474774
rect 199292 474710 199344 474716
rect 199304 453286 199332 474710
rect 199292 453280 199344 453286
rect 199292 453222 199344 453228
rect 199200 453076 199252 453082
rect 199200 453018 199252 453024
rect 198740 452192 198792 452198
rect 198740 452134 198792 452140
rect 199396 448322 199424 575146
rect 199844 575000 199896 575006
rect 199844 574942 199896 574948
rect 199752 574388 199804 574394
rect 199752 574330 199804 574336
rect 199568 572688 199620 572694
rect 199568 572630 199620 572636
rect 199476 571940 199528 571946
rect 199476 571882 199528 571888
rect 199384 448316 199436 448322
rect 199384 448258 199436 448264
rect 198648 447772 198700 447778
rect 198648 447714 198700 447720
rect 198464 445528 198516 445534
rect 198464 445470 198516 445476
rect 199488 445262 199516 571882
rect 199580 445466 199608 572630
rect 199660 571872 199712 571878
rect 199660 571814 199712 571820
rect 199568 445460 199620 445466
rect 199568 445402 199620 445408
rect 199672 445330 199700 571814
rect 199764 448254 199792 574330
rect 199752 448248 199804 448254
rect 199752 448190 199804 448196
rect 199856 445738 199884 574942
rect 237208 570654 237236 591631
rect 237196 570648 237248 570654
rect 237196 570590 237248 570596
rect 237300 543017 237328 654463
rect 336738 603800 336794 603809
rect 336738 603735 336794 603744
rect 238666 594688 238722 594697
rect 238666 594623 238722 594632
rect 238574 593056 238630 593065
rect 238574 592991 238630 593000
rect 238588 544406 238616 592991
rect 238576 544400 238628 544406
rect 238576 544342 238628 544348
rect 238680 543046 238708 594623
rect 253110 576192 253166 576201
rect 253110 576127 253166 576136
rect 292486 576192 292542 576201
rect 292486 576127 292542 576136
rect 253124 567866 253152 576127
rect 284206 575376 284262 575385
rect 284206 575311 284262 575320
rect 285310 575376 285366 575385
rect 285310 575311 285366 575320
rect 286598 575376 286654 575385
rect 286598 575311 286654 575320
rect 287886 575376 287942 575385
rect 287886 575311 287942 575320
rect 280158 575104 280214 575113
rect 280158 575039 280214 575048
rect 280172 575006 280200 575039
rect 280160 575000 280212 575006
rect 280160 574942 280212 574948
rect 280250 574968 280306 574977
rect 280250 574903 280252 574912
rect 280304 574903 280306 574912
rect 281538 574968 281594 574977
rect 281538 574903 281594 574912
rect 280252 574874 280304 574880
rect 281552 574870 281580 574903
rect 281540 574864 281592 574870
rect 281540 574806 281592 574812
rect 253754 574424 253810 574433
rect 253754 574359 253810 574368
rect 273258 574424 273314 574433
rect 273258 574359 273314 574368
rect 276018 574424 276074 574433
rect 276018 574359 276074 574368
rect 253768 569226 253796 574359
rect 254582 574288 254638 574297
rect 254582 574223 254638 574232
rect 269210 574288 269266 574297
rect 269210 574223 269266 574232
rect 253846 574152 253902 574161
rect 253846 574087 253902 574096
rect 253756 569220 253808 569226
rect 253756 569162 253808 569168
rect 253112 567860 253164 567866
rect 253112 567802 253164 567808
rect 253860 562358 253888 574087
rect 253848 562352 253900 562358
rect 253848 562294 253900 562300
rect 254596 545766 254624 574223
rect 269118 574152 269174 574161
rect 269118 574087 269174 574096
rect 269132 573442 269160 574087
rect 269120 573436 269172 573442
rect 269120 573378 269172 573384
rect 269224 569362 269252 574223
rect 270498 574152 270554 574161
rect 270498 574087 270554 574096
rect 271878 574152 271934 574161
rect 271878 574087 271934 574096
rect 270512 569430 270540 574087
rect 270500 569424 270552 569430
rect 270500 569366 270552 569372
rect 269212 569356 269264 569362
rect 269212 569298 269264 569304
rect 271892 569294 271920 574087
rect 273272 571878 273300 574359
rect 274638 574288 274694 574297
rect 274638 574223 274694 574232
rect 274652 571946 274680 574223
rect 276032 572694 276060 574359
rect 284220 574326 284248 575311
rect 284390 575240 284446 575249
rect 284390 575175 284446 575184
rect 284298 574832 284354 574841
rect 284298 574767 284300 574776
rect 284352 574767 284354 574776
rect 284300 574738 284352 574744
rect 284404 574734 284432 575175
rect 284392 574728 284444 574734
rect 284392 574670 284444 574676
rect 285324 574666 285352 575311
rect 285312 574660 285364 574666
rect 285312 574602 285364 574608
rect 284208 574320 284260 574326
rect 278778 574288 278834 574297
rect 284208 574262 284260 574268
rect 285678 574288 285734 574297
rect 278778 574223 278834 574232
rect 285678 574223 285734 574232
rect 277674 574152 277730 574161
rect 277674 574087 277730 574096
rect 278686 574152 278742 574161
rect 278686 574087 278742 574096
rect 276020 572688 276072 572694
rect 276020 572630 276072 572636
rect 277688 572626 277716 574087
rect 277676 572620 277728 572626
rect 277676 572562 277728 572568
rect 274640 571940 274692 571946
rect 274640 571882 274692 571888
rect 273260 571872 273312 571878
rect 273260 571814 273312 571820
rect 271880 569288 271932 569294
rect 271880 569230 271932 569236
rect 254584 545760 254636 545766
rect 254584 545702 254636 545708
rect 238668 543040 238720 543046
rect 237286 543008 237342 543017
rect 238668 542982 238720 542988
rect 237286 542943 237342 542952
rect 278700 540394 278728 574087
rect 278792 572558 278820 574223
rect 285692 574190 285720 574223
rect 286612 574190 286640 575311
rect 287518 574968 287574 574977
rect 287518 574903 287574 574912
rect 287532 574598 287560 574903
rect 287520 574592 287572 574598
rect 287520 574534 287572 574540
rect 287900 574530 287928 575311
rect 289818 575240 289874 575249
rect 289818 575175 289874 575184
rect 289832 575142 289860 575175
rect 289820 575136 289872 575142
rect 289820 575078 289872 575084
rect 291198 575104 291254 575113
rect 291198 575039 291254 575048
rect 291106 574968 291162 574977
rect 291106 574903 291162 574912
rect 288438 574832 288494 574841
rect 288438 574767 288494 574776
rect 291014 574832 291070 574841
rect 291014 574767 291070 574776
rect 287888 574524 287940 574530
rect 287888 574466 287940 574472
rect 288452 574258 288480 574767
rect 289726 574560 289782 574569
rect 289726 574495 289782 574504
rect 288440 574252 288492 574258
rect 288440 574194 288492 574200
rect 285680 574184 285732 574190
rect 280066 574152 280122 574161
rect 280066 574087 280122 574096
rect 281446 574152 281502 574161
rect 281446 574087 281502 574096
rect 282826 574152 282882 574161
rect 282826 574087 282882 574096
rect 284206 574152 284262 574161
rect 285680 574126 285732 574132
rect 286600 574184 286652 574190
rect 286600 574126 286652 574132
rect 284206 574087 284262 574096
rect 278780 572552 278832 572558
rect 278780 572494 278832 572500
rect 280080 540462 280108 574087
rect 280068 540456 280120 540462
rect 280068 540398 280120 540404
rect 278688 540388 278740 540394
rect 278688 540330 278740 540336
rect 218060 540320 218112 540326
rect 218060 540262 218112 540268
rect 217600 540252 217652 540258
rect 217600 540194 217652 540200
rect 205732 539980 205784 539986
rect 205732 539922 205784 539928
rect 205744 539209 205772 539922
rect 217612 539753 217640 540194
rect 218072 539918 218100 540262
rect 218060 539912 218112 539918
rect 218060 539854 218112 539860
rect 217598 539744 217654 539753
rect 217598 539679 217654 539688
rect 218072 539617 218100 539854
rect 218058 539608 218114 539617
rect 218058 539543 218114 539552
rect 205730 539200 205786 539209
rect 205730 539135 205786 539144
rect 281460 538898 281488 574087
rect 282840 538966 282868 574087
rect 284220 539034 284248 574087
rect 289740 572558 289768 574495
rect 291028 572694 291056 574767
rect 291016 572688 291068 572694
rect 291016 572630 291068 572636
rect 291120 572626 291148 574903
rect 291212 574462 291240 575039
rect 291200 574456 291252 574462
rect 291200 574398 291252 574404
rect 292500 574258 292528 576127
rect 330208 575476 330260 575482
rect 330208 575418 330260 575424
rect 330220 575385 330248 575418
rect 297914 575376 297970 575385
rect 297914 575311 297970 575320
rect 300674 575376 300730 575385
rect 300674 575311 300730 575320
rect 301870 575376 301926 575385
rect 301870 575311 301926 575320
rect 302882 575376 302938 575385
rect 302882 575311 302938 575320
rect 304630 575376 304686 575385
rect 304630 575311 304686 575320
rect 305550 575376 305606 575385
rect 305550 575311 305606 575320
rect 306286 575376 306342 575385
rect 306286 575311 306342 575320
rect 307574 575376 307630 575385
rect 307574 575311 307630 575320
rect 320454 575376 320510 575385
rect 320454 575311 320510 575320
rect 330206 575376 330262 575385
rect 330206 575311 330262 575320
rect 330482 575376 330538 575385
rect 330482 575311 330538 575320
rect 293958 575240 294014 575249
rect 293958 575175 293960 575184
rect 294012 575175 294014 575184
rect 293960 575146 294012 575152
rect 293958 575104 294014 575113
rect 293958 575039 293960 575048
rect 294012 575039 294014 575048
rect 293960 575010 294012 575016
rect 292578 574832 292634 574841
rect 292578 574767 292634 574776
rect 292592 574394 292620 574767
rect 296534 574560 296590 574569
rect 296534 574495 296590 574504
rect 293774 574424 293830 574433
rect 292580 574388 292632 574394
rect 293774 574359 293830 574368
rect 294694 574424 294750 574433
rect 294694 574359 294750 574368
rect 292580 574330 292632 574336
rect 292488 574252 292540 574258
rect 292488 574194 292540 574200
rect 291108 572620 291160 572626
rect 291108 572562 291160 572568
rect 289728 572552 289780 572558
rect 289728 572494 289780 572500
rect 293788 571946 293816 574359
rect 293776 571940 293828 571946
rect 293776 571882 293828 571888
rect 294708 571878 294736 574359
rect 295338 574152 295394 574161
rect 295338 574087 295394 574096
rect 295352 572490 295380 574087
rect 296548 572490 296576 574495
rect 297928 574394 297956 575311
rect 298926 574560 298982 574569
rect 298926 574495 298982 574504
rect 299202 574560 299258 574569
rect 299202 574495 299258 574504
rect 299478 574560 299534 574569
rect 299478 574495 299534 574504
rect 297916 574388 297968 574394
rect 297916 574330 297968 574336
rect 298190 574288 298246 574297
rect 298190 574223 298246 574232
rect 298098 574152 298154 574161
rect 298098 574087 298154 574096
rect 295340 572484 295392 572490
rect 295340 572426 295392 572432
rect 296536 572484 296588 572490
rect 296536 572426 296588 572432
rect 298112 572422 298140 574087
rect 298100 572416 298152 572422
rect 298100 572358 298152 572364
rect 298204 572286 298232 574223
rect 298940 572286 298968 574495
rect 299216 572422 299244 574495
rect 299204 572416 299256 572422
rect 299204 572358 299256 572364
rect 299492 572354 299520 574495
rect 300688 574462 300716 575311
rect 301884 575074 301912 575311
rect 301872 575068 301924 575074
rect 301872 575010 301924 575016
rect 302896 574598 302924 575311
rect 304644 574870 304672 575311
rect 304632 574864 304684 574870
rect 304632 574806 304684 574812
rect 305564 574802 305592 575311
rect 305552 574796 305604 574802
rect 305552 574738 305604 574744
rect 306300 574734 306328 575311
rect 307588 574938 307616 575311
rect 320468 575006 320496 575311
rect 330496 575006 330524 575311
rect 320456 575000 320508 575006
rect 320456 574942 320508 574948
rect 330484 575000 330536 575006
rect 330484 574942 330536 574948
rect 307576 574932 307628 574938
rect 307576 574874 307628 574880
rect 306288 574728 306340 574734
rect 306288 574670 306340 574676
rect 302884 574592 302936 574598
rect 302884 574534 302936 574540
rect 300676 574456 300728 574462
rect 300676 574398 300728 574404
rect 303618 574288 303674 574297
rect 303618 574223 303674 574232
rect 300858 574152 300914 574161
rect 300858 574087 300914 574096
rect 302238 574152 302294 574161
rect 302238 574087 302294 574096
rect 299480 572348 299532 572354
rect 299480 572290 299532 572296
rect 298192 572280 298244 572286
rect 298192 572222 298244 572228
rect 298928 572280 298980 572286
rect 298928 572222 298980 572228
rect 300872 572150 300900 574087
rect 302252 572218 302280 574087
rect 302240 572212 302292 572218
rect 302240 572154 302292 572160
rect 300860 572144 300912 572150
rect 300860 572086 300912 572092
rect 303632 572082 303660 574223
rect 304998 574152 305054 574161
rect 304998 574087 305054 574096
rect 306470 574152 306526 574161
rect 306470 574087 306472 574096
rect 303620 572076 303672 572082
rect 303620 572018 303672 572024
rect 305012 572014 305040 574087
rect 306524 574087 306526 574096
rect 318706 574152 318762 574161
rect 318706 574087 318762 574096
rect 306472 574058 306524 574064
rect 305000 572008 305052 572014
rect 305000 571950 305052 571956
rect 294696 571872 294748 571878
rect 294696 571814 294748 571820
rect 318720 539102 318748 574087
rect 318708 539096 318760 539102
rect 318708 539038 318760 539044
rect 284208 539028 284260 539034
rect 284208 538970 284260 538976
rect 282828 538960 282880 538966
rect 282828 538902 282880 538908
rect 281448 538892 281500 538898
rect 281448 538834 281500 538840
rect 336280 453892 336332 453898
rect 336280 453834 336332 453840
rect 288898 453792 288954 453801
rect 294786 453792 294842 453801
rect 288898 453727 288954 453736
rect 291016 453756 291068 453762
rect 213182 453656 213238 453665
rect 213182 453591 213238 453600
rect 284298 453656 284354 453665
rect 284298 453591 284354 453600
rect 286782 453656 286838 453665
rect 286782 453591 286838 453600
rect 201776 451648 201828 451654
rect 201776 451590 201828 451596
rect 200212 451580 200264 451586
rect 200212 451522 200264 451528
rect 199844 445732 199896 445738
rect 199844 445674 199896 445680
rect 199660 445324 199712 445330
rect 199660 445266 199712 445272
rect 199476 445256 199528 445262
rect 199476 445198 199528 445204
rect 198556 431384 198608 431390
rect 198556 431326 198608 431332
rect 198372 431248 198424 431254
rect 198372 431190 198424 431196
rect 198004 252486 198056 252492
rect 198278 252512 198334 252521
rect 198278 252447 198334 252456
rect 197542 251560 197598 251569
rect 197542 251495 197598 251504
rect 197358 251288 197414 251297
rect 197358 251223 197414 251232
rect 197266 248840 197322 248849
rect 197266 248775 197322 248784
rect 197360 247036 197412 247042
rect 197360 246978 197412 246984
rect 197372 246401 197400 246978
rect 197358 246392 197414 246401
rect 197358 246327 197414 246336
rect 197360 245608 197412 245614
rect 197360 245550 197412 245556
rect 197372 245041 197400 245550
rect 197358 245032 197414 245041
rect 197358 244967 197414 244976
rect 197360 244248 197412 244254
rect 197360 244190 197412 244196
rect 197372 243817 197400 244190
rect 197358 243808 197414 243817
rect 197358 243743 197414 243752
rect 197360 242888 197412 242894
rect 197360 242830 197412 242836
rect 197372 242593 197400 242830
rect 197358 242584 197414 242593
rect 197358 242519 197414 242528
rect 196900 242208 196952 242214
rect 196900 242150 196952 242156
rect 196808 215416 196860 215422
rect 196808 215358 196860 215364
rect 196912 180794 196940 242150
rect 197542 241360 197598 241369
rect 197542 241295 197598 241304
rect 197450 239592 197506 239601
rect 197450 239527 197506 239536
rect 197360 238944 197412 238950
rect 197358 238912 197360 238921
rect 197412 238912 197414 238921
rect 197358 238847 197414 238856
rect 197360 238060 197412 238066
rect 197360 238002 197412 238008
rect 197372 236473 197400 238002
rect 197464 236706 197492 239527
rect 197452 236700 197504 236706
rect 197452 236642 197504 236648
rect 197358 236464 197414 236473
rect 197358 236399 197414 236408
rect 197556 235278 197584 241295
rect 197728 235952 197780 235958
rect 197728 235894 197780 235900
rect 197544 235272 197596 235278
rect 197740 235249 197768 235894
rect 197544 235214 197596 235220
rect 197726 235240 197782 235249
rect 197726 235175 197782 235184
rect 197358 233880 197414 233889
rect 197358 233815 197414 233824
rect 197372 233306 197400 233815
rect 197360 233300 197412 233306
rect 197360 233242 197412 233248
rect 197358 232656 197414 232665
rect 197358 232591 197414 232600
rect 197818 232656 197874 232665
rect 197818 232591 197874 232600
rect 197372 232558 197400 232591
rect 197360 232552 197412 232558
rect 197360 232494 197412 232500
rect 197360 231804 197412 231810
rect 197360 231746 197412 231752
rect 197372 231713 197400 231746
rect 197358 231704 197414 231713
rect 197358 231639 197414 231648
rect 197542 230208 197598 230217
rect 197542 230143 197598 230152
rect 197556 229770 197584 230143
rect 197544 229764 197596 229770
rect 197544 229706 197596 229712
rect 197556 229094 197584 229706
rect 197464 229066 197584 229094
rect 197360 224256 197412 224262
rect 197360 224198 197412 224204
rect 197372 224097 197400 224198
rect 197358 224088 197414 224097
rect 197358 224023 197414 224032
rect 197358 220280 197414 220289
rect 197358 220215 197414 220224
rect 197372 220114 197400 220215
rect 197360 220108 197412 220114
rect 197360 220050 197412 220056
rect 197360 218000 197412 218006
rect 197360 217942 197412 217948
rect 197372 217841 197400 217942
rect 197358 217832 197414 217841
rect 197358 217767 197414 217776
rect 197358 216608 197414 216617
rect 197358 216543 197414 216552
rect 197372 215966 197400 216543
rect 197360 215960 197412 215966
rect 197360 215902 197412 215908
rect 197358 214160 197414 214169
rect 197358 214095 197414 214104
rect 197372 213994 197400 214095
rect 197360 213988 197412 213994
rect 197360 213930 197412 213936
rect 197358 212936 197414 212945
rect 197358 212871 197414 212880
rect 197372 212566 197400 212871
rect 197360 212560 197412 212566
rect 197360 212502 197412 212508
rect 197360 211132 197412 211138
rect 197360 211074 197412 211080
rect 197372 210361 197400 211074
rect 197358 210352 197414 210361
rect 197358 210287 197414 210296
rect 197360 210248 197412 210254
rect 197360 210190 197412 210196
rect 197372 209234 197400 210190
rect 197360 209228 197412 209234
rect 197360 209170 197412 209176
rect 197360 208344 197412 208350
rect 197358 208312 197360 208321
rect 197412 208312 197414 208321
rect 197358 208247 197414 208256
rect 197358 206680 197414 206689
rect 197358 206615 197414 206624
rect 197372 206378 197400 206615
rect 197360 206372 197412 206378
rect 197360 206314 197412 206320
rect 197358 205456 197414 205465
rect 197358 205391 197414 205400
rect 197372 204338 197400 205391
rect 197360 204332 197412 204338
rect 197360 204274 197412 204280
rect 197358 204232 197414 204241
rect 197358 204167 197360 204176
rect 197412 204167 197414 204176
rect 197360 204138 197412 204144
rect 197358 201784 197414 201793
rect 197358 201719 197414 201728
rect 197372 201550 197400 201719
rect 197360 201544 197412 201550
rect 197360 201486 197412 201492
rect 197360 200796 197412 200802
rect 197360 200738 197412 200744
rect 197372 200569 197400 200738
rect 197358 200560 197414 200569
rect 197358 200495 197414 200504
rect 197360 199436 197412 199442
rect 197360 199378 197412 199384
rect 197372 199209 197400 199378
rect 197358 199200 197414 199209
rect 197358 199135 197414 199144
rect 197360 198008 197412 198014
rect 197358 197976 197360 197985
rect 197412 197976 197414 197985
rect 197358 197911 197414 197920
rect 197360 197328 197412 197334
rect 197360 197270 197412 197276
rect 197372 196761 197400 197270
rect 197358 196752 197414 196761
rect 197358 196687 197414 196696
rect 197360 195968 197412 195974
rect 197360 195910 197412 195916
rect 197372 195537 197400 195910
rect 197358 195528 197414 195537
rect 197358 195463 197414 195472
rect 197360 194540 197412 194546
rect 197360 194482 197412 194488
rect 197372 194313 197400 194482
rect 197358 194304 197414 194313
rect 197358 194239 197414 194248
rect 197358 193080 197414 193089
rect 197358 193015 197414 193024
rect 197372 191894 197400 193015
rect 197360 191888 197412 191894
rect 197360 191830 197412 191836
rect 197360 191140 197412 191146
rect 197360 191082 197412 191088
rect 197372 190641 197400 191082
rect 197358 190632 197414 190641
rect 197358 190567 197414 190576
rect 197360 189780 197412 189786
rect 197360 189722 197412 189728
rect 197372 189417 197400 189722
rect 197358 189408 197414 189417
rect 197358 189343 197414 189352
rect 197360 188352 197412 188358
rect 197360 188294 197412 188300
rect 197372 188193 197400 188294
rect 197358 188184 197414 188193
rect 197358 188119 197414 188128
rect 197360 186992 197412 186998
rect 197360 186934 197412 186940
rect 197372 186833 197400 186934
rect 197358 186824 197414 186833
rect 197358 186759 197414 186768
rect 197360 185632 197412 185638
rect 197358 185600 197360 185609
rect 197412 185600 197414 185609
rect 197358 185535 197414 185544
rect 197358 184240 197414 184249
rect 197358 184175 197360 184184
rect 197412 184175 197414 184184
rect 197360 184146 197412 184152
rect 197358 182880 197414 182889
rect 197358 182815 197360 182824
rect 197412 182815 197414 182824
rect 197360 182786 197412 182792
rect 197360 182164 197412 182170
rect 197360 182106 197412 182112
rect 197372 181937 197400 182106
rect 197358 181928 197414 181937
rect 197358 181863 197414 181872
rect 196820 180766 196940 180794
rect 196820 178294 196848 180766
rect 197358 180704 197414 180713
rect 197358 180639 197414 180648
rect 197372 180130 197400 180639
rect 197360 180124 197412 180130
rect 197360 180066 197412 180072
rect 197360 179512 197412 179518
rect 197358 179480 197360 179489
rect 197412 179480 197414 179489
rect 197358 179415 197414 179424
rect 196808 178288 196860 178294
rect 196808 178230 196860 178236
rect 196716 115252 196768 115258
rect 196716 115194 196768 115200
rect 196624 113824 196676 113830
rect 196624 113766 196676 113772
rect 196624 57860 196676 57866
rect 196624 57802 196676 57808
rect 195980 32428 196032 32434
rect 195980 32370 196032 32376
rect 195244 22704 195296 22710
rect 195244 22646 195296 22652
rect 195992 16574 196020 32370
rect 194612 16546 195192 16574
rect 195992 16546 196572 16574
rect 194416 3596 194468 3602
rect 194416 3538 194468 3544
rect 193232 3454 193352 3482
rect 193232 480 193260 3454
rect 194428 480 194456 3538
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196544 3482 196572 16546
rect 196636 3602 196664 57802
rect 196820 26353 196848 178230
rect 197360 177336 197412 177342
rect 197360 177278 197412 177284
rect 197372 177041 197400 177278
rect 197358 177032 197414 177041
rect 197358 176967 197414 176976
rect 197360 175704 197412 175710
rect 197358 175672 197360 175681
rect 197412 175672 197414 175681
rect 197358 175607 197414 175616
rect 197360 175228 197412 175234
rect 197360 175170 197412 175176
rect 197372 174457 197400 175170
rect 197358 174448 197414 174457
rect 197358 174383 197414 174392
rect 197360 173256 197412 173262
rect 197358 173224 197360 173233
rect 197412 173224 197414 173233
rect 197358 173159 197414 173168
rect 197360 172508 197412 172514
rect 197360 172450 197412 172456
rect 197372 172009 197400 172450
rect 197358 172000 197414 172009
rect 197358 171935 197414 171944
rect 197358 170776 197414 170785
rect 197358 170711 197414 170720
rect 197372 170474 197400 170711
rect 197360 170468 197412 170474
rect 197360 170410 197412 170416
rect 197360 169720 197412 169726
rect 197360 169662 197412 169668
rect 197372 169561 197400 169662
rect 197358 169552 197414 169561
rect 197358 169487 197414 169496
rect 197358 167784 197414 167793
rect 197358 167719 197414 167728
rect 197372 167686 197400 167719
rect 197360 167680 197412 167686
rect 197360 167622 197412 167628
rect 197360 167000 197412 167006
rect 197360 166942 197412 166948
rect 197372 165889 197400 166942
rect 197358 165880 197414 165889
rect 197358 165815 197414 165824
rect 197360 164960 197412 164966
rect 197360 164902 197412 164908
rect 197372 164529 197400 164902
rect 197358 164520 197414 164529
rect 197358 164455 197414 164464
rect 197360 164212 197412 164218
rect 197360 164154 197412 164160
rect 197372 163305 197400 164154
rect 197358 163296 197414 163305
rect 197358 163231 197414 163240
rect 197360 162172 197412 162178
rect 197360 162114 197412 162120
rect 197372 162081 197400 162114
rect 197358 162072 197414 162081
rect 197358 162007 197414 162016
rect 197360 161424 197412 161430
rect 197360 161366 197412 161372
rect 197372 160857 197400 161366
rect 197358 160848 197414 160857
rect 197358 160783 197414 160792
rect 197358 159488 197414 159497
rect 197358 159423 197414 159432
rect 197372 159390 197400 159423
rect 197360 159384 197412 159390
rect 197360 159326 197412 159332
rect 197358 158400 197414 158409
rect 197358 158335 197360 158344
rect 197412 158335 197414 158344
rect 197360 158306 197412 158312
rect 197358 157176 197414 157185
rect 197358 157111 197414 157120
rect 197372 156670 197400 157111
rect 197360 156664 197412 156670
rect 197360 156606 197412 156612
rect 197358 155952 197414 155961
rect 197358 155887 197414 155896
rect 197372 155242 197400 155887
rect 197360 155236 197412 155242
rect 197360 155178 197412 155184
rect 197360 154556 197412 154562
rect 197360 154498 197412 154504
rect 197372 153513 197400 154498
rect 197358 153504 197414 153513
rect 197358 153439 197414 153448
rect 197360 153196 197412 153202
rect 197360 153138 197412 153144
rect 197372 152833 197400 153138
rect 197358 152824 197414 152833
rect 197358 152759 197414 152768
rect 197358 150512 197414 150521
rect 197358 150447 197360 150456
rect 197412 150447 197414 150456
rect 197360 150418 197412 150424
rect 197358 149696 197414 149705
rect 197358 149631 197414 149640
rect 197372 149122 197400 149631
rect 197360 149116 197412 149122
rect 197360 149058 197412 149064
rect 197360 147620 197412 147626
rect 197360 147562 197412 147568
rect 197372 147257 197400 147562
rect 197358 147248 197414 147257
rect 197358 147183 197414 147192
rect 197358 146024 197414 146033
rect 197358 145959 197414 145968
rect 197372 144974 197400 145959
rect 197360 144968 197412 144974
rect 197360 144910 197412 144916
rect 197358 144800 197414 144809
rect 197358 144735 197360 144744
rect 197412 144735 197414 144744
rect 197360 144706 197412 144712
rect 197360 143608 197412 143614
rect 197358 143576 197360 143585
rect 197412 143576 197414 143585
rect 197358 143511 197414 143520
rect 197358 142352 197414 142361
rect 197358 142287 197414 142296
rect 197372 142186 197400 142287
rect 197360 142180 197412 142186
rect 197360 142122 197412 142128
rect 197464 141438 197492 229066
rect 197542 226536 197598 226545
rect 197542 226471 197598 226480
rect 197556 170406 197584 226471
rect 197728 215416 197780 215422
rect 197728 215358 197780 215364
rect 197636 212492 197688 212498
rect 197636 212434 197688 212440
rect 197648 211721 197676 212434
rect 197634 211712 197690 211721
rect 197634 211647 197690 211656
rect 197636 211608 197688 211614
rect 197636 211550 197688 211556
rect 197648 175982 197676 211550
rect 197740 210254 197768 215358
rect 197832 210362 197860 232591
rect 198384 229090 198412 431190
rect 198464 428596 198516 428602
rect 198464 428538 198516 428544
rect 198372 229084 198424 229090
rect 198372 229026 198424 229032
rect 198384 228993 198412 229026
rect 198370 228984 198426 228993
rect 198370 228919 198426 228928
rect 198476 226302 198504 428538
rect 198568 227730 198596 431326
rect 199200 431316 199252 431322
rect 199200 431258 199252 431264
rect 198740 430160 198792 430166
rect 198740 430102 198792 430108
rect 198648 429956 198700 429962
rect 198648 429898 198700 429904
rect 198556 227724 198608 227730
rect 198556 227666 198608 227672
rect 198568 226545 198596 227666
rect 198554 226536 198610 226545
rect 198554 226471 198610 226480
rect 198464 226296 198516 226302
rect 198464 226238 198516 226244
rect 198476 225321 198504 226238
rect 198462 225312 198518 225321
rect 198462 225247 198518 225256
rect 198660 224097 198688 429898
rect 198752 345710 198780 430102
rect 198924 430092 198976 430098
rect 198924 430034 198976 430040
rect 198832 428664 198884 428670
rect 198832 428606 198884 428612
rect 198844 427650 198872 428606
rect 198832 427644 198884 427650
rect 198832 427586 198884 427592
rect 198844 351286 198872 427586
rect 198832 351280 198884 351286
rect 198832 351222 198884 351228
rect 198740 345704 198792 345710
rect 198740 345646 198792 345652
rect 198646 224088 198702 224097
rect 198646 224023 198702 224032
rect 198752 220289 198780 345646
rect 198936 229022 198964 430034
rect 199016 430024 199068 430030
rect 199016 429966 199068 429972
rect 198924 229016 198976 229022
rect 198924 228958 198976 228964
rect 198936 221513 198964 228958
rect 199028 223582 199056 429966
rect 199108 429888 199160 429894
rect 199108 429830 199160 429836
rect 199120 228478 199148 429830
rect 199212 230217 199240 431258
rect 199290 425776 199346 425785
rect 199290 425711 199346 425720
rect 199304 237697 199332 425711
rect 199384 422952 199436 422958
rect 199384 422894 199436 422900
rect 199396 259593 199424 422894
rect 199568 421592 199620 421598
rect 199568 421534 199620 421540
rect 200118 421560 200174 421569
rect 199476 420232 199528 420238
rect 199476 420174 199528 420180
rect 199382 259584 199438 259593
rect 199382 259519 199438 259528
rect 199488 258777 199516 420174
rect 199580 365090 199608 421534
rect 200118 421495 200174 421504
rect 199568 365084 199620 365090
rect 199568 365026 199620 365032
rect 200132 365022 200160 421495
rect 200224 419139 200252 451522
rect 200224 419111 200598 419139
rect 201788 419125 201816 451590
rect 213196 451489 213224 453591
rect 278044 453552 278096 453558
rect 278044 453494 278096 453500
rect 231766 452568 231822 452577
rect 231766 452503 231822 452512
rect 234526 452568 234582 452577
rect 234526 452503 234582 452512
rect 235906 452568 235962 452577
rect 235906 452503 235962 452512
rect 238666 452568 238722 452577
rect 238666 452503 238722 452512
rect 241426 452568 241482 452577
rect 241426 452503 241482 452512
rect 243174 452568 243230 452577
rect 243174 452503 243230 452512
rect 245566 452568 245622 452577
rect 245566 452503 245622 452512
rect 253846 452568 253902 452577
rect 253846 452503 253902 452512
rect 255686 452568 255742 452577
rect 255686 452503 255742 452512
rect 260746 452568 260802 452577
rect 260746 452503 260802 452512
rect 263506 452568 263562 452577
rect 263506 452503 263562 452512
rect 265622 452568 265678 452577
rect 265622 452503 265678 452512
rect 269026 452568 269082 452577
rect 269026 452503 269082 452512
rect 271786 452568 271842 452577
rect 271786 452503 271842 452512
rect 273166 452568 273222 452577
rect 273166 452503 273222 452512
rect 275834 452568 275890 452577
rect 275834 452503 275890 452512
rect 213366 452432 213422 452441
rect 213366 452367 213422 452376
rect 213182 451480 213238 451489
rect 213182 451415 213238 451424
rect 203064 450968 203116 450974
rect 203064 450910 203116 450916
rect 203076 419125 203104 450910
rect 204534 447944 204590 447953
rect 204534 447879 204590 447888
rect 204260 447704 204312 447710
rect 204260 447646 204312 447652
rect 204272 419125 204300 447646
rect 204548 447166 204576 447879
rect 213092 447772 213144 447778
rect 213092 447714 213144 447720
rect 205548 447636 205600 447642
rect 205548 447578 205600 447584
rect 204536 447160 204588 447166
rect 204536 447102 204588 447108
rect 205560 419125 205588 447578
rect 206834 445360 206890 445369
rect 206834 445295 206890 445304
rect 206848 419125 206876 445295
rect 208030 445224 208086 445233
rect 208030 445159 208086 445168
rect 208044 419125 208072 445159
rect 209318 445088 209374 445097
rect 209318 445023 209374 445032
rect 209332 419125 209360 445023
rect 211804 444916 211856 444922
rect 211804 444858 211856 444864
rect 210608 444848 210660 444854
rect 210608 444790 210660 444796
rect 210620 419125 210648 444790
rect 211816 419125 211844 444858
rect 213104 419125 213132 447714
rect 213196 420238 213224 451415
rect 213380 422958 213408 452367
rect 214380 448316 214432 448322
rect 214380 448258 214432 448264
rect 213368 422952 213420 422958
rect 213368 422894 213420 422900
rect 213184 420232 213236 420238
rect 213184 420174 213236 420180
rect 214392 419125 214420 448258
rect 215576 448248 215628 448254
rect 215576 448190 215628 448196
rect 215588 419125 215616 448190
rect 216864 448180 216916 448186
rect 216864 448122 216916 448128
rect 216876 419125 216904 448122
rect 219348 448112 219400 448118
rect 219348 448054 219400 448060
rect 218152 448044 218204 448050
rect 218152 447986 218204 447992
rect 218164 419125 218192 447986
rect 219360 419125 219388 448054
rect 220636 447976 220688 447982
rect 220636 447918 220688 447924
rect 220648 419125 220676 447918
rect 221924 447908 221976 447914
rect 221924 447850 221976 447856
rect 221936 419125 221964 447850
rect 223120 447840 223172 447846
rect 223120 447782 223172 447788
rect 223132 419125 223160 447782
rect 226892 445732 226944 445738
rect 226892 445674 226944 445680
rect 225696 445664 225748 445670
rect 225696 445606 225748 445612
rect 224408 444984 224460 444990
rect 224408 444926 224460 444932
rect 224420 419125 224448 444926
rect 225708 419125 225736 445606
rect 226904 419125 226932 445674
rect 228180 445596 228232 445602
rect 228180 445538 228232 445544
rect 228192 419125 228220 445538
rect 230664 445528 230716 445534
rect 230664 445470 230716 445476
rect 229468 445392 229520 445398
rect 229468 445334 229520 445340
rect 229480 419125 229508 445334
rect 230676 419125 230704 445470
rect 231780 424386 231808 452503
rect 231952 445460 232004 445466
rect 231952 445402 232004 445408
rect 231768 424380 231820 424386
rect 231768 424322 231820 424328
rect 231964 419125 231992 445402
rect 234436 445324 234488 445330
rect 234436 445266 234488 445272
rect 233240 445256 233292 445262
rect 233240 445198 233292 445204
rect 233252 419125 233280 445198
rect 234448 419125 234476 445266
rect 234540 442270 234568 452503
rect 235724 445188 235776 445194
rect 235724 445130 235776 445136
rect 234528 442264 234580 442270
rect 234528 442206 234580 442212
rect 235736 419125 235764 445130
rect 235920 424454 235948 452503
rect 237012 445120 237064 445126
rect 237012 445062 237064 445068
rect 235908 424448 235960 424454
rect 235908 424390 235960 424396
rect 237024 419125 237052 445062
rect 238208 445052 238260 445058
rect 238208 444994 238260 445000
rect 238220 419125 238248 444994
rect 238680 424522 238708 452503
rect 240782 447808 240838 447817
rect 240782 447743 240838 447752
rect 239496 442400 239548 442406
rect 239496 442342 239548 442348
rect 238668 424516 238720 424522
rect 238668 424458 238720 424464
rect 239508 419125 239536 442342
rect 240796 419125 240824 447743
rect 241440 424590 241468 452503
rect 243188 449206 243216 452503
rect 243176 449200 243228 449206
rect 243176 449142 243228 449148
rect 244556 446616 244608 446622
rect 244556 446558 244608 446564
rect 243268 445120 243320 445126
rect 243268 445062 243320 445068
rect 241980 431520 242032 431526
rect 241980 431462 242032 431468
rect 241428 424584 241480 424590
rect 241428 424526 241480 424532
rect 241992 419125 242020 431462
rect 243280 419125 243308 445062
rect 244568 419125 244596 446558
rect 245580 432614 245608 452503
rect 248234 451344 248290 451353
rect 248234 451279 248290 451288
rect 251086 451344 251142 451353
rect 251086 451279 251142 451288
rect 247040 449472 247092 449478
rect 247040 449414 247092 449420
rect 245568 432608 245620 432614
rect 245568 432550 245620 432556
rect 245752 423088 245804 423094
rect 245752 423030 245804 423036
rect 245764 419125 245792 423030
rect 247052 419125 247080 449414
rect 248248 436762 248276 451279
rect 249522 447944 249578 447953
rect 249522 447879 249578 447888
rect 248326 439512 248382 439521
rect 248326 439447 248382 439456
rect 248236 436756 248288 436762
rect 248236 436698 248288 436704
rect 248340 419125 248368 439447
rect 249536 419125 249564 447879
rect 250810 447672 250866 447681
rect 250810 447607 250866 447616
rect 250824 419125 250852 447607
rect 251100 435402 251128 451279
rect 252100 447976 252152 447982
rect 252100 447918 252152 447924
rect 251088 435396 251140 435402
rect 251088 435338 251140 435344
rect 252112 419125 252140 447918
rect 253296 445392 253348 445398
rect 253296 445334 253348 445340
rect 253308 419125 253336 445334
rect 253860 434042 253888 452503
rect 255700 447846 255728 452503
rect 259366 451344 259422 451353
rect 259366 451279 259422 451288
rect 255688 447840 255740 447846
rect 255688 447782 255740 447788
rect 258356 445460 258408 445466
rect 258356 445402 258408 445408
rect 254584 445324 254636 445330
rect 254584 445266 254636 445272
rect 253848 434036 253900 434042
rect 253848 433978 253900 433984
rect 254596 419125 254624 445266
rect 257068 445256 257120 445262
rect 257068 445198 257120 445204
rect 255872 445188 255924 445194
rect 255872 445130 255924 445136
rect 255884 419125 255912 445130
rect 257080 419125 257108 445198
rect 258368 419125 258396 445402
rect 259380 431458 259408 451279
rect 259644 445528 259696 445534
rect 259644 445470 259696 445476
rect 259368 431452 259420 431458
rect 259368 431394 259420 431400
rect 259656 419125 259684 445470
rect 260760 440978 260788 452503
rect 262128 445664 262180 445670
rect 262128 445606 262180 445612
rect 260840 445596 260892 445602
rect 260840 445538 260892 445544
rect 260748 440972 260800 440978
rect 260748 440914 260800 440920
rect 260852 419125 260880 445538
rect 262140 419125 262168 445606
rect 263520 443766 263548 452503
rect 264612 448180 264664 448186
rect 264612 448122 264664 448128
rect 263508 443760 263560 443766
rect 263508 443702 263560 443708
rect 263416 442604 263468 442610
rect 263416 442546 263468 442552
rect 263428 419125 263456 442546
rect 264624 419125 264652 448122
rect 265636 445058 265664 452503
rect 268384 445732 268436 445738
rect 268384 445674 268436 445680
rect 265624 445052 265676 445058
rect 265624 444994 265676 445000
rect 267188 442536 267240 442542
rect 267188 442478 267240 442484
rect 265900 442468 265952 442474
rect 265900 442410 265952 442416
rect 265912 419125 265940 442410
rect 267200 419125 267228 442478
rect 268396 419125 268424 445674
rect 269040 422958 269068 452503
rect 269672 444984 269724 444990
rect 269672 444926 269724 444932
rect 269028 422952 269080 422958
rect 269028 422894 269080 422900
rect 269684 419125 269712 444926
rect 270960 444848 271012 444854
rect 270960 444790 271012 444796
rect 270972 419125 271000 444790
rect 271800 423026 271828 452503
rect 273180 446486 273208 452503
rect 273168 446480 273220 446486
rect 273168 446422 273220 446428
rect 274732 442808 274784 442814
rect 274732 442750 274784 442756
rect 273444 442740 273496 442746
rect 273444 442682 273496 442688
rect 272156 442672 272208 442678
rect 272156 442614 272208 442620
rect 271788 423020 271840 423026
rect 271788 422962 271840 422968
rect 272168 419125 272196 442614
rect 273456 419125 273484 442682
rect 274744 419125 274772 442750
rect 275848 438258 275876 452503
rect 278056 452130 278084 453494
rect 281448 453484 281500 453490
rect 281448 453426 281500 453432
rect 278686 452568 278742 452577
rect 278686 452503 278742 452512
rect 280158 452568 280214 452577
rect 280158 452503 280214 452512
rect 278044 452124 278096 452130
rect 278044 452066 278096 452072
rect 277216 442944 277268 442950
rect 277216 442886 277268 442892
rect 275928 442876 275980 442882
rect 275928 442818 275980 442824
rect 275836 438252 275888 438258
rect 275836 438194 275888 438200
rect 275940 419125 275968 442818
rect 277228 419125 277256 442886
rect 278700 442406 278728 452503
rect 280172 449342 280200 452503
rect 281460 452169 281488 453426
rect 284312 453150 284340 453591
rect 284300 453144 284352 453150
rect 284300 453086 284352 453092
rect 286796 453014 286824 453591
rect 288912 453354 288940 453727
rect 294786 453727 294842 453736
rect 291016 453698 291068 453704
rect 289820 453688 289872 453694
rect 289820 453630 289872 453636
rect 290186 453656 290242 453665
rect 288900 453348 288952 453354
rect 288900 453290 288952 453296
rect 286784 453008 286836 453014
rect 286784 452950 286836 452956
rect 282090 452568 282146 452577
rect 282090 452503 282146 452512
rect 284206 452568 284262 452577
rect 284206 452503 284262 452512
rect 285586 452568 285642 452577
rect 285586 452503 285642 452512
rect 288346 452568 288402 452577
rect 288346 452503 288402 452512
rect 282104 452266 282132 452503
rect 283194 452296 283250 452305
rect 282092 452260 282144 452266
rect 283194 452231 283250 452240
rect 282092 452202 282144 452208
rect 283208 452198 283236 452231
rect 283196 452192 283248 452198
rect 281446 452160 281502 452169
rect 283196 452134 283248 452140
rect 281446 452095 281502 452104
rect 280988 451852 281040 451858
rect 280988 451794 281040 451800
rect 280160 449336 280212 449342
rect 280160 449278 280212 449284
rect 278688 442400 278740 442406
rect 278688 442342 278740 442348
rect 278504 442196 278556 442202
rect 278504 442138 278556 442144
rect 278516 419125 278544 442138
rect 279700 442128 279752 442134
rect 279700 442070 279752 442076
rect 279712 419125 279740 442070
rect 281000 419125 281028 451794
rect 282276 451784 282328 451790
rect 282276 451726 282328 451732
rect 282288 419125 282316 451726
rect 283472 451716 283524 451722
rect 283472 451658 283524 451664
rect 283484 419125 283512 451658
rect 284220 436830 284248 452503
rect 285600 441046 285628 452503
rect 285588 441040 285640 441046
rect 285588 440982 285640 440988
rect 288360 438326 288388 452503
rect 288348 438320 288400 438326
rect 288348 438262 288400 438268
rect 284208 436824 284260 436830
rect 284208 436766 284260 436772
rect 288532 424992 288584 424998
rect 288532 424934 288584 424940
rect 287244 424924 287296 424930
rect 287244 424866 287296 424872
rect 286048 424856 286100 424862
rect 286048 424798 286100 424804
rect 284760 421864 284812 421870
rect 284760 421806 284812 421812
rect 284772 419125 284800 421806
rect 286060 419125 286088 424798
rect 287256 419125 287284 424866
rect 288544 419125 288572 424934
rect 289832 419125 289860 453630
rect 290186 453591 290242 453600
rect 290200 452878 290228 453591
rect 290188 452872 290240 452878
rect 290188 452814 290240 452820
rect 291028 419125 291056 453698
rect 291198 453656 291254 453665
rect 291198 453591 291254 453600
rect 293682 453656 293738 453665
rect 293682 453591 293738 453600
rect 291212 452810 291240 453591
rect 293696 452946 293724 453591
rect 294800 453422 294828 453727
rect 297086 453656 297142 453665
rect 297086 453591 297142 453600
rect 298466 453656 298522 453665
rect 298466 453591 298522 453600
rect 299570 453656 299626 453665
rect 299570 453591 299626 453600
rect 311070 453656 311126 453665
rect 311070 453591 311126 453600
rect 312358 453656 312414 453665
rect 312358 453591 312414 453600
rect 324964 453620 325016 453626
rect 294788 453416 294840 453422
rect 294788 453358 294840 453364
rect 293684 452940 293736 452946
rect 293684 452882 293736 452888
rect 291200 452804 291252 452810
rect 291200 452746 291252 452752
rect 292580 452736 292632 452742
rect 297100 452713 297128 453591
rect 298480 453286 298508 453591
rect 298560 453416 298612 453422
rect 298560 453358 298612 453364
rect 298468 453280 298520 453286
rect 298468 453222 298520 453228
rect 292580 452678 292632 452684
rect 297086 452704 297142 452713
rect 292592 452577 292620 452678
rect 297086 452639 297142 452648
rect 291106 452568 291162 452577
rect 291106 452503 291162 452512
rect 292578 452568 292634 452577
rect 292578 452503 292634 452512
rect 293038 452568 293094 452577
rect 293038 452503 293094 452512
rect 296626 452568 296682 452577
rect 296626 452503 296682 452512
rect 291120 430234 291148 452503
rect 293052 446554 293080 452503
rect 294786 452024 294842 452033
rect 294786 451959 294842 451968
rect 293590 451888 293646 451897
rect 293590 451823 293646 451832
rect 293040 446548 293092 446554
rect 293040 446490 293092 446496
rect 292304 432676 292356 432682
rect 292304 432618 292356 432624
rect 291108 430228 291160 430234
rect 291108 430170 291160 430176
rect 292316 419125 292344 432618
rect 293604 419125 293632 451823
rect 294800 419125 294828 451959
rect 296076 447908 296128 447914
rect 296076 447850 296128 447856
rect 296088 419125 296116 447850
rect 296640 424658 296668 452503
rect 297362 452160 297418 452169
rect 297362 452095 297418 452104
rect 296628 424652 296680 424658
rect 296628 424594 296680 424600
rect 297376 419125 297404 452095
rect 298572 419125 298600 453358
rect 299584 453218 299612 453591
rect 301228 453484 301280 453490
rect 301228 453426 301280 453432
rect 299848 453348 299900 453354
rect 299848 453290 299900 453296
rect 299572 453212 299624 453218
rect 299572 453154 299624 453160
rect 299386 452568 299442 452577
rect 299386 452503 299442 452512
rect 299400 424726 299428 452503
rect 299388 424720 299440 424726
rect 299388 424662 299440 424668
rect 299860 419125 299888 453290
rect 300766 452568 300822 452577
rect 300766 452503 300822 452512
rect 300122 452296 300178 452305
rect 300122 452231 300178 452240
rect 300136 449750 300164 452231
rect 300124 449744 300176 449750
rect 300124 449686 300176 449692
rect 300780 424794 300808 452503
rect 301240 431954 301268 453426
rect 311084 453082 311112 453591
rect 311164 453552 311216 453558
rect 311164 453494 311216 453500
rect 311072 453076 311124 453082
rect 311072 453018 311124 453024
rect 305276 452600 305328 452606
rect 301962 452568 302018 452577
rect 301962 452503 302018 452512
rect 303066 452568 303122 452577
rect 303066 452503 303122 452512
rect 304170 452568 304226 452577
rect 304170 452503 304226 452512
rect 305274 452568 305276 452577
rect 305328 452568 305330 452577
rect 305274 452503 305330 452512
rect 306378 452568 306434 452577
rect 306378 452503 306434 452512
rect 307850 452568 307906 452577
rect 307850 452503 307906 452512
rect 308954 452568 309010 452577
rect 308954 452503 309010 452512
rect 309874 452568 309930 452577
rect 309874 452503 309930 452512
rect 301976 452130 302004 452503
rect 301964 452124 302016 452130
rect 301964 452066 302016 452072
rect 302332 451988 302384 451994
rect 302332 451930 302384 451936
rect 301148 431926 301268 431954
rect 300768 424788 300820 424794
rect 300768 424730 300820 424736
rect 301148 419125 301176 431926
rect 302344 419125 302372 451930
rect 303080 451518 303108 452503
rect 304184 452334 304212 452503
rect 304172 452328 304224 452334
rect 303526 452296 303582 452305
rect 304172 452270 304224 452276
rect 306286 452296 306342 452305
rect 303526 452231 303582 452240
rect 306286 452231 306342 452240
rect 303068 451512 303120 451518
rect 303068 451454 303120 451460
rect 303540 428738 303568 452231
rect 306104 452124 306156 452130
rect 306104 452066 306156 452072
rect 303620 452056 303672 452062
rect 303620 451998 303672 452004
rect 303528 428732 303580 428738
rect 303528 428674 303580 428680
rect 303632 419125 303660 451998
rect 304908 427168 304960 427174
rect 304908 427110 304960 427116
rect 304920 419125 304948 427110
rect 306116 419125 306144 452066
rect 306300 439618 306328 452231
rect 306392 451382 306420 452503
rect 307864 452402 307892 452503
rect 307852 452396 307904 452402
rect 307852 452338 307904 452344
rect 308680 452192 308732 452198
rect 308680 452134 308732 452140
rect 306380 451376 306432 451382
rect 306380 451318 306432 451324
rect 307390 445088 307446 445097
rect 307390 445023 307446 445032
rect 306288 439612 306340 439618
rect 306288 439554 306340 439560
rect 307404 419125 307432 445023
rect 308692 419125 308720 452134
rect 308968 451450 308996 452503
rect 309888 451926 309916 452503
rect 309968 452260 310020 452266
rect 309968 452202 310020 452208
rect 309876 451920 309928 451926
rect 309876 451862 309928 451868
rect 308956 451444 309008 451450
rect 308956 451386 309008 451392
rect 309046 451344 309102 451353
rect 309046 451279 309102 451288
rect 309060 435470 309088 451279
rect 309048 435464 309100 435470
rect 309048 435406 309100 435412
rect 309980 431954 310008 452202
rect 309888 431926 310008 431954
rect 309888 419125 309916 431926
rect 311176 419125 311204 453494
rect 312372 452674 312400 453591
rect 324964 453562 325016 453568
rect 312360 452668 312412 452674
rect 312360 452610 312412 452616
rect 313370 452568 313426 452577
rect 313370 452503 313372 452512
rect 313424 452503 313426 452512
rect 314658 452568 314714 452577
rect 314658 452503 314714 452512
rect 320178 452568 320234 452577
rect 320178 452503 320234 452512
rect 313372 452474 313424 452480
rect 314672 452470 314700 452503
rect 314660 452464 314712 452470
rect 314660 452406 314712 452412
rect 317420 452464 317472 452470
rect 317420 452406 317472 452412
rect 316224 452396 316276 452402
rect 316224 452338 316276 452344
rect 312452 452328 312504 452334
rect 312452 452270 312504 452276
rect 312464 419125 312492 452270
rect 314936 436892 314988 436898
rect 314936 436834 314988 436840
rect 313648 425740 313700 425746
rect 313648 425682 313700 425688
rect 313660 419125 313688 425682
rect 314948 419125 314976 436834
rect 316236 419125 316264 452338
rect 317432 419125 317460 452406
rect 319442 452296 319498 452305
rect 319442 452231 319498 452240
rect 319456 451382 319484 452231
rect 320192 451926 320220 452503
rect 320180 451920 320232 451926
rect 320180 451862 320232 451868
rect 318800 451376 318852 451382
rect 318800 451318 318852 451324
rect 319444 451376 319496 451382
rect 319444 451318 319496 451324
rect 318812 449818 318840 451318
rect 320192 451314 320220 451862
rect 320180 451308 320232 451314
rect 320180 451250 320232 451256
rect 318800 449812 318852 449818
rect 318800 449754 318852 449760
rect 322480 448112 322532 448118
rect 322480 448054 322532 448060
rect 319996 448044 320048 448050
rect 319996 447986 320048 447992
rect 318708 425808 318760 425814
rect 318708 425750 318760 425756
rect 318720 419125 318748 425750
rect 320008 419125 320036 447986
rect 321192 425876 321244 425882
rect 321192 425818 321244 425824
rect 321204 419125 321232 425818
rect 322492 419125 322520 448054
rect 323768 430296 323820 430302
rect 323768 430238 323820 430244
rect 323780 419125 323808 430238
rect 324976 419125 325004 453562
rect 335084 452736 335136 452742
rect 335084 452678 335136 452684
rect 330024 452532 330076 452538
rect 330024 452474 330076 452480
rect 327540 444916 327592 444922
rect 327540 444858 327592 444864
rect 326252 432744 326304 432750
rect 326252 432686 326304 432692
rect 326264 419125 326292 432686
rect 327552 419125 327580 444858
rect 328736 425944 328788 425950
rect 328736 425886 328788 425892
rect 328748 419125 328776 425886
rect 330036 419125 330064 452474
rect 333796 439816 333848 439822
rect 333796 439758 333848 439764
rect 331312 431588 331364 431594
rect 331312 431530 331364 431536
rect 331324 419125 331352 431530
rect 332508 425060 332560 425066
rect 332508 425002 332560 425008
rect 332520 419125 332548 425002
rect 333808 419125 333836 439758
rect 335096 419125 335124 452678
rect 336292 419125 336320 453834
rect 336752 431526 336780 603735
rect 336922 585304 336978 585313
rect 336922 585239 336978 585248
rect 336832 574864 336884 574870
rect 336832 574806 336884 574812
rect 336844 442610 336872 574806
rect 336936 453898 336964 585239
rect 337120 575482 337148 659670
rect 340142 659631 340198 659640
rect 339406 612232 339462 612241
rect 339406 612167 339462 612176
rect 339420 612066 339448 612167
rect 339408 612060 339460 612066
rect 339408 612002 339460 612008
rect 339406 611008 339462 611017
rect 339406 610943 339462 610952
rect 339420 610638 339448 610943
rect 339408 610632 339460 610638
rect 339408 610574 339460 610580
rect 338302 609240 338358 609249
rect 338302 609175 338358 609184
rect 338316 608666 338344 609175
rect 338304 608660 338356 608666
rect 338304 608602 338356 608608
rect 338118 608152 338174 608161
rect 338118 608087 338174 608096
rect 338132 607238 338160 608087
rect 338120 607232 338172 607238
rect 338120 607174 338172 607180
rect 337382 583672 337438 583681
rect 337382 583607 337438 583616
rect 337108 575476 337160 575482
rect 337108 575418 337160 575424
rect 337014 574288 337070 574297
rect 337014 574223 337070 574232
rect 336924 453892 336976 453898
rect 336924 453834 336976 453840
rect 337028 445398 337056 574223
rect 337120 574161 337148 575418
rect 337106 574152 337162 574161
rect 337106 574087 337162 574096
rect 337108 572688 337160 572694
rect 337108 572630 337160 572636
rect 337016 445392 337068 445398
rect 337016 445334 337068 445340
rect 337120 442950 337148 572630
rect 337200 572620 337252 572626
rect 337200 572562 337252 572568
rect 337108 442944 337160 442950
rect 337108 442886 337160 442892
rect 336832 442604 336884 442610
rect 336832 442546 336884 442552
rect 337212 442202 337240 572562
rect 337292 572552 337344 572558
rect 337292 572494 337344 572500
rect 337200 442196 337252 442202
rect 337200 442138 337252 442144
rect 337304 442134 337332 572494
rect 337396 452742 337424 583607
rect 338028 575544 338080 575550
rect 338028 575486 338080 575492
rect 338040 575385 338068 575486
rect 338026 575376 338082 575385
rect 338026 575311 338082 575320
rect 337566 575240 337622 575249
rect 337566 575175 337622 575184
rect 337476 574592 337528 574598
rect 337476 574534 337528 574540
rect 337384 452736 337436 452742
rect 337384 452678 337436 452684
rect 337488 448186 337516 574534
rect 337476 448180 337528 448186
rect 337476 448122 337528 448128
rect 337580 447982 337608 575175
rect 337568 447976 337620 447982
rect 337568 447918 337620 447924
rect 337292 442128 337344 442134
rect 337292 442070 337344 442076
rect 336740 431520 336792 431526
rect 336740 431462 336792 431468
rect 338132 423094 338160 607174
rect 338212 604512 338264 604518
rect 338212 604454 338264 604460
rect 338224 445126 338252 604454
rect 338316 449478 338344 608602
rect 338394 606520 338450 606529
rect 338394 606455 338450 606464
rect 338408 605878 338436 606455
rect 338396 605872 338448 605878
rect 338396 605814 338448 605820
rect 338304 449472 338356 449478
rect 338304 449414 338356 449420
rect 338408 446622 338436 605814
rect 339406 605568 339462 605577
rect 339406 605503 339462 605512
rect 339420 604518 339448 605503
rect 339408 604512 339460 604518
rect 339408 604454 339460 604460
rect 339222 603800 339278 603809
rect 339222 603735 339224 603744
rect 339276 603735 339278 603744
rect 339224 603706 339276 603712
rect 339224 585812 339276 585818
rect 339224 585754 339276 585760
rect 339236 585313 339264 585754
rect 339222 585304 339278 585313
rect 339222 585239 339278 585248
rect 339406 583672 339462 583681
rect 339406 583607 339462 583616
rect 339420 583030 339448 583607
rect 339408 583024 339460 583030
rect 339408 582966 339460 582972
rect 338486 575104 338542 575113
rect 338486 575039 338542 575048
rect 342352 575068 342404 575074
rect 338396 446616 338448 446622
rect 338396 446558 338448 446564
rect 338500 445330 338528 575039
rect 342352 575010 342404 575016
rect 340144 575000 340196 575006
rect 340144 574942 340196 574948
rect 341246 574968 341302 574977
rect 339592 574932 339644 574938
rect 339592 574874 339644 574880
rect 339500 574252 339552 574258
rect 339500 574194 339552 574200
rect 338580 571940 338632 571946
rect 338580 571882 338632 571888
rect 338488 445324 338540 445330
rect 338488 445266 338540 445272
rect 338212 445120 338264 445126
rect 338212 445062 338264 445068
rect 338592 442814 338620 571882
rect 338764 540456 338816 540462
rect 338764 540398 338816 540404
rect 338672 540388 338724 540394
rect 338672 540330 338724 540336
rect 338684 453762 338712 540330
rect 338672 453756 338724 453762
rect 338672 453698 338724 453704
rect 338776 453694 338804 540398
rect 338856 539844 338908 539850
rect 338856 539786 338908 539792
rect 338868 487150 338896 539786
rect 339316 491292 339368 491298
rect 339316 491234 339368 491240
rect 339328 489977 339356 491234
rect 339408 491224 339460 491230
rect 339408 491166 339460 491172
rect 339420 490929 339448 491166
rect 339406 490920 339462 490929
rect 339406 490855 339462 490864
rect 339314 489968 339370 489977
rect 339314 489903 339370 489912
rect 338856 487144 338908 487150
rect 338856 487086 338908 487092
rect 338868 486849 338896 487086
rect 338854 486840 338910 486849
rect 338854 486775 338910 486784
rect 339406 485072 339462 485081
rect 339406 485007 339462 485016
rect 339420 484430 339448 485007
rect 339408 484424 339460 484430
rect 339408 484366 339460 484372
rect 338854 482216 338910 482225
rect 338854 482151 338910 482160
rect 338868 481710 338896 482151
rect 338856 481704 338908 481710
rect 338856 481646 338908 481652
rect 338764 453688 338816 453694
rect 338764 453630 338816 453636
rect 338868 449410 338896 481646
rect 339406 463992 339462 464001
rect 339406 463927 339462 463936
rect 339420 463758 339448 463927
rect 339408 463752 339460 463758
rect 339408 463694 339460 463700
rect 339132 463004 339184 463010
rect 339132 462946 339184 462952
rect 339144 462369 339172 462946
rect 339130 462360 339186 462369
rect 339130 462295 339186 462304
rect 339040 461644 339092 461650
rect 339040 461586 339092 461592
rect 339052 461553 339080 461586
rect 339038 461544 339094 461553
rect 339038 461479 339094 461488
rect 339144 451274 339172 462295
rect 339052 451246 339172 451274
rect 338856 449404 338908 449410
rect 338856 449346 338908 449352
rect 339052 448390 339080 451246
rect 339040 448384 339092 448390
rect 339040 448326 339092 448332
rect 339512 442882 339540 574194
rect 339604 445534 339632 574874
rect 339684 574796 339736 574802
rect 339684 574738 339736 574744
rect 339696 445670 339724 574738
rect 339776 574728 339828 574734
rect 339776 574670 339828 574676
rect 339684 445664 339736 445670
rect 339684 445606 339736 445612
rect 339788 445602 339816 574670
rect 339960 574660 340012 574666
rect 339960 574602 340012 574608
rect 339868 571872 339920 571878
rect 339868 571814 339920 571820
rect 339776 445596 339828 445602
rect 339776 445538 339828 445544
rect 339592 445528 339644 445534
rect 339592 445470 339644 445476
rect 339500 442876 339552 442882
rect 339500 442818 339552 442824
rect 338580 442808 338632 442814
rect 338580 442750 338632 442756
rect 339880 442746 339908 571814
rect 339972 451722 340000 574602
rect 340052 539776 340104 539782
rect 340052 539718 340104 539724
rect 340064 488510 340092 539718
rect 340052 488504 340104 488510
rect 340052 488446 340104 488452
rect 340064 487801 340092 488446
rect 340050 487792 340106 487801
rect 340050 487727 340106 487736
rect 340050 483984 340106 483993
rect 340050 483919 340106 483928
rect 340064 483070 340092 483919
rect 340052 483064 340104 483070
rect 340052 483006 340104 483012
rect 339960 451716 340012 451722
rect 339960 451658 340012 451664
rect 340064 449886 340092 483006
rect 340052 449880 340104 449886
rect 340052 449822 340104 449828
rect 339868 442740 339920 442746
rect 339868 442682 339920 442688
rect 340156 431594 340184 574942
rect 341246 574903 341302 574912
rect 341062 574832 341118 574841
rect 341062 574767 341118 574776
rect 340972 574388 341024 574394
rect 340972 574330 341024 574336
rect 340880 572484 340932 572490
rect 340880 572426 340932 572432
rect 340328 539708 340380 539714
rect 340328 539650 340380 539656
rect 340236 539640 340288 539646
rect 340236 539582 340288 539588
rect 340248 491230 340276 539582
rect 340340 491298 340368 539650
rect 340328 491292 340380 491298
rect 340328 491234 340380 491240
rect 340236 491224 340288 491230
rect 340236 491166 340288 491172
rect 340236 484424 340288 484430
rect 340236 484366 340288 484372
rect 340248 451110 340276 484366
rect 340328 463752 340380 463758
rect 340328 463694 340380 463700
rect 340236 451104 340288 451110
rect 340236 451046 340288 451052
rect 340340 448458 340368 463694
rect 340328 448452 340380 448458
rect 340328 448394 340380 448400
rect 340892 442678 340920 572426
rect 340984 444854 341012 574330
rect 341076 445262 341104 574767
rect 341154 574696 341210 574705
rect 341154 574631 341210 574640
rect 341168 445466 341196 574631
rect 341156 445460 341208 445466
rect 341156 445402 341208 445408
rect 341064 445256 341116 445262
rect 341064 445198 341116 445204
rect 341260 445194 341288 574903
rect 341432 574524 341484 574530
rect 341432 574466 341484 574472
rect 341340 572416 341392 572422
rect 341340 572358 341392 572364
rect 341352 445738 341380 572358
rect 341444 451858 341472 574466
rect 342260 574320 342312 574326
rect 342260 574262 342312 574268
rect 341524 574184 341576 574190
rect 341524 574126 341576 574132
rect 341432 451852 341484 451858
rect 341432 451794 341484 451800
rect 341536 451790 341564 574126
rect 341614 543144 341670 543153
rect 341614 543079 341670 543088
rect 341628 543046 341656 543079
rect 341616 543040 341668 543046
rect 341616 542982 341668 542988
rect 341708 538892 341760 538898
rect 341708 538834 341760 538840
rect 341524 451784 341576 451790
rect 341524 451726 341576 451732
rect 341522 450936 341578 450945
rect 341522 450871 341578 450880
rect 341340 445732 341392 445738
rect 341340 445674 341392 445680
rect 341248 445188 341300 445194
rect 341248 445130 341300 445136
rect 340972 444848 341024 444854
rect 340972 444790 341024 444796
rect 340880 442672 340932 442678
rect 340880 442614 340932 442620
rect 340144 431588 340196 431594
rect 340144 431530 340196 431536
rect 338120 423088 338172 423094
rect 338120 423030 338172 423036
rect 337382 421832 337438 421841
rect 337382 421767 337438 421776
rect 338854 421832 338910 421841
rect 338854 421767 338910 421776
rect 340050 421832 340106 421841
rect 341536 421802 341564 450871
rect 341614 428088 341670 428097
rect 341614 428023 341670 428032
rect 340050 421767 340106 421776
rect 341524 421796 341576 421802
rect 337396 419139 337424 421767
rect 337396 419111 337586 419139
rect 338868 419125 338896 421767
rect 340064 419125 340092 421767
rect 341524 421738 341576 421744
rect 341628 419139 341656 428023
rect 341720 424998 341748 538834
rect 341708 424992 341760 424998
rect 341708 424934 341760 424940
rect 342272 421870 342300 574262
rect 342364 442474 342392 575010
rect 342444 574456 342496 574462
rect 342444 574398 342496 574404
rect 342456 442542 342484 574398
rect 342536 572280 342588 572286
rect 342536 572222 342588 572228
rect 342548 444990 342576 572222
rect 343824 545080 343876 545086
rect 343824 545022 343876 545028
rect 342628 544400 342680 544406
rect 342628 544342 342680 544348
rect 342640 543726 342668 544342
rect 342628 543720 342680 543726
rect 342628 543662 342680 543668
rect 342536 444984 342588 444990
rect 342536 444926 342588 444932
rect 342444 442536 342496 442542
rect 342444 442478 342496 442484
rect 342352 442468 342404 442474
rect 342352 442410 342404 442416
rect 342260 421864 342312 421870
rect 342260 421806 342312 421812
rect 341366 419111 341656 419139
rect 342640 419125 342668 543662
rect 342720 539096 342772 539102
rect 342720 539038 342772 539044
rect 342732 425066 342760 539038
rect 342812 539028 342864 539034
rect 342812 538970 342864 538976
rect 342720 425060 342772 425066
rect 342720 425002 342772 425008
rect 342824 424862 342852 538970
rect 342904 538960 342956 538966
rect 342904 538902 342956 538908
rect 342916 424930 342944 538902
rect 342904 424924 342956 424930
rect 342904 424866 342956 424872
rect 342812 424856 342864 424862
rect 342812 424798 342864 424804
rect 343836 419125 343864 545022
rect 344296 445126 344324 700606
rect 351184 700528 351236 700534
rect 351184 700470 351236 700476
rect 348424 700392 348476 700398
rect 348424 700334 348476 700340
rect 344376 570648 344428 570654
rect 344376 570590 344428 570596
rect 344388 545086 344416 570590
rect 347044 569220 347096 569226
rect 347044 569162 347096 569168
rect 347056 547874 347084 569162
rect 347136 567860 347188 567866
rect 347136 567802 347188 567808
rect 347148 549234 347176 567802
rect 347136 549228 347188 549234
rect 347136 549170 347188 549176
rect 347596 549228 347648 549234
rect 347596 549170 347648 549176
rect 347044 547868 347096 547874
rect 347044 547810 347096 547816
rect 347056 546514 347084 547810
rect 346400 546508 346452 546514
rect 346400 546450 346452 546456
rect 347044 546508 347096 546514
rect 347044 546450 347096 546456
rect 345112 545760 345164 545766
rect 345112 545702 345164 545708
rect 344376 545080 344428 545086
rect 344376 545022 344428 545028
rect 344284 445120 344336 445126
rect 344284 445062 344336 445068
rect 345124 419125 345152 545702
rect 346412 419125 346440 546450
rect 347608 419125 347636 549170
rect 348436 443834 348464 700334
rect 348516 562352 348568 562358
rect 348516 562294 348568 562300
rect 348528 550594 348556 562294
rect 348516 550588 348568 550594
rect 348516 550530 348568 550536
rect 348528 547874 348556 550530
rect 348528 547846 348924 547874
rect 348424 443828 348476 443834
rect 348424 443770 348476 443776
rect 348896 419125 348924 547846
rect 350172 539028 350224 539034
rect 350172 538970 350224 538976
rect 350184 419125 350212 538970
rect 351196 447982 351224 700470
rect 353944 700324 353996 700330
rect 353944 700266 353996 700272
rect 351368 562352 351420 562358
rect 351368 562294 351420 562300
rect 351184 447976 351236 447982
rect 351184 447918 351236 447924
rect 351380 419125 351408 562294
rect 352656 540524 352708 540530
rect 352656 540466 352708 540472
rect 352668 419125 352696 540466
rect 353300 540388 353352 540394
rect 353300 540330 353352 540336
rect 353312 441614 353340 540330
rect 353312 441586 353616 441614
rect 353588 419139 353616 441586
rect 353956 431526 353984 700266
rect 356428 566500 356480 566506
rect 356428 566442 356480 566448
rect 355140 556844 355192 556850
rect 355140 556786 355192 556792
rect 353944 431520 353996 431526
rect 353944 431462 353996 431468
rect 353588 419111 353962 419139
rect 355152 419125 355180 556786
rect 356440 419125 356468 566442
rect 356716 439754 356744 700674
rect 358084 700460 358136 700466
rect 358084 700402 358136 700408
rect 357716 563780 357768 563786
rect 357716 563722 357768 563728
rect 356704 439748 356756 439754
rect 356704 439690 356756 439696
rect 357728 419125 357756 563722
rect 358096 441114 358124 700402
rect 364996 700330 365024 703520
rect 396724 700664 396776 700670
rect 396724 700606 396776 700612
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 393964 700324 394016 700330
rect 393964 700266 394016 700272
rect 391204 574184 391256 574190
rect 391204 574126 391256 574132
rect 360200 573436 360252 573442
rect 360200 573378 360252 573384
rect 358912 541748 358964 541754
rect 358912 541690 358964 541696
rect 358084 441108 358136 441114
rect 358084 441050 358136 441056
rect 358924 419125 358952 541690
rect 360212 419125 360240 573378
rect 365260 570648 365312 570654
rect 365260 570590 365312 570596
rect 361488 541680 361540 541686
rect 361488 541622 361540 541628
rect 361500 419125 361528 541622
rect 362684 539164 362736 539170
rect 362684 539106 362736 539112
rect 362696 419125 362724 539106
rect 363972 539096 364024 539102
rect 363972 539038 364024 539044
rect 363984 419125 364012 539038
rect 365272 419125 365300 570590
rect 367744 569220 367796 569226
rect 367744 569162 367796 569168
rect 366456 538960 366508 538966
rect 366456 538902 366508 538908
rect 366468 419125 366496 538902
rect 367756 419125 367784 569162
rect 374000 567860 374052 567866
rect 374000 567802 374052 567808
rect 369032 551336 369084 551342
rect 369032 551278 369084 551284
rect 369044 419125 369072 551278
rect 370228 539368 370280 539374
rect 370228 539310 370280 539316
rect 370240 419125 370268 539310
rect 371516 539300 371568 539306
rect 371516 539242 371568 539248
rect 371528 419125 371556 539242
rect 372804 539232 372856 539238
rect 372804 539174 372856 539180
rect 372816 419125 372844 539174
rect 374012 419125 374040 567802
rect 375288 560992 375340 560998
rect 375288 560934 375340 560940
rect 375300 419125 375328 560934
rect 377772 559564 377824 559570
rect 377772 559506 377824 559512
rect 376576 552696 376628 552702
rect 376576 552638 376628 552644
rect 376588 419125 376616 552638
rect 377784 419125 377812 559506
rect 379060 558204 379112 558210
rect 379060 558146 379112 558152
rect 379072 419125 379100 558146
rect 381544 555484 381596 555490
rect 381544 555426 381596 555432
rect 380348 554056 380400 554062
rect 380348 553998 380400 554004
rect 380360 419125 380388 553998
rect 381556 419125 381584 555426
rect 384120 540864 384172 540870
rect 384120 540806 384172 540812
rect 382832 540456 382884 540462
rect 382832 540398 382884 540404
rect 382844 419125 382872 540398
rect 384132 419125 384160 540806
rect 385316 540796 385368 540802
rect 385316 540738 385368 540744
rect 385328 419125 385356 540738
rect 386604 540728 386656 540734
rect 386604 540670 386656 540676
rect 386616 419125 386644 540670
rect 387892 540660 387944 540666
rect 387892 540602 387944 540608
rect 387904 419125 387932 540602
rect 389088 540592 389140 540598
rect 389088 540534 389140 540540
rect 389100 419125 389128 540534
rect 391216 430302 391244 574126
rect 393976 438394 394004 700266
rect 396736 449410 396764 700606
rect 396816 574252 396868 574258
rect 396816 574194 396868 574200
rect 396724 449404 396776 449410
rect 396724 449346 396776 449352
rect 393964 438388 394016 438394
rect 393964 438330 394016 438336
rect 391204 430296 391256 430302
rect 391204 430238 391256 430244
rect 392860 426488 392912 426494
rect 392860 426430 392912 426436
rect 390098 421696 390154 421705
rect 390098 421631 390154 421640
rect 390112 419139 390140 421631
rect 391386 419656 391442 419665
rect 391386 419591 391442 419600
rect 391400 419139 391428 419591
rect 390112 419111 390394 419139
rect 391400 419111 391682 419139
rect 392872 419125 392900 426430
rect 396828 425950 396856 574194
rect 397472 446622 397500 703520
rect 405004 700596 405056 700602
rect 405004 700538 405056 700544
rect 400864 574388 400916 574394
rect 400864 574330 400916 574336
rect 398104 574320 398156 574326
rect 398104 574262 398156 574268
rect 397460 446616 397512 446622
rect 397460 446558 397512 446564
rect 398116 432750 398144 574262
rect 399760 572348 399812 572354
rect 399760 572290 399812 572296
rect 399576 572280 399628 572286
rect 399576 572222 399628 572228
rect 399484 572076 399536 572082
rect 399484 572018 399536 572024
rect 399496 444922 399524 572018
rect 399588 448050 399616 572222
rect 399668 572212 399720 572218
rect 399668 572154 399720 572160
rect 399680 448118 399708 572154
rect 399772 452470 399800 572290
rect 399944 572144 399996 572150
rect 399944 572086 399996 572092
rect 399852 572008 399904 572014
rect 399852 571950 399904 571956
rect 399864 452538 399892 571950
rect 399956 453626 399984 572086
rect 399944 453620 399996 453626
rect 399944 453562 399996 453568
rect 399852 452532 399904 452538
rect 399852 452474 399904 452480
rect 399760 452464 399812 452470
rect 399760 452406 399812 452412
rect 399668 448112 399720 448118
rect 399668 448054 399720 448060
rect 399576 448044 399628 448050
rect 399576 447986 399628 447992
rect 399484 444916 399536 444922
rect 399484 444858 399536 444864
rect 398104 432744 398156 432750
rect 398104 432686 398156 432692
rect 396816 425944 396868 425950
rect 396816 425886 396868 425892
rect 400876 425882 400904 574330
rect 402244 572688 402296 572694
rect 402244 572630 402296 572636
rect 400956 565888 401008 565894
rect 400956 565830 401008 565836
rect 400968 442474 400996 565830
rect 402256 452130 402284 572630
rect 402428 572620 402480 572626
rect 402428 572562 402480 572568
rect 402336 572484 402388 572490
rect 402336 572426 402388 572432
rect 402348 452334 402376 572426
rect 402336 452328 402388 452334
rect 402336 452270 402388 452276
rect 402440 452198 402468 572562
rect 402704 572552 402756 572558
rect 402704 572494 402756 572500
rect 402612 572416 402664 572422
rect 402612 572358 402664 572364
rect 402520 571940 402572 571946
rect 402520 571882 402572 571888
rect 402428 452192 402480 452198
rect 402428 452134 402480 452140
rect 402244 452124 402296 452130
rect 402244 452066 402296 452072
rect 402532 452062 402560 571882
rect 402624 452402 402652 572358
rect 402612 452396 402664 452402
rect 402612 452338 402664 452344
rect 402716 452266 402744 572494
rect 402704 452260 402756 452266
rect 402704 452202 402756 452208
rect 402520 452056 402572 452062
rect 402520 451998 402572 452004
rect 400956 442468 401008 442474
rect 400956 442410 401008 442416
rect 405016 430302 405044 700538
rect 408408 700460 408460 700466
rect 408408 700402 408460 700408
rect 408316 700324 408368 700330
rect 408316 700266 408368 700272
rect 407764 698964 407816 698970
rect 407764 698906 407816 698912
rect 407118 612232 407174 612241
rect 407118 612167 407174 612176
rect 407132 612066 407160 612167
rect 407120 612060 407172 612066
rect 407120 612002 407172 612008
rect 407118 611008 407174 611017
rect 407118 610943 407174 610952
rect 407132 610638 407160 610943
rect 407120 610632 407172 610638
rect 407120 610574 407172 610580
rect 407118 609240 407174 609249
rect 407118 609175 407174 609184
rect 407132 608666 407160 609175
rect 407120 608660 407172 608666
rect 407120 608602 407172 608608
rect 407118 608152 407174 608161
rect 407118 608087 407174 608096
rect 407132 607238 407160 608087
rect 407120 607232 407172 607238
rect 407120 607174 407172 607180
rect 407118 606520 407174 606529
rect 407118 606455 407174 606464
rect 407132 605878 407160 606455
rect 407120 605872 407172 605878
rect 407120 605814 407172 605820
rect 407118 605568 407174 605577
rect 407118 605503 407174 605512
rect 407132 604518 407160 605503
rect 407120 604512 407172 604518
rect 407120 604454 407172 604460
rect 407118 603800 407174 603809
rect 407118 603735 407120 603744
rect 407172 603735 407174 603744
rect 407120 603706 407172 603712
rect 407120 585812 407172 585818
rect 407120 585754 407172 585760
rect 407132 585313 407160 585754
rect 407118 585304 407174 585313
rect 407118 585239 407174 585248
rect 407118 583672 407174 583681
rect 407118 583607 407174 583616
rect 407132 583030 407160 583607
rect 407120 583024 407172 583030
rect 407120 582966 407172 582972
rect 406568 574796 406620 574802
rect 406568 574738 406620 574744
rect 406476 574728 406528 574734
rect 406476 574670 406528 574676
rect 405280 574592 405332 574598
rect 405280 574534 405332 574540
rect 405096 574524 405148 574530
rect 405096 574466 405148 574472
rect 405004 430296 405056 430302
rect 405004 430238 405056 430244
rect 400864 425876 400916 425882
rect 400864 425818 400916 425824
rect 405108 425746 405136 574466
rect 405186 572248 405242 572257
rect 405186 572183 405242 572192
rect 405200 447914 405228 572183
rect 405292 453558 405320 574534
rect 406384 574456 406436 574462
rect 406384 574398 406436 574404
rect 405554 572384 405610 572393
rect 405554 572319 405610 572328
rect 405370 572112 405426 572121
rect 405370 572047 405426 572056
rect 405280 453552 405332 453558
rect 405280 453494 405332 453500
rect 405384 452169 405412 572047
rect 405464 571872 405516 571878
rect 405464 571814 405516 571820
rect 405370 452160 405426 452169
rect 405370 452095 405426 452104
rect 405476 451994 405504 571814
rect 405568 452033 405596 572319
rect 405648 571804 405700 571810
rect 405648 571746 405700 571752
rect 405660 453422 405688 571746
rect 405648 453416 405700 453422
rect 405648 453358 405700 453364
rect 405554 452024 405610 452033
rect 405464 451988 405516 451994
rect 405554 451959 405610 451968
rect 405464 451930 405516 451936
rect 405188 447908 405240 447914
rect 405188 447850 405240 447856
rect 406396 425814 406424 574398
rect 406488 445097 406516 574670
rect 406580 453490 406608 574738
rect 407672 538892 407724 538898
rect 407672 538834 407724 538840
rect 407212 491292 407264 491298
rect 407212 491234 407264 491240
rect 407120 491224 407172 491230
rect 407120 491166 407172 491172
rect 407132 490929 407160 491166
rect 407118 490920 407174 490929
rect 407118 490855 407174 490864
rect 407224 489977 407252 491234
rect 407210 489968 407266 489977
rect 407210 489903 407266 489912
rect 407120 488504 407172 488510
rect 407120 488446 407172 488452
rect 407132 487801 407160 488446
rect 407118 487792 407174 487801
rect 407118 487727 407174 487736
rect 407120 487144 407172 487150
rect 407120 487086 407172 487092
rect 407132 486849 407160 487086
rect 407118 486840 407174 486849
rect 407118 486775 407174 486784
rect 407118 485072 407174 485081
rect 407118 485007 407174 485016
rect 407132 484430 407160 485007
rect 407120 484424 407172 484430
rect 407120 484366 407172 484372
rect 407118 483984 407174 483993
rect 407118 483919 407174 483928
rect 407132 483070 407160 483919
rect 407120 483064 407172 483070
rect 407120 483006 407172 483012
rect 407118 482216 407174 482225
rect 407118 482151 407174 482160
rect 407132 481710 407160 482151
rect 407120 481704 407172 481710
rect 407120 481646 407172 481652
rect 407118 463992 407174 464001
rect 407118 463927 407174 463936
rect 407132 463758 407160 463927
rect 407120 463752 407172 463758
rect 407120 463694 407172 463700
rect 407684 463010 407712 538834
rect 407120 463004 407172 463010
rect 407120 462946 407172 462952
rect 407672 463004 407724 463010
rect 407672 462946 407724 462952
rect 407132 462369 407160 462946
rect 407118 462360 407174 462369
rect 407118 462295 407174 462304
rect 407118 462088 407174 462097
rect 407118 462023 407174 462032
rect 407132 461650 407160 462023
rect 407120 461644 407172 461650
rect 407120 461586 407172 461592
rect 406568 453484 406620 453490
rect 406568 453426 406620 453432
rect 406474 445088 406530 445097
rect 406474 445023 406530 445032
rect 406384 425808 406436 425814
rect 406384 425750 406436 425756
rect 405096 425740 405148 425746
rect 405096 425682 405148 425688
rect 407776 421870 407804 698906
rect 408224 659728 408276 659734
rect 408224 659670 408276 659676
rect 408236 575482 408264 659670
rect 408224 575476 408276 575482
rect 408224 575418 408276 575424
rect 408222 574832 408278 574841
rect 408222 574767 408278 574776
rect 407856 573368 407908 573374
rect 407856 573310 407908 573316
rect 407868 422142 407896 573310
rect 407946 571976 408002 571985
rect 407946 571911 408002 571920
rect 407856 422136 407908 422142
rect 407856 422078 407908 422084
rect 407960 422006 407988 571911
rect 408040 565140 408092 565146
rect 408040 565082 408092 565088
rect 407948 422000 408000 422006
rect 407948 421942 408000 421948
rect 408052 421938 408080 565082
rect 408132 563712 408184 563718
rect 408132 563654 408184 563660
rect 408144 422074 408172 563654
rect 408236 451897 408264 574767
rect 408222 451888 408278 451897
rect 408222 451823 408278 451832
rect 408132 422068 408184 422074
rect 408132 422010 408184 422016
rect 408040 421932 408092 421938
rect 408040 421874 408092 421880
rect 407764 421864 407816 421870
rect 407764 421806 407816 421812
rect 397644 421728 397696 421734
rect 397644 421670 397696 421676
rect 396354 421560 396410 421569
rect 396354 421495 396410 421504
rect 395066 421424 395122 421433
rect 395066 421359 395122 421368
rect 393780 421252 393832 421258
rect 393780 421194 393832 421200
rect 393792 419139 393820 421194
rect 395080 419139 395108 421359
rect 396368 419139 396396 421495
rect 397656 419139 397684 421670
rect 408328 421666 408356 700266
rect 400220 421660 400272 421666
rect 400220 421602 400272 421608
rect 408316 421660 408368 421666
rect 408316 421602 408368 421608
rect 398932 421184 398984 421190
rect 398932 421126 398984 421132
rect 398944 419139 398972 421126
rect 400232 419139 400260 421602
rect 408420 421598 408448 700402
rect 409788 700392 409840 700398
rect 409788 700334 409840 700340
rect 409696 699712 409748 699718
rect 409696 699654 409748 699660
rect 409142 575104 409198 575113
rect 409142 575039 409198 575048
rect 409156 427174 409184 575039
rect 409326 574968 409382 574977
rect 409326 574903 409382 574912
rect 409420 574932 409472 574938
rect 409236 574660 409288 574666
rect 409236 574602 409288 574608
rect 409248 436898 409276 574602
rect 409236 436892 409288 436898
rect 409236 436834 409288 436840
rect 409340 432682 409368 574903
rect 409420 574874 409472 574880
rect 409432 439822 409460 574874
rect 409512 574864 409564 574870
rect 409512 574806 409564 574812
rect 409524 453354 409552 574806
rect 409708 453354 409736 699654
rect 409512 453348 409564 453354
rect 409512 453290 409564 453296
rect 409696 453348 409748 453354
rect 409696 453290 409748 453296
rect 409420 439816 409472 439822
rect 409420 439758 409472 439764
rect 409328 432676 409380 432682
rect 409328 432618 409380 432624
rect 409144 427168 409196 427174
rect 409144 427110 409196 427116
rect 409800 421734 409828 700334
rect 413664 699718 413692 703520
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 462332 700398 462360 703520
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 478524 700330 478552 703520
rect 494808 700330 494836 703520
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 478512 700324 478564 700330
rect 478512 700266 478564 700272
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 543476 699718 543504 703520
rect 546684 700392 546736 700398
rect 546684 700334 546736 700340
rect 413652 699712 413704 699718
rect 413652 699654 413704 699660
rect 543464 699712 543516 699718
rect 543464 699654 543516 699660
rect 488908 660340 488960 660346
rect 488908 660282 488960 660288
rect 488920 659705 488948 660282
rect 499856 659728 499908 659734
rect 488906 659696 488962 659705
rect 488906 659631 488962 659640
rect 499854 659696 499856 659705
rect 499908 659696 499910 659705
rect 499854 659631 499910 659640
rect 507858 654528 507914 654537
rect 507858 654463 507914 654472
rect 506570 594688 506626 594697
rect 506570 594623 506626 594632
rect 506478 593056 506534 593065
rect 506478 592991 506534 593000
rect 492678 577824 492734 577833
rect 492678 577759 492734 577768
rect 441802 577008 441858 577017
rect 441802 576943 441858 576952
rect 462870 577008 462926 577017
rect 462870 576943 462926 576952
rect 425060 575544 425112 575550
rect 425060 575486 425112 575492
rect 415400 575476 415452 575482
rect 415400 575418 415452 575424
rect 415412 575385 415440 575418
rect 425072 575385 425100 575486
rect 415398 575376 415454 575385
rect 415398 575311 415454 575320
rect 425058 575376 425114 575385
rect 425058 575311 425114 575320
rect 426438 575240 426494 575249
rect 426438 575175 426494 575184
rect 437478 575240 437534 575249
rect 437478 575175 437534 575184
rect 426452 574938 426480 575175
rect 426440 574932 426492 574938
rect 426440 574874 426492 574880
rect 437492 574870 437520 575175
rect 437480 574864 437532 574870
rect 437480 574806 437532 574812
rect 438858 574832 438914 574841
rect 438858 574767 438860 574776
rect 438912 574767 438914 574776
rect 438860 574738 438912 574744
rect 433338 574424 433394 574433
rect 433338 574359 433394 574368
rect 433352 572393 433380 574359
rect 436098 574288 436154 574297
rect 436098 574223 436154 574232
rect 440330 574288 440386 574297
rect 440330 574223 440386 574232
rect 434718 574152 434774 574161
rect 434718 574087 434774 574096
rect 433338 572384 433394 572393
rect 433338 572319 433394 572328
rect 434732 572257 434760 574087
rect 434718 572248 434774 572257
rect 434718 572183 434774 572192
rect 436112 572121 436140 574223
rect 436190 574152 436246 574161
rect 436190 574087 436246 574096
rect 437570 574152 437626 574161
rect 437570 574087 437626 574096
rect 438950 574152 439006 574161
rect 438950 574087 439006 574096
rect 440238 574152 440294 574161
rect 440238 574087 440294 574096
rect 436098 572112 436154 572121
rect 436098 572047 436154 572056
rect 436204 571810 436232 574087
rect 436192 571804 436244 571810
rect 436192 571746 436244 571752
rect 437584 539034 437612 574087
rect 438964 562358 438992 574087
rect 438952 562352 439004 562358
rect 438952 562294 439004 562300
rect 440252 540530 440280 574087
rect 440344 571878 440372 574223
rect 441618 574152 441674 574161
rect 441618 574087 441674 574096
rect 440332 571872 440384 571878
rect 440332 571814 440384 571820
rect 440240 540524 440292 540530
rect 440240 540466 440292 540472
rect 441632 540394 441660 574087
rect 441816 571946 441844 576943
rect 455510 576192 455566 576201
rect 455510 576127 455566 576136
rect 459282 576192 459338 576201
rect 459282 576127 459338 576136
rect 448518 575104 448574 575113
rect 448518 575039 448574 575048
rect 444378 574832 444434 574841
rect 444378 574767 444434 574776
rect 444392 574734 444420 574767
rect 444380 574728 444432 574734
rect 444380 574670 444432 574676
rect 448532 574598 448560 575039
rect 451278 574696 451334 574705
rect 451278 574631 451280 574640
rect 451332 574631 451334 574640
rect 451280 574602 451332 574608
rect 448520 574592 448572 574598
rect 448520 574534 448572 574540
rect 451278 574560 451334 574569
rect 451278 574495 451280 574504
rect 451332 574495 451334 574504
rect 455418 574560 455474 574569
rect 455418 574495 455474 574504
rect 451280 574466 451332 574472
rect 455432 574462 455460 574495
rect 455420 574456 455472 574462
rect 455420 574398 455472 574404
rect 443090 574288 443146 574297
rect 443090 574223 443146 574232
rect 444562 574288 444618 574297
rect 444562 574223 444618 574232
rect 445850 574288 445906 574297
rect 445850 574223 445906 574232
rect 447230 574288 447286 574297
rect 447230 574223 447286 574232
rect 449990 574288 450046 574297
rect 449990 574223 450046 574232
rect 452750 574288 452806 574297
rect 452750 574223 452806 574232
rect 454130 574288 454186 574297
rect 454130 574223 454186 574232
rect 442998 574152 443054 574161
rect 442998 574087 443054 574096
rect 441804 571940 441856 571946
rect 441804 571882 441856 571888
rect 443012 556850 443040 574087
rect 443104 572694 443132 574223
rect 444470 574152 444526 574161
rect 444470 574087 444526 574096
rect 443092 572688 443144 572694
rect 443092 572630 443144 572636
rect 444484 566506 444512 574087
rect 444472 566500 444524 566506
rect 444472 566442 444524 566448
rect 444576 563786 444604 574223
rect 445758 574152 445814 574161
rect 445758 574087 445814 574096
rect 444564 563780 444616 563786
rect 444564 563722 444616 563728
rect 443000 556844 443052 556850
rect 443000 556786 443052 556792
rect 445772 541754 445800 574087
rect 445864 572626 445892 574223
rect 447138 574152 447194 574161
rect 447138 574087 447194 574096
rect 447152 573442 447180 574087
rect 447140 573436 447192 573442
rect 447140 573378 447192 573384
rect 445852 572620 445904 572626
rect 445852 572562 445904 572568
rect 447244 572558 447272 574223
rect 448610 574152 448666 574161
rect 448610 574087 448666 574096
rect 449898 574152 449954 574161
rect 449898 574087 449954 574096
rect 447232 572552 447284 572558
rect 447232 572494 447284 572500
rect 445760 541748 445812 541754
rect 445760 541690 445812 541696
rect 448624 541686 448652 574087
rect 448612 541680 448664 541686
rect 448612 541622 448664 541628
rect 441620 540388 441672 540394
rect 441620 540330 441672 540336
rect 449912 539170 449940 574087
rect 450004 572490 450032 574223
rect 451278 574152 451334 574161
rect 451278 574087 451334 574096
rect 452658 574152 452714 574161
rect 452658 574087 452714 574096
rect 449992 572484 450044 572490
rect 449992 572426 450044 572432
rect 449900 539164 449952 539170
rect 449900 539106 449952 539112
rect 451292 539102 451320 574087
rect 452672 572422 452700 574087
rect 452660 572416 452712 572422
rect 452660 572358 452712 572364
rect 452764 570654 452792 574223
rect 454038 574152 454094 574161
rect 454038 574087 454094 574096
rect 452752 570648 452804 570654
rect 452752 570590 452804 570596
rect 451280 539096 451332 539102
rect 451280 539038 451332 539044
rect 437572 539028 437624 539034
rect 437572 538970 437624 538976
rect 454052 538966 454080 574087
rect 454144 572354 454172 574223
rect 454132 572348 454184 572354
rect 454132 572290 454184 572296
rect 455524 569226 455552 576127
rect 458178 574424 458234 574433
rect 458178 574359 458180 574368
rect 458232 574359 458234 574368
rect 458180 574330 458232 574336
rect 456890 574288 456946 574297
rect 456890 574223 456946 574232
rect 455602 574152 455658 574161
rect 455602 574087 455658 574096
rect 456798 574152 456854 574161
rect 456798 574087 456854 574096
rect 455512 569220 455564 569226
rect 455512 569162 455564 569168
rect 455616 551342 455644 574087
rect 455604 551336 455656 551342
rect 455604 551278 455656 551284
rect 456812 539374 456840 574087
rect 456904 572286 456932 574223
rect 458362 574152 458418 574161
rect 458362 574087 458418 574096
rect 456892 572280 456944 572286
rect 456892 572222 456944 572228
rect 456800 539368 456852 539374
rect 456800 539310 456852 539316
rect 458376 539306 458404 574087
rect 459296 572218 459324 576127
rect 459558 574424 459614 574433
rect 459558 574359 459614 574368
rect 459572 574190 459600 574359
rect 462884 574326 462912 576943
rect 468482 576192 468538 576201
rect 468482 576127 468538 576136
rect 466458 575240 466514 575249
rect 466458 575175 466514 575184
rect 466472 575006 466500 575175
rect 466460 575000 466512 575006
rect 466460 574942 466512 574948
rect 463790 574560 463846 574569
rect 463790 574495 463846 574504
rect 462872 574320 462924 574326
rect 461122 574288 461178 574297
rect 462872 574262 462924 574268
rect 461122 574223 461178 574232
rect 459560 574184 459612 574190
rect 459560 574126 459612 574132
rect 459650 574152 459706 574161
rect 459650 574087 459706 574096
rect 459284 572212 459336 572218
rect 459284 572154 459336 572160
rect 458364 539300 458416 539306
rect 458364 539242 458416 539248
rect 459664 539238 459692 574087
rect 461136 567866 461164 574223
rect 461306 574152 461362 574161
rect 461306 574087 461362 574096
rect 462410 574152 462466 574161
rect 462410 574087 462466 574096
rect 463698 574152 463754 574161
rect 463698 574087 463754 574096
rect 461320 572150 461348 574087
rect 461308 572144 461360 572150
rect 461308 572086 461360 572092
rect 461124 567860 461176 567866
rect 461124 567802 461176 567808
rect 462424 560998 462452 574087
rect 462412 560992 462464 560998
rect 462412 560934 462464 560940
rect 463712 552702 463740 574087
rect 463804 572082 463832 574495
rect 465078 574424 465134 574433
rect 465078 574359 465134 574368
rect 464342 574288 464398 574297
rect 465092 574258 465120 574359
rect 464342 574223 464398 574232
rect 465080 574252 465132 574258
rect 463792 572076 463844 572082
rect 463792 572018 463844 572024
rect 464356 559570 464384 574223
rect 465080 574194 465132 574200
rect 466458 574152 466514 574161
rect 466458 574087 466514 574096
rect 466642 574152 466698 574161
rect 466642 574087 466698 574096
rect 467838 574152 467894 574161
rect 467838 574087 467894 574096
rect 466472 572014 466500 574087
rect 466460 572008 466512 572014
rect 466460 571950 466512 571956
rect 464344 559564 464396 559570
rect 464344 559506 464396 559512
rect 466656 558210 466684 574087
rect 466644 558204 466696 558210
rect 466644 558146 466696 558152
rect 467852 554062 467880 574087
rect 468496 555490 468524 576127
rect 492692 574530 492720 577759
rect 492954 576872 493010 576881
rect 492954 576807 493010 576816
rect 490564 574524 490616 574530
rect 490564 574466 490616 574472
rect 492680 574524 492732 574530
rect 492680 574466 492732 574472
rect 480904 574320 480956 574326
rect 470690 574288 470746 574297
rect 480904 574262 480956 574268
rect 470690 574223 470746 574232
rect 470598 574152 470654 574161
rect 470598 574087 470654 574096
rect 468484 555484 468536 555490
rect 468484 555426 468536 555432
rect 467840 554056 467892 554062
rect 467840 553998 467892 554004
rect 463700 552696 463752 552702
rect 463700 552638 463752 552644
rect 470612 540462 470640 574087
rect 470704 540870 470732 574223
rect 471978 574152 472034 574161
rect 471978 574087 472034 574096
rect 473358 574152 473414 574161
rect 473358 574087 473414 574096
rect 474738 574152 474794 574161
rect 474738 574087 474794 574096
rect 476118 574152 476174 574161
rect 476118 574087 476174 574096
rect 470692 540864 470744 540870
rect 470692 540806 470744 540812
rect 471992 540802 472020 574087
rect 471980 540796 472032 540802
rect 471980 540738 472032 540744
rect 473372 540734 473400 574087
rect 473360 540728 473412 540734
rect 473360 540670 473412 540676
rect 474752 540666 474780 574087
rect 474740 540660 474792 540666
rect 474740 540602 474792 540608
rect 476132 540598 476160 574087
rect 480916 545766 480944 574262
rect 487804 574252 487856 574258
rect 487804 574194 487856 574200
rect 485044 574184 485096 574190
rect 485044 574126 485096 574132
rect 485056 550594 485084 574126
rect 485044 550588 485096 550594
rect 485044 550530 485096 550536
rect 487816 549234 487844 574194
rect 487804 549228 487856 549234
rect 487804 549170 487856 549176
rect 490576 547874 490604 574466
rect 492678 574424 492734 574433
rect 492678 574359 492734 574368
rect 492692 574326 492720 574359
rect 492680 574320 492732 574326
rect 492680 574262 492732 574268
rect 492770 574288 492826 574297
rect 492770 574223 492772 574232
rect 492824 574223 492826 574232
rect 492772 574194 492824 574200
rect 492968 574190 492996 576807
rect 492956 574184 493008 574190
rect 492956 574126 493008 574132
rect 490564 547868 490616 547874
rect 490564 547810 490616 547816
rect 480904 545760 480956 545766
rect 480904 545702 480956 545708
rect 506492 543726 506520 592991
rect 506584 576065 506612 594623
rect 506570 576056 506626 576065
rect 506570 575991 506626 576000
rect 506480 543720 506532 543726
rect 506480 543662 506532 543668
rect 507872 543017 507900 654463
rect 507950 591696 508006 591705
rect 507950 591631 508006 591640
rect 507964 545086 507992 591631
rect 507952 545080 508004 545086
rect 507952 545022 508004 545028
rect 507858 543008 507914 543017
rect 507858 542943 507914 542952
rect 476120 540592 476172 540598
rect 476120 540534 476172 540540
rect 470600 540456 470652 540462
rect 470600 540398 470652 540404
rect 527180 540320 527232 540326
rect 527178 540288 527180 540297
rect 527232 540288 527234 540297
rect 527178 540223 527234 540232
rect 528836 540252 528888 540258
rect 528836 540194 528888 540200
rect 528848 539753 528876 540194
rect 528834 539744 528890 539753
rect 528834 539679 528890 539688
rect 459652 539232 459704 539238
rect 459652 539174 459704 539180
rect 454040 538960 454092 538966
rect 454040 538902 454092 538908
rect 540796 538892 540848 538898
rect 540796 538834 540848 538840
rect 540808 538801 540836 538834
rect 540794 538792 540850 538801
rect 540794 538727 540850 538736
rect 443642 453656 443698 453665
rect 443642 453591 443698 453600
rect 425426 452568 425482 452577
rect 425426 452503 425482 452512
rect 426898 452568 426954 452577
rect 426898 452503 426954 452512
rect 428462 452568 428518 452577
rect 428462 452503 428518 452512
rect 432050 452568 432106 452577
rect 432050 452503 432106 452512
rect 433706 452568 433762 452577
rect 433706 452503 433762 452512
rect 434718 452568 434774 452577
rect 434718 452503 434774 452512
rect 436282 452568 436338 452577
rect 436282 452503 436338 452512
rect 425440 451926 425468 452503
rect 425428 451920 425480 451926
rect 425428 451862 425480 451868
rect 426912 451382 426940 452503
rect 426900 451376 426952 451382
rect 426900 451318 426952 451324
rect 421840 450152 421892 450158
rect 421840 450094 421892 450100
rect 410524 450016 410576 450022
rect 410524 449958 410576 449964
rect 410536 422210 410564 449958
rect 413284 449948 413336 449954
rect 413284 449890 413336 449896
rect 410524 422204 410576 422210
rect 410524 422146 410576 422152
rect 409788 421728 409840 421734
rect 409788 421670 409840 421676
rect 407580 421592 407632 421598
rect 407580 421534 407632 421540
rect 408408 421592 408460 421598
rect 408408 421534 408460 421540
rect 403900 421524 403952 421530
rect 403900 421466 403952 421472
rect 401598 421288 401654 421297
rect 401598 421223 401654 421232
rect 401612 419139 401640 421223
rect 402980 419756 403032 419762
rect 402980 419698 403032 419704
rect 393792 419111 394166 419139
rect 395080 419111 395454 419139
rect 396368 419111 396650 419139
rect 397656 419111 397938 419139
rect 398944 419111 399226 419139
rect 400232 419111 400422 419139
rect 401612 419111 401710 419139
rect 402992 419125 403020 419698
rect 403912 419139 403940 421466
rect 405186 421152 405242 421161
rect 405186 421087 405242 421096
rect 406476 421116 406528 421122
rect 405200 419139 405228 421087
rect 406476 421058 406528 421064
rect 406488 419139 406516 421058
rect 407592 419139 407620 421534
rect 408868 421456 408920 421462
rect 408868 421398 408920 421404
rect 408880 419139 408908 421398
rect 413296 421054 413324 449890
rect 415400 421388 415452 421394
rect 415400 421330 415452 421336
rect 412824 421048 412876 421054
rect 411442 421016 411498 421025
rect 412824 420990 412876 420996
rect 413284 421048 413336 421054
rect 413284 420990 413336 420996
rect 411442 420951 411498 420960
rect 410156 419620 410208 419626
rect 410156 419562 410208 419568
rect 410168 419139 410196 419562
rect 411456 419139 411484 420951
rect 412836 419139 412864 420990
rect 414020 420980 414072 420986
rect 414020 420922 414072 420928
rect 414032 419139 414060 420922
rect 415412 419139 415440 421330
rect 416780 421320 416832 421326
rect 416780 421262 416832 421268
rect 403912 419111 404194 419139
rect 405200 419111 405482 419139
rect 406488 419111 406770 419139
rect 407592 419111 407966 419139
rect 408880 419111 409254 419139
rect 410168 419111 410542 419139
rect 411456 419111 411738 419139
rect 412836 419111 413026 419139
rect 414032 419111 414314 419139
rect 415412 419111 415510 419139
rect 416792 419125 416820 421262
rect 420276 421048 420328 421054
rect 420276 420990 420328 420996
rect 418988 419688 419040 419694
rect 418988 419630 419040 419636
rect 417700 419552 417752 419558
rect 417700 419494 417752 419500
rect 417712 419139 417740 419494
rect 419000 419139 419028 419630
rect 420288 419139 420316 420990
rect 417712 419111 418086 419139
rect 419000 419111 419282 419139
rect 420288 419111 420570 419139
rect 421852 419125 421880 450094
rect 423036 450084 423088 450090
rect 423036 450026 423088 450032
rect 423048 419125 423076 450026
rect 424324 449268 424376 449274
rect 424324 449210 424376 449216
rect 424336 419125 424364 449210
rect 426808 434104 426860 434110
rect 426808 434046 426860 434052
rect 425244 422204 425296 422210
rect 425244 422146 425296 422152
rect 425256 419139 425284 422146
rect 425256 419111 425630 419139
rect 426820 419125 426848 434046
rect 428476 429010 428504 452503
rect 429384 450628 429436 450634
rect 429384 450570 429436 450576
rect 428464 429004 428516 429010
rect 428464 428946 428516 428952
rect 427820 421796 427872 421802
rect 427820 421738 427872 421744
rect 427832 419139 427860 421738
rect 427832 419111 428114 419139
rect 429396 419125 429424 450570
rect 430580 450560 430632 450566
rect 430580 450502 430632 450508
rect 430592 419125 430620 450502
rect 431866 444952 431922 444961
rect 431866 444887 431922 444896
rect 431880 419125 431908 444887
rect 432064 438190 432092 452503
rect 433154 450800 433210 450809
rect 433720 450770 433748 452503
rect 434732 450838 434760 452503
rect 436296 450906 436324 452503
rect 438674 452296 438730 452305
rect 438674 452231 438730 452240
rect 437662 451616 437718 451625
rect 437662 451551 437718 451560
rect 437570 451344 437626 451353
rect 437570 451279 437626 451288
rect 436284 450900 436336 450906
rect 436284 450842 436336 450848
rect 434720 450832 434772 450838
rect 434720 450774 434772 450780
rect 433154 450735 433210 450744
rect 433708 450764 433760 450770
rect 432052 438184 432104 438190
rect 432052 438126 432104 438132
rect 433168 419125 433196 450735
rect 433708 450706 433760 450712
rect 436744 446548 436796 446554
rect 436744 446490 436796 446496
rect 434352 442468 434404 442474
rect 434352 442410 434404 442416
rect 434364 419125 434392 442410
rect 435364 422136 435416 422142
rect 435364 422078 435416 422084
rect 435376 419139 435404 422078
rect 436652 422068 436704 422074
rect 436652 422010 436704 422016
rect 436664 419139 436692 422010
rect 436756 421802 436784 446490
rect 437584 423570 437612 451279
rect 437676 440230 437704 451551
rect 438122 450664 438178 450673
rect 438122 450599 438178 450608
rect 437664 440224 437716 440230
rect 437664 440166 437716 440172
rect 437572 423564 437624 423570
rect 437572 423506 437624 423512
rect 436744 421796 436796 421802
rect 436744 421738 436796 421744
rect 435376 419111 435658 419139
rect 436664 419111 436946 419139
rect 438136 419125 438164 450599
rect 438688 450566 438716 452231
rect 441618 452160 441674 452169
rect 441618 452095 441674 452104
rect 442998 452160 443054 452169
rect 442998 452095 443054 452104
rect 440238 451616 440294 451625
rect 440238 451551 440294 451560
rect 438950 451344 439006 451353
rect 438950 451279 439006 451288
rect 438676 450560 438728 450566
rect 438676 450502 438728 450508
rect 438964 440162 438992 451279
rect 439412 443692 439464 443698
rect 439412 443634 439464 443640
rect 438952 440156 439004 440162
rect 438952 440098 439004 440104
rect 439424 419125 439452 443634
rect 440252 423638 440280 451551
rect 441526 451344 441582 451353
rect 441526 451279 441582 451288
rect 441540 427174 441568 451279
rect 441528 427168 441580 427174
rect 441528 427110 441580 427116
rect 441632 425649 441660 452095
rect 443012 441590 443040 452095
rect 443656 450634 443684 453591
rect 468300 453348 468352 453354
rect 468300 453290 468352 453296
rect 450266 452568 450322 452577
rect 450266 452503 450322 452512
rect 452842 452568 452898 452577
rect 452842 452503 452898 452512
rect 466182 452568 466238 452577
rect 466182 452503 466184 452512
rect 445758 452160 445814 452169
rect 445758 452095 445814 452104
rect 447046 452160 447102 452169
rect 447046 452095 447102 452104
rect 448610 452160 448666 452169
rect 448610 452095 448666 452104
rect 444470 451344 444526 451353
rect 444470 451279 444526 451288
rect 443644 450628 443696 450634
rect 443644 450570 443696 450576
rect 443000 441584 443052 441590
rect 443000 441526 443052 441532
rect 444484 439686 444512 451279
rect 445666 450528 445722 450537
rect 445666 450463 445722 450472
rect 444472 439680 444524 439686
rect 444472 439622 444524 439628
rect 444472 439544 444524 439550
rect 444472 439486 444524 439492
rect 443182 438152 443238 438161
rect 443182 438087 443238 438096
rect 441618 425640 441674 425649
rect 441618 425575 441674 425584
rect 440240 423632 440292 423638
rect 440240 423574 440292 423580
rect 440332 422000 440384 422006
rect 440332 421942 440384 421948
rect 440344 419139 440372 421942
rect 441712 421932 441764 421938
rect 441712 421874 441764 421880
rect 441724 419139 441752 421874
rect 440344 419111 440718 419139
rect 441724 419111 441914 419139
rect 443196 419125 443224 438087
rect 444484 419125 444512 439486
rect 445680 419125 445708 450463
rect 445772 426426 445800 452095
rect 445850 451344 445906 451353
rect 445850 451279 445906 451288
rect 445864 427786 445892 451279
rect 447060 439550 447088 452095
rect 447230 451344 447286 451353
rect 447230 451279 447286 451288
rect 448518 451344 448574 451353
rect 448518 451279 448574 451288
rect 447048 439544 447100 439550
rect 447048 439486 447100 439492
rect 445852 427780 445904 427786
rect 445852 427722 445904 427728
rect 447244 427718 447272 451279
rect 448532 447914 448560 451279
rect 448520 447908 448572 447914
rect 448520 447850 448572 447856
rect 448244 440904 448296 440910
rect 448244 440846 448296 440852
rect 447784 430228 447836 430234
rect 447784 430170 447836 430176
rect 447232 427712 447284 427718
rect 447232 427654 447284 427660
rect 445760 426420 445812 426426
rect 445760 426362 445812 426368
rect 447796 421870 447824 430170
rect 446588 421864 446640 421870
rect 446588 421806 446640 421812
rect 447784 421864 447836 421870
rect 447784 421806 447836 421812
rect 446600 419139 446628 421806
rect 446600 419111 446974 419139
rect 448256 419125 448284 440846
rect 448624 427106 448652 452095
rect 450280 451178 450308 452503
rect 451370 452160 451426 452169
rect 451370 452095 451426 452104
rect 451186 451344 451242 451353
rect 451186 451279 451242 451288
rect 450268 451172 450320 451178
rect 450268 451114 450320 451120
rect 449440 447160 449492 447166
rect 449440 447102 449492 447108
rect 448612 427100 448664 427106
rect 448612 427042 448664 427048
rect 449452 419125 449480 447102
rect 450728 442332 450780 442338
rect 450728 442274 450780 442280
rect 450740 419125 450768 442274
rect 451200 434110 451228 451279
rect 451188 434104 451240 434110
rect 451188 434046 451240 434052
rect 451384 429146 451412 452095
rect 452750 451344 452806 451353
rect 452750 451279 452806 451288
rect 452016 446412 452068 446418
rect 452016 446354 452068 446360
rect 451372 429140 451424 429146
rect 451372 429082 451424 429088
rect 452028 419125 452056 446354
rect 452764 429078 452792 451279
rect 452856 451246 452884 452503
rect 466236 452503 466238 452512
rect 466550 452568 466606 452577
rect 467930 452568 467986 452577
rect 466550 452503 466606 452512
rect 467104 452532 467156 452538
rect 466184 452474 466236 452480
rect 454130 452296 454186 452305
rect 454130 452231 454186 452240
rect 462318 452296 462374 452305
rect 462318 452231 462374 452240
rect 453670 452160 453726 452169
rect 453670 452095 453726 452104
rect 452844 451240 452896 451246
rect 452844 451182 452896 451188
rect 453684 446418 453712 452095
rect 454144 450702 454172 452231
rect 456706 452160 456762 452169
rect 456706 452095 456762 452104
rect 459742 452160 459798 452169
rect 459742 452095 459798 452104
rect 455510 451344 455566 451353
rect 455510 451279 455566 451288
rect 454132 450696 454184 450702
rect 454132 450638 454184 450644
rect 453672 446412 453724 446418
rect 453672 446354 453724 446360
rect 454500 441108 454552 441114
rect 454500 441050 454552 441056
rect 453210 432576 453266 432585
rect 453210 432511 453266 432520
rect 452752 429072 452804 429078
rect 452752 429014 452804 429020
rect 453224 419125 453252 432511
rect 454512 419125 454540 441050
rect 455524 428534 455552 451279
rect 456720 443698 456748 452095
rect 459466 451616 459522 451625
rect 459466 451551 459522 451560
rect 456890 451344 456946 451353
rect 456890 451279 456946 451288
rect 458270 451344 458326 451353
rect 458270 451279 458326 451288
rect 456708 443692 456760 443698
rect 456708 443634 456760 443640
rect 455788 431520 455840 431526
rect 455788 431462 455840 431468
rect 455512 428528 455564 428534
rect 455512 428470 455564 428476
rect 455800 419125 455828 431462
rect 456904 428466 456932 451279
rect 456984 443828 457036 443834
rect 456984 443770 457036 443776
rect 456892 428460 456944 428466
rect 456892 428402 456944 428408
rect 456996 419125 457024 443770
rect 458180 439748 458232 439754
rect 458180 439690 458232 439696
rect 458192 419139 458220 439690
rect 458284 428670 458312 451279
rect 459480 438190 459508 451551
rect 459560 447976 459612 447982
rect 459560 447918 459612 447924
rect 459468 438184 459520 438190
rect 459468 438126 459520 438132
rect 458272 428664 458324 428670
rect 458272 428606 458324 428612
rect 458192 419111 458290 419139
rect 459572 419125 459600 447918
rect 459756 430166 459784 452095
rect 461030 449304 461086 449313
rect 461030 449239 461086 449248
rect 460756 445120 460808 445126
rect 460756 445062 460808 445068
rect 459744 430160 459796 430166
rect 459744 430102 459796 430108
rect 460768 419125 460796 445062
rect 461044 430098 461072 449239
rect 462226 449168 462282 449177
rect 462226 449103 462282 449112
rect 462044 438388 462096 438394
rect 462044 438330 462096 438336
rect 461032 430092 461084 430098
rect 461032 430034 461084 430040
rect 462056 419125 462084 438330
rect 462240 431526 462268 449103
rect 462228 431520 462280 431526
rect 462228 431462 462280 431468
rect 462332 429962 462360 452231
rect 462410 452160 462466 452169
rect 462410 452095 462466 452104
rect 463606 452160 463662 452169
rect 463606 452095 463662 452104
rect 465078 452160 465134 452169
rect 465078 452095 465134 452104
rect 462424 430030 462452 452095
rect 463620 445126 463648 452095
rect 463790 451344 463846 451353
rect 463790 451279 463846 451288
rect 463608 445120 463660 445126
rect 463608 445062 463660 445068
rect 463332 430296 463384 430302
rect 463332 430238 463384 430244
rect 462412 430024 462464 430030
rect 462412 429966 462464 429972
rect 462320 429956 462372 429962
rect 462320 429898 462372 429904
rect 463344 419125 463372 430238
rect 463804 428602 463832 451279
rect 464528 449404 464580 449410
rect 464528 449346 464580 449352
rect 463792 428596 463844 428602
rect 463792 428538 463844 428544
rect 464540 419125 464568 449346
rect 465092 431390 465120 452095
rect 466460 446616 466512 446622
rect 466460 446558 466512 446564
rect 465080 431384 465132 431390
rect 465080 431326 465132 431332
rect 466472 422294 466500 446558
rect 466564 429894 466592 452503
rect 467930 452503 467986 452512
rect 467104 452474 467156 452480
rect 467116 432682 467144 452474
rect 467104 432676 467156 432682
rect 467104 432618 467156 432624
rect 467944 431254 467972 452503
rect 468022 452296 468078 452305
rect 468022 452231 468078 452240
rect 468036 431322 468064 452231
rect 468024 431316 468076 431322
rect 468024 431258 468076 431264
rect 467932 431248 467984 431254
rect 467932 431190 467984 431196
rect 466552 429888 466604 429894
rect 466552 429830 466604 429836
rect 466472 422266 466776 422294
rect 465540 421592 465592 421598
rect 465540 421534 465592 421540
rect 465552 419139 465580 421534
rect 466748 419139 466776 422266
rect 465552 419111 465834 419139
rect 466748 419111 467122 419139
rect 468312 419125 468340 453290
rect 468666 452568 468722 452577
rect 468666 452503 468722 452512
rect 471886 452568 471942 452577
rect 471886 452503 471942 452512
rect 473542 452568 473598 452577
rect 473542 452503 473544 452512
rect 468680 451314 468708 452503
rect 468668 451308 468720 451314
rect 468668 451250 468720 451256
rect 471244 441040 471296 441046
rect 471244 440982 471296 440988
rect 471256 421938 471284 440982
rect 471900 440910 471928 452503
rect 473596 452503 473598 452512
rect 476026 452568 476082 452577
rect 478418 452568 478474 452577
rect 476026 452503 476082 452512
rect 476764 452532 476816 452538
rect 473544 452474 473596 452480
rect 476040 451314 476068 452503
rect 478418 452503 478474 452512
rect 481086 452568 481142 452577
rect 481086 452503 481088 452512
rect 476764 452474 476816 452480
rect 474004 451308 474056 451314
rect 474004 451250 474056 451256
rect 476028 451308 476080 451314
rect 476028 451250 476080 451256
rect 471888 440904 471940 440910
rect 471888 440846 471940 440852
rect 473360 435532 473412 435538
rect 473360 435474 473412 435480
rect 471244 421932 471296 421938
rect 471244 421874 471296 421880
rect 470692 421728 470744 421734
rect 470692 421670 470744 421676
rect 469588 421592 469640 421598
rect 469588 421534 469640 421540
rect 469600 419125 469628 421534
rect 470704 419139 470732 421670
rect 471980 421660 472032 421666
rect 471980 421602 472032 421608
rect 471992 419139 472020 421602
rect 470704 419111 470894 419139
rect 471992 419111 472090 419139
rect 473372 419125 473400 435474
rect 474016 428466 474044 451250
rect 476776 439686 476804 452474
rect 478432 449274 478460 452503
rect 481140 452503 481142 452512
rect 483478 452568 483534 452577
rect 487066 452568 487122 452577
rect 483478 452503 483534 452512
rect 485136 452532 485188 452538
rect 481088 452474 481140 452480
rect 483492 452470 483520 452503
rect 487066 452503 487122 452512
rect 488446 452568 488502 452577
rect 488446 452503 488502 452512
rect 491022 452568 491078 452577
rect 491022 452503 491078 452512
rect 493598 452568 493654 452577
rect 493598 452503 493600 452512
rect 485136 452474 485188 452480
rect 483480 452464 483532 452470
rect 483480 452406 483532 452412
rect 480904 451308 480956 451314
rect 480904 451250 480956 451256
rect 478420 449268 478472 449274
rect 478420 449210 478472 449216
rect 476764 439680 476816 439686
rect 476764 439622 476816 439628
rect 478420 439612 478472 439618
rect 478420 439554 478472 439560
rect 477132 435464 477184 435470
rect 477132 435406 477184 435412
rect 474004 428460 474056 428466
rect 474004 428402 474056 428408
rect 474648 421728 474700 421734
rect 474648 421670 474700 421676
rect 474660 419125 474688 421670
rect 475844 421660 475896 421666
rect 475844 421602 475896 421608
rect 475856 419125 475884 421602
rect 477144 419125 477172 435406
rect 478432 419125 478460 439554
rect 479616 428732 479668 428738
rect 479616 428674 479668 428680
rect 479628 419125 479656 428674
rect 480916 425746 480944 451250
rect 485044 438320 485096 438326
rect 485044 438262 485096 438268
rect 480904 425740 480956 425746
rect 480904 425682 480956 425688
rect 480628 424788 480680 424794
rect 480628 424730 480680 424736
rect 480640 419139 480668 424730
rect 481916 424720 481968 424726
rect 481916 424662 481968 424668
rect 481928 419139 481956 424662
rect 483204 424652 483256 424658
rect 483204 424594 483256 424600
rect 483216 419139 483244 424594
rect 484400 421796 484452 421802
rect 484400 421738 484452 421744
rect 484412 419139 484440 421738
rect 485056 420986 485084 438262
rect 485148 436898 485176 452474
rect 487080 442338 487108 452503
rect 487804 452464 487856 452470
rect 487804 452406 487856 452412
rect 487068 442332 487120 442338
rect 487068 442274 487120 442280
rect 485136 436892 485188 436898
rect 485136 436834 485188 436840
rect 487816 423094 487844 452406
rect 488460 427106 488488 452503
rect 490932 449336 490984 449342
rect 490932 449278 490984 449284
rect 489736 436824 489788 436830
rect 489736 436766 489788 436772
rect 488448 427100 488500 427106
rect 488448 427042 488500 427048
rect 487804 423088 487856 423094
rect 487804 423030 487856 423036
rect 488172 421932 488224 421938
rect 488172 421874 488224 421880
rect 485780 421864 485832 421870
rect 485780 421806 485832 421812
rect 485044 420980 485096 420986
rect 485044 420922 485096 420928
rect 485792 419139 485820 421806
rect 487160 420980 487212 420986
rect 487160 420922 487212 420928
rect 480640 419111 480922 419139
rect 481928 419111 482210 419139
rect 483216 419111 483406 419139
rect 484412 419111 484694 419139
rect 485792 419111 485982 419139
rect 487172 419125 487200 420922
rect 488184 419139 488212 421874
rect 488184 419111 488466 419139
rect 489748 419125 489776 436766
rect 490944 419125 490972 449278
rect 491036 446554 491064 452503
rect 493652 452503 493654 452512
rect 495990 452568 496046 452577
rect 499486 452568 499542 452577
rect 495990 452503 496046 452512
rect 497464 452532 497516 452538
rect 493600 452474 493652 452480
rect 496004 451382 496032 452503
rect 499486 452503 499542 452512
rect 501234 452568 501290 452577
rect 501234 452503 501290 452512
rect 503534 452568 503590 452577
rect 505926 452568 505982 452577
rect 503534 452503 503536 452512
rect 497464 452474 497516 452480
rect 495992 451376 496044 451382
rect 495992 451318 496044 451324
rect 491024 446548 491076 446554
rect 491024 446490 491076 446496
rect 494704 446480 494756 446486
rect 494704 446422 494756 446428
rect 492220 442400 492272 442406
rect 492220 442342 492272 442348
rect 492232 419125 492260 442342
rect 493508 438252 493560 438258
rect 493508 438194 493560 438200
rect 493520 419125 493548 438194
rect 494716 419125 494744 446422
rect 497476 438258 497504 452474
rect 498476 445052 498528 445058
rect 498476 444994 498528 445000
rect 497464 438252 497516 438258
rect 497464 438194 497516 438200
rect 495716 423020 495768 423026
rect 495716 422962 495768 422968
rect 495728 419139 495756 422962
rect 497004 422952 497056 422958
rect 497004 422894 497056 422900
rect 497016 419139 497044 422894
rect 495728 419111 496010 419139
rect 497016 419111 497298 419139
rect 498488 419125 498516 444994
rect 499500 421802 499528 452503
rect 501248 447982 501276 452503
rect 503588 452503 503590 452512
rect 504364 452532 504416 452538
rect 503536 452474 503588 452480
rect 509146 452568 509202 452577
rect 505926 452503 505928 452512
rect 504364 452474 504416 452480
rect 505980 452503 505982 452512
rect 507124 452532 507176 452538
rect 505928 452474 505980 452480
rect 509146 452503 509202 452512
rect 511906 452568 511962 452577
rect 511906 452503 511962 452512
rect 514666 452568 514722 452577
rect 514666 452503 514722 452512
rect 516046 452568 516102 452577
rect 516046 452503 516102 452512
rect 507124 452474 507176 452480
rect 501236 447976 501288 447982
rect 501236 447918 501288 447924
rect 503536 447840 503588 447846
rect 503536 447782 503588 447788
rect 499764 443760 499816 443766
rect 499764 443702 499816 443708
rect 499488 421796 499540 421802
rect 499488 421738 499540 421744
rect 499776 419125 499804 443702
rect 501052 440972 501104 440978
rect 501052 440914 501104 440920
rect 501064 419125 501092 440914
rect 502248 431452 502300 431458
rect 502248 431394 502300 431400
rect 502260 419125 502288 431394
rect 503548 419125 503576 447782
rect 504376 425814 504404 452474
rect 507136 443766 507164 452474
rect 507124 443760 507176 443766
rect 507124 443702 507176 443708
rect 507308 436756 507360 436762
rect 507308 436698 507360 436704
rect 506020 435396 506072 435402
rect 506020 435338 506072 435344
rect 504824 434036 504876 434042
rect 504824 433978 504876 433984
rect 504364 425808 504416 425814
rect 504364 425750 504416 425756
rect 504836 419125 504864 433978
rect 506032 419125 506060 435338
rect 507320 419125 507348 436698
rect 508596 432608 508648 432614
rect 508596 432550 508648 432556
rect 508608 419125 508636 432550
rect 509160 421870 509188 452503
rect 509792 449200 509844 449206
rect 509792 449142 509844 449148
rect 509148 421864 509200 421870
rect 509148 421806 509200 421812
rect 509804 419125 509832 449142
rect 511920 434042 511948 452503
rect 511908 434036 511960 434042
rect 511908 433978 511960 433984
rect 510804 424584 510856 424590
rect 510804 424526 510856 424532
rect 510816 419139 510844 424526
rect 512184 424516 512236 424522
rect 512184 424458 512236 424464
rect 512196 419139 512224 424458
rect 513380 424448 513432 424454
rect 513380 424390 513432 424396
rect 513392 419139 513420 424390
rect 514680 421938 514708 452503
rect 516060 450702 516088 452503
rect 530584 451376 530636 451382
rect 530584 451318 530636 451324
rect 516048 450696 516100 450702
rect 516048 450638 516100 450644
rect 519912 450628 519964 450634
rect 519912 450570 519964 450576
rect 517336 450560 517388 450566
rect 517336 450502 517388 450508
rect 514852 442264 514904 442270
rect 514852 442206 514904 442212
rect 514668 421932 514720 421938
rect 514668 421874 514720 421880
rect 510816 419111 511098 419139
rect 512196 419111 512386 419139
rect 513392 419111 513582 419139
rect 514864 419125 514892 442206
rect 516140 424380 516192 424386
rect 516140 424322 516192 424328
rect 516152 419125 516180 424322
rect 517348 419125 517376 450502
rect 518624 427168 518676 427174
rect 518624 427110 518676 427116
rect 518636 419125 518664 427110
rect 519924 419125 519952 450570
rect 522396 447908 522448 447914
rect 522396 447850 522448 447856
rect 521108 439544 521160 439550
rect 521108 439486 521160 439492
rect 521120 419125 521148 439486
rect 522408 419125 522436 447850
rect 524880 446412 524932 446418
rect 524880 446354 524932 446360
rect 523684 434104 523736 434110
rect 523684 434046 523736 434052
rect 523696 419125 523724 434046
rect 524892 419125 524920 446354
rect 529940 445120 529992 445126
rect 529940 445062 529992 445068
rect 526168 443692 526220 443698
rect 526168 443634 526220 443640
rect 526180 419125 526208 443634
rect 527456 438184 527508 438190
rect 527456 438126 527508 438132
rect 527468 419125 527496 438126
rect 528652 431520 528704 431526
rect 528652 431462 528704 431468
rect 528664 419125 528692 431462
rect 529952 419125 529980 445062
rect 530596 422006 530624 451318
rect 537484 449268 537536 449274
rect 537484 449210 537536 449216
rect 533712 440904 533764 440910
rect 533712 440846 533764 440852
rect 531228 432676 531280 432682
rect 531228 432618 531280 432624
rect 530584 422000 530636 422006
rect 530584 421942 530636 421948
rect 531240 419125 531268 432618
rect 532424 428460 532476 428466
rect 532424 428402 532476 428408
rect 532436 419125 532464 428402
rect 533724 419125 533752 440846
rect 535000 439680 535052 439686
rect 535000 439622 535052 439628
rect 535012 419125 535040 439622
rect 536196 425740 536248 425746
rect 536196 425682 536248 425688
rect 536208 419125 536236 425682
rect 537496 419125 537524 449210
rect 543740 446548 543792 446554
rect 543740 446490 543792 446496
rect 541256 442332 541308 442338
rect 541256 442274 541308 442280
rect 538772 436892 538824 436898
rect 538772 436834 538824 436840
rect 538784 419125 538812 436834
rect 539692 423088 539744 423094
rect 539692 423030 539744 423036
rect 539704 419139 539732 423030
rect 539704 419111 539986 419139
rect 541268 419125 541296 442274
rect 542544 427100 542596 427106
rect 542544 427042 542596 427048
rect 542556 419125 542584 427042
rect 543752 419125 543780 446490
rect 545028 438252 545080 438258
rect 545028 438194 545080 438200
rect 545040 419125 545068 438194
rect 545948 422000 546000 422006
rect 545948 421942 546000 421948
rect 545960 419139 545988 421942
rect 546696 421734 546724 700334
rect 559668 700330 559696 703520
rect 546776 700324 546828 700330
rect 546776 700266 546828 700272
rect 548524 700324 548576 700330
rect 548524 700266 548576 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 546684 421728 546736 421734
rect 546684 421670 546736 421676
rect 546788 421598 546816 700266
rect 547880 699712 547932 699718
rect 547880 699654 547932 699660
rect 547236 421796 547288 421802
rect 547236 421738 547288 421744
rect 546776 421592 546828 421598
rect 546776 421534 546828 421540
rect 547248 419139 547276 421738
rect 547892 421666 547920 699654
rect 548536 435538 548564 700266
rect 580446 697232 580502 697241
rect 580446 697167 580502 697176
rect 580460 696998 580488 697167
rect 577504 696992 577556 696998
rect 577504 696934 577556 696940
rect 580448 696992 580500 696998
rect 580448 696934 580500 696940
rect 570604 670744 570656 670750
rect 570604 670686 570656 670692
rect 560944 643136 560996 643142
rect 560944 643078 560996 643084
rect 549258 533216 549314 533225
rect 549258 533151 549314 533160
rect 548800 447976 548852 447982
rect 548800 447918 548852 447924
rect 548524 435532 548576 435538
rect 548524 435474 548576 435480
rect 547880 421660 547932 421666
rect 547880 421602 547932 421608
rect 545960 419111 546334 419139
rect 547248 419111 547530 419139
rect 548812 419125 548840 447918
rect 549272 422929 549300 533151
rect 549350 473376 549406 473385
rect 549350 473311 549406 473320
rect 549364 448089 549392 473311
rect 549442 471744 549498 471753
rect 549442 471679 549498 471688
rect 549456 448225 549484 471679
rect 549534 470384 549590 470393
rect 549534 470319 549590 470328
rect 549548 448361 549576 470319
rect 549626 468888 549682 468897
rect 549626 468823 549682 468832
rect 549640 448497 549668 468823
rect 549718 467664 549774 467673
rect 549718 467599 549774 467608
rect 549732 448526 549760 467599
rect 556344 450696 556396 450702
rect 556344 450638 556396 450644
rect 549720 448520 549772 448526
rect 549626 448488 549682 448497
rect 549720 448462 549772 448468
rect 549626 448423 549682 448432
rect 549534 448352 549590 448361
rect 549534 448287 549590 448296
rect 549442 448216 549498 448225
rect 549442 448151 549498 448160
rect 549350 448080 549406 448089
rect 549350 448015 549406 448024
rect 551284 443760 551336 443766
rect 551284 443702 551336 443708
rect 550088 425808 550140 425814
rect 550088 425750 550140 425756
rect 549258 422920 549314 422929
rect 549258 422855 549314 422864
rect 550100 419125 550128 425750
rect 551296 419125 551324 443702
rect 553860 434036 553912 434042
rect 553860 433978 553912 433984
rect 552204 421864 552256 421870
rect 552204 421806 552256 421812
rect 552216 419139 552244 421806
rect 552216 419111 552590 419139
rect 553872 419125 553900 433978
rect 554780 421932 554832 421938
rect 554780 421874 554832 421880
rect 554792 419139 554820 421874
rect 554792 419111 555074 419139
rect 556356 419125 556384 450638
rect 560208 415404 560260 415410
rect 560208 415346 560260 415352
rect 560220 415177 560248 415346
rect 560206 415168 560262 415177
rect 560206 415103 560262 415112
rect 560116 408468 560168 408474
rect 560116 408410 560168 408416
rect 560128 407153 560156 408410
rect 560114 407144 560170 407153
rect 560114 407079 560170 407088
rect 560024 400172 560076 400178
rect 560024 400114 560076 400120
rect 560036 399129 560064 400114
rect 560022 399120 560078 399129
rect 560022 399055 560078 399064
rect 560208 391944 560260 391950
rect 560208 391886 560260 391892
rect 560220 391241 560248 391886
rect 560206 391232 560262 391241
rect 560206 391167 560262 391176
rect 560956 383450 560984 643078
rect 567844 616888 567896 616894
rect 567844 616830 567896 616836
rect 565084 576904 565136 576910
rect 565084 576846 565136 576852
rect 561036 456816 561088 456822
rect 561036 456758 561088 456764
rect 559196 383444 559248 383450
rect 559196 383386 559248 383392
rect 560944 383444 560996 383450
rect 560944 383386 560996 383392
rect 559208 383217 559236 383386
rect 559194 383208 559250 383217
rect 559194 383143 559250 383152
rect 560208 375352 560260 375358
rect 560208 375294 560260 375300
rect 560220 375193 560248 375294
rect 560206 375184 560262 375193
rect 560206 375119 560262 375128
rect 559196 367464 559248 367470
rect 559196 367406 559248 367412
rect 559208 367305 559236 367406
rect 559194 367296 559250 367305
rect 559194 367231 559250 367240
rect 200120 365016 200172 365022
rect 200120 364958 200172 364964
rect 559564 364404 559616 364410
rect 559564 364346 559616 364352
rect 559380 320136 559432 320142
rect 559380 320078 559432 320084
rect 559392 319433 559420 320078
rect 559378 319424 559434 319433
rect 559378 319359 559434 319368
rect 559288 303476 559340 303482
rect 559288 303418 559340 303424
rect 559300 303385 559328 303418
rect 559286 303376 559342 303385
rect 559286 303311 559342 303320
rect 559012 296676 559064 296682
rect 559012 296618 559064 296624
rect 559024 295361 559052 296618
rect 559010 295352 559066 295361
rect 559010 295287 559066 295296
rect 559576 271425 559604 364346
rect 560208 360188 560260 360194
rect 560208 360130 560260 360136
rect 560220 359281 560248 360130
rect 560206 359272 560262 359281
rect 560206 359207 560262 359216
rect 559656 351892 559708 351898
rect 559656 351834 559708 351840
rect 559668 351257 559696 351834
rect 559654 351248 559710 351257
rect 559654 351183 559710 351192
rect 560208 343596 560260 343602
rect 560208 343538 560260 343544
rect 560220 343369 560248 343538
rect 560206 343360 560262 343369
rect 560206 343295 560262 343304
rect 560206 335336 560262 335345
rect 560206 335271 560208 335280
rect 560260 335271 560262 335280
rect 560208 335242 560260 335248
rect 559932 328432 559984 328438
rect 559932 328374 559984 328380
rect 559944 327321 559972 328374
rect 559930 327312 559986 327321
rect 559930 327247 559986 327256
rect 560208 311840 560260 311846
rect 560208 311782 560260 311788
rect 560220 311409 560248 311782
rect 560206 311400 560262 311409
rect 560206 311335 560262 311344
rect 561048 303482 561076 456758
rect 565096 367470 565124 576846
rect 566464 563100 566516 563106
rect 566464 563042 566516 563048
rect 565176 510672 565228 510678
rect 565176 510614 565228 510620
rect 565084 367464 565136 367470
rect 565084 367406 565136 367412
rect 565188 328438 565216 510614
rect 566476 351898 566504 563042
rect 566556 470620 566608 470626
rect 566556 470562 566608 470568
rect 566464 351892 566516 351898
rect 566464 351834 566516 351840
rect 565176 328432 565228 328438
rect 565176 328374 565228 328380
rect 565084 324352 565136 324358
rect 565084 324294 565136 324300
rect 561036 303476 561088 303482
rect 561036 303418 561088 303424
rect 560944 298172 560996 298178
rect 560944 298114 560996 298120
rect 560208 288380 560260 288386
rect 560208 288322 560260 288328
rect 560220 287473 560248 288322
rect 560206 287464 560262 287473
rect 560206 287399 560262 287408
rect 559932 280152 559984 280158
rect 559932 280094 559984 280100
rect 559944 279449 559972 280094
rect 559930 279440 559986 279449
rect 559930 279375 559986 279384
rect 559562 271416 559618 271425
rect 559562 271351 559618 271360
rect 560208 263560 560260 263566
rect 560206 263528 560208 263537
rect 560260 263528 560262 263537
rect 560206 263463 560262 263472
rect 199474 258768 199530 258777
rect 199474 258703 199530 258712
rect 560024 256692 560076 256698
rect 560024 256634 560076 256640
rect 560036 255513 560064 256634
rect 560022 255504 560078 255513
rect 560022 255439 560078 255448
rect 560208 248396 560260 248402
rect 560208 248338 560260 248344
rect 560220 247489 560248 248338
rect 560206 247480 560262 247489
rect 560206 247415 560262 247424
rect 560208 239624 560260 239630
rect 560206 239592 560208 239601
rect 560260 239592 560262 239601
rect 560206 239527 560262 239536
rect 199290 237688 199346 237697
rect 199290 237623 199346 237632
rect 560956 231742 560984 298114
rect 565096 239630 565124 324294
rect 566568 320142 566596 470562
rect 567856 375358 567884 616830
rect 567936 430636 567988 430642
rect 567936 430578 567988 430584
rect 567844 375352 567896 375358
rect 567844 375294 567896 375300
rect 566556 320136 566608 320142
rect 566556 320078 566608 320084
rect 567948 288386 567976 430578
rect 570616 400178 570644 670686
rect 574744 590708 574796 590714
rect 574744 590650 574796 590656
rect 570696 524476 570748 524482
rect 570696 524418 570748 524424
rect 570604 400172 570656 400178
rect 570604 400114 570656 400120
rect 570604 378208 570656 378214
rect 570604 378150 570656 378156
rect 567936 288380 567988 288386
rect 567936 288322 567988 288328
rect 566464 271924 566516 271930
rect 566464 271866 566516 271872
rect 565084 239624 565136 239630
rect 565084 239566 565136 239572
rect 565084 231872 565136 231878
rect 565084 231814 565136 231820
rect 559196 231736 559248 231742
rect 559196 231678 559248 231684
rect 560944 231736 560996 231742
rect 560944 231678 560996 231684
rect 559208 231577 559236 231678
rect 559194 231568 559250 231577
rect 559194 231503 559250 231512
rect 199198 230208 199254 230217
rect 199198 230143 199254 230152
rect 199108 228472 199160 228478
rect 199108 228414 199160 228420
rect 199120 227769 199148 228414
rect 199106 227760 199162 227769
rect 199106 227695 199162 227704
rect 199016 223576 199068 223582
rect 199016 223518 199068 223524
rect 199568 223576 199620 223582
rect 560208 223576 560260 223582
rect 199568 223518 199620 223524
rect 560206 223544 560208 223553
rect 560260 223544 560262 223553
rect 199580 222941 199608 223518
rect 560206 223479 560262 223488
rect 199566 222932 199622 222941
rect 199566 222867 199622 222876
rect 198922 221504 198978 221513
rect 198922 221439 198978 221448
rect 198936 220862 198964 221439
rect 198924 220856 198976 220862
rect 198924 220798 198976 220804
rect 198738 220280 198794 220289
rect 198738 220215 198794 220224
rect 197910 219056 197966 219065
rect 197910 218991 197966 219000
rect 197924 218822 197952 218991
rect 197912 218816 197964 218822
rect 197912 218758 197964 218764
rect 197924 211614 197952 218758
rect 559564 218068 559616 218074
rect 559564 218010 559616 218016
rect 198004 215960 198056 215966
rect 198004 215902 198056 215908
rect 197912 211608 197964 211614
rect 197912 211550 197964 211556
rect 197832 210334 197952 210362
rect 197728 210248 197780 210254
rect 197728 210190 197780 210196
rect 197728 210112 197780 210118
rect 197728 210054 197780 210060
rect 197740 209234 197768 210054
rect 197924 209930 197952 210334
rect 198016 210118 198044 215902
rect 559196 215824 559248 215830
rect 559196 215766 559248 215772
rect 559208 215665 559236 215766
rect 559194 215656 559250 215665
rect 559194 215591 559250 215600
rect 198096 215416 198148 215422
rect 198094 215384 198096 215393
rect 198148 215384 198150 215393
rect 198094 215319 198150 215328
rect 198004 210112 198056 210118
rect 198004 210054 198056 210060
rect 197832 209902 197952 209930
rect 197728 209228 197780 209234
rect 197728 209170 197780 209176
rect 197726 209128 197782 209137
rect 197726 209063 197782 209072
rect 197740 206310 197768 209063
rect 197728 206304 197780 206310
rect 197728 206246 197780 206252
rect 197728 204264 197780 204270
rect 197728 204206 197780 204212
rect 197740 203017 197768 204206
rect 197726 203008 197782 203017
rect 197726 202943 197782 202952
rect 197728 192500 197780 192506
rect 197728 192442 197780 192448
rect 197740 192409 197768 192442
rect 197726 192400 197782 192409
rect 197726 192335 197782 192344
rect 197636 175976 197688 175982
rect 197636 175918 197688 175924
rect 197544 170400 197596 170406
rect 197544 170342 197596 170348
rect 197544 168360 197596 168366
rect 197544 168302 197596 168308
rect 197556 167657 197584 168302
rect 197542 167648 197598 167657
rect 197542 167583 197598 167592
rect 197544 155916 197596 155922
rect 197544 155858 197596 155864
rect 197556 154737 197584 155858
rect 197542 154728 197598 154737
rect 197542 154663 197598 154672
rect 197542 148472 197598 148481
rect 197542 148407 197598 148416
rect 197556 147694 197584 148407
rect 197544 147688 197596 147694
rect 197544 147630 197596 147636
rect 197832 141506 197860 209902
rect 197912 209228 197964 209234
rect 197912 209170 197964 209176
rect 197924 202842 197952 209170
rect 197912 202836 197964 202842
rect 197912 202778 197964 202784
rect 559576 199617 559604 218010
rect 560208 208344 560260 208350
rect 560208 208286 560260 208292
rect 560220 207641 560248 208286
rect 560206 207632 560262 207641
rect 560206 207567 560262 207576
rect 559562 199608 559618 199617
rect 559562 199543 559618 199552
rect 560944 191888 560996 191894
rect 560944 191830 560996 191836
rect 560208 191752 560260 191758
rect 560206 191720 560208 191729
rect 560260 191720 560262 191729
rect 560206 191655 560262 191664
rect 560024 184884 560076 184890
rect 560024 184826 560076 184832
rect 560036 183705 560064 184826
rect 560022 183696 560078 183705
rect 560022 183631 560078 183640
rect 197912 178288 197964 178294
rect 197910 178256 197912 178265
rect 197964 178256 197966 178265
rect 197910 178191 197966 178200
rect 560208 176656 560260 176662
rect 560208 176598 560260 176604
rect 560220 175681 560248 176598
rect 560206 175672 560262 175681
rect 560206 175607 560262 175616
rect 560956 168298 560984 191830
rect 565096 191758 565124 231814
rect 566476 215830 566504 271866
rect 570616 263566 570644 378150
rect 570708 343602 570736 524418
rect 574756 360194 574784 590650
rect 577516 408474 577544 696934
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 578882 630864 578938 630873
rect 578882 630799 578938 630808
rect 577596 484424 577648 484430
rect 577596 484366 577648 484372
rect 577504 408468 577556 408474
rect 577504 408410 577556 408416
rect 574836 404388 574888 404394
rect 574836 404330 574888 404336
rect 574744 360188 574796 360194
rect 574744 360130 574796 360136
rect 570696 343596 570748 343602
rect 570696 343538 570748 343544
rect 574848 280158 574876 404330
rect 577504 311908 577556 311914
rect 577504 311850 577556 311856
rect 574836 280152 574888 280158
rect 574836 280094 574888 280100
rect 570604 263560 570656 263566
rect 570604 263502 570656 263508
rect 567844 258120 567896 258126
rect 567844 258062 567896 258068
rect 567856 223582 567884 258062
rect 577516 248402 577544 311850
rect 577608 311846 577636 484366
rect 578896 391950 578924 630799
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 578974 537840 579030 537849
rect 578974 537775 579030 537784
rect 578884 391944 578936 391950
rect 578884 391886 578936 391892
rect 578882 351928 578938 351937
rect 578882 351863 578938 351872
rect 577596 311840 577648 311846
rect 577596 311782 577648 311788
rect 578896 256698 578924 351863
rect 578988 335306 579016 537775
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 579908 430642 579936 431559
rect 579896 430636 579948 430642
rect 579896 430578 579948 430584
rect 580276 415410 580304 683839
rect 580630 484664 580686 484673
rect 580630 484599 580686 484608
rect 580644 484430 580672 484599
rect 580632 484424 580684 484430
rect 580632 484366 580684 484372
rect 580354 418296 580410 418305
rect 580354 418231 580410 418240
rect 580264 415404 580316 415410
rect 580264 415346 580316 415352
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 578976 335300 579028 335306
rect 578976 335242 579028 335248
rect 580078 325272 580134 325281
rect 580078 325207 580134 325216
rect 580092 324358 580120 325207
rect 580080 324352 580132 324358
rect 580080 324294 580132 324300
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580368 296682 580396 418231
rect 580446 312080 580502 312089
rect 580446 312015 580502 312024
rect 580460 311914 580488 312015
rect 580448 311908 580500 311914
rect 580448 311850 580500 311856
rect 580356 296676 580408 296682
rect 580356 296618 580408 296624
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 578884 256692 578936 256698
rect 578884 256634 578936 256640
rect 577504 248396 577556 248402
rect 577504 248338 577556 248344
rect 580262 245576 580318 245585
rect 580262 245511 580318 245520
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579816 231878 579844 232319
rect 579804 231872 579856 231878
rect 579804 231814 579856 231820
rect 567844 223576 567896 223582
rect 567844 223518 567896 223524
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 579908 218074 579936 218991
rect 579896 218068 579948 218074
rect 579896 218010 579948 218016
rect 566464 215824 566516 215830
rect 566464 215766 566516 215772
rect 580276 208350 580304 245511
rect 580264 208344 580316 208350
rect 580264 208286 580316 208292
rect 580262 205728 580318 205737
rect 580262 205663 580318 205672
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 565084 191752 565136 191758
rect 565084 191694 565136 191700
rect 580276 184890 580304 205663
rect 580264 184884 580316 184890
rect 580264 184826 580316 184832
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 176662 580212 179143
rect 580172 176656 580224 176662
rect 580172 176598 580224 176604
rect 559012 168292 559064 168298
rect 559012 168234 559064 168240
rect 560944 168292 560996 168298
rect 560944 168234 560996 168240
rect 559024 167657 559052 168234
rect 559010 167648 559066 167657
rect 559010 167583 559066 167592
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 559564 165640 559616 165646
rect 559564 165582 559616 165588
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 559576 159769 559604 165582
rect 559562 159760 559618 159769
rect 559562 159695 559618 159704
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 559562 151736 559618 151745
rect 559562 151671 559618 151680
rect 197820 141500 197872 141506
rect 197820 141442 197872 141448
rect 197452 141432 197504 141438
rect 197452 141374 197504 141380
rect 197266 140992 197322 141001
rect 197266 140927 197322 140936
rect 197280 139942 197308 140927
rect 197360 140004 197412 140010
rect 197360 139946 197412 139952
rect 197268 139936 197320 139942
rect 197268 139878 197320 139884
rect 197372 139777 197400 139946
rect 197358 139768 197414 139777
rect 197358 139703 197414 139712
rect 559576 139398 559604 151671
rect 580276 144906 580304 152623
rect 560024 144900 560076 144906
rect 560024 144842 560076 144848
rect 580264 144900 580316 144906
rect 580264 144842 580316 144848
rect 560036 143721 560064 144842
rect 560022 143712 560078 143721
rect 560022 143647 560078 143656
rect 559564 139392 559616 139398
rect 580172 139392 580224 139398
rect 559564 139334 559616 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 197450 138544 197506 138553
rect 197450 138479 197506 138488
rect 197360 137896 197412 137902
rect 197360 137838 197412 137844
rect 197372 137329 197400 137838
rect 197464 137834 197492 138479
rect 197452 137828 197504 137834
rect 197452 137770 197504 137776
rect 197358 137320 197414 137329
rect 197358 137255 197414 137264
rect 197360 136604 197412 136610
rect 197360 136546 197412 136552
rect 197372 136377 197400 136546
rect 197358 136368 197414 136377
rect 197358 136303 197414 136312
rect 559286 135824 559342 135833
rect 559286 135759 559342 135768
rect 559300 135386 559328 135759
rect 559288 135380 559340 135386
rect 559288 135322 559340 135328
rect 560944 135380 560996 135386
rect 560944 135322 560996 135328
rect 197360 135244 197412 135250
rect 197360 135186 197412 135192
rect 197372 134881 197400 135186
rect 197358 134872 197414 134881
rect 197358 134807 197414 134816
rect 197360 133884 197412 133890
rect 197360 133826 197412 133832
rect 197372 133657 197400 133826
rect 197358 133648 197414 133657
rect 197358 133583 197414 133592
rect 197360 132456 197412 132462
rect 197358 132424 197360 132433
rect 197412 132424 197414 132433
rect 197358 132359 197414 132368
rect 197452 132388 197504 132394
rect 197452 132330 197504 132336
rect 197464 131209 197492 132330
rect 197450 131200 197506 131209
rect 197450 131135 197506 131144
rect 197360 131096 197412 131102
rect 197360 131038 197412 131044
rect 197372 129849 197400 131038
rect 197358 129840 197414 129849
rect 197358 129775 197414 129784
rect 197360 129736 197412 129742
rect 197360 129678 197412 129684
rect 197372 129305 197400 129678
rect 197358 129296 197414 129305
rect 197358 129231 197414 129240
rect 197360 128308 197412 128314
rect 197360 128250 197412 128256
rect 197372 128081 197400 128250
rect 197358 128072 197414 128081
rect 197358 128007 197414 128016
rect 559562 127800 559618 127809
rect 559562 127735 559618 127744
rect 197360 126948 197412 126954
rect 197360 126890 197412 126896
rect 197372 126177 197400 126890
rect 197358 126168 197414 126177
rect 197358 126103 197414 126112
rect 197360 125588 197412 125594
rect 197360 125530 197412 125536
rect 197372 124953 197400 125530
rect 197358 124944 197414 124953
rect 197358 124879 197414 124888
rect 197360 124160 197412 124166
rect 197360 124102 197412 124108
rect 197372 123729 197400 124102
rect 197358 123720 197414 123729
rect 197358 123655 197414 123664
rect 197360 122800 197412 122806
rect 197360 122742 197412 122748
rect 197372 122505 197400 122742
rect 197358 122496 197414 122505
rect 197358 122431 197414 122440
rect 197360 121440 197412 121446
rect 197360 121382 197412 121388
rect 197372 121281 197400 121382
rect 197358 121272 197414 121281
rect 197358 121207 197414 121216
rect 197360 120080 197412 120086
rect 197358 120048 197360 120057
rect 197412 120048 197414 120057
rect 197358 119983 197414 119992
rect 197452 120012 197504 120018
rect 197452 119954 197504 119960
rect 197464 118833 197492 119954
rect 558918 119776 558974 119785
rect 558918 119711 558974 119720
rect 197450 118824 197506 118833
rect 197450 118759 197506 118768
rect 558932 118726 558960 119711
rect 558920 118720 558972 118726
rect 558920 118662 558972 118668
rect 197360 118652 197412 118658
rect 197360 118594 197412 118600
rect 197372 117473 197400 118594
rect 197358 117464 197414 117473
rect 197358 117399 197414 117408
rect 197360 117224 197412 117230
rect 197360 117166 197412 117172
rect 197372 116249 197400 117166
rect 197358 116240 197414 116249
rect 197358 116175 197414 116184
rect 197360 115932 197412 115938
rect 197360 115874 197412 115880
rect 197372 115025 197400 115874
rect 197358 115016 197414 115025
rect 197358 114951 197414 114960
rect 197360 114504 197412 114510
rect 197360 114446 197412 114452
rect 197372 113801 197400 114446
rect 197358 113792 197414 113801
rect 197358 113727 197414 113736
rect 197360 113144 197412 113150
rect 197358 113112 197360 113121
rect 197412 113112 197414 113121
rect 197358 113047 197414 113056
rect 559194 111888 559250 111897
rect 559194 111823 559196 111832
rect 559248 111823 559250 111832
rect 559196 111794 559248 111800
rect 197360 111784 197412 111790
rect 197358 111752 197360 111761
rect 197412 111752 197414 111761
rect 197358 111687 197414 111696
rect 197360 110424 197412 110430
rect 197360 110366 197412 110372
rect 197372 110129 197400 110366
rect 197358 110120 197414 110129
rect 197358 110055 197414 110064
rect 197544 108996 197596 109002
rect 197544 108938 197596 108944
rect 197360 108928 197412 108934
rect 197358 108896 197360 108905
rect 197412 108896 197414 108905
rect 197358 108831 197414 108840
rect 197556 107681 197584 108938
rect 197542 107672 197598 107681
rect 197452 107636 197504 107642
rect 197542 107607 197598 107616
rect 197452 107578 197504 107584
rect 197464 106321 197492 107578
rect 197450 106312 197506 106321
rect 197360 106276 197412 106282
rect 197450 106247 197506 106256
rect 197360 106218 197412 106224
rect 197372 105097 197400 106218
rect 197358 105088 197414 105097
rect 197358 105023 197414 105032
rect 197360 104848 197412 104854
rect 197360 104790 197412 104796
rect 197372 103873 197400 104790
rect 197358 103864 197414 103873
rect 197358 103799 197414 103808
rect 197360 103488 197412 103494
rect 197360 103430 197412 103436
rect 197372 102649 197400 103430
rect 197358 102640 197414 102649
rect 197358 102575 197414 102584
rect 197360 102128 197412 102134
rect 197360 102070 197412 102076
rect 197372 101425 197400 102070
rect 197358 101416 197414 101425
rect 197358 101351 197414 101360
rect 559576 100706 559604 127735
rect 560956 126954 560984 135322
rect 560944 126948 560996 126954
rect 560944 126890 560996 126896
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 561036 118720 561088 118726
rect 561036 118662 561088 118668
rect 561048 113150 561076 118662
rect 561036 113144 561088 113150
rect 561036 113086 561088 113092
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 560944 111852 560996 111858
rect 560944 111794 560996 111800
rect 560206 103864 560262 103873
rect 560206 103799 560208 103808
rect 560260 103799 560262 103808
rect 560208 103770 560260 103776
rect 197360 100700 197412 100706
rect 197360 100642 197412 100648
rect 559564 100700 559616 100706
rect 559564 100642 559616 100648
rect 197372 100201 197400 100642
rect 197358 100192 197414 100201
rect 197358 100127 197414 100136
rect 197358 98968 197414 98977
rect 197358 98903 197414 98912
rect 197372 98054 197400 98903
rect 197360 98048 197412 98054
rect 197360 97990 197412 97996
rect 198002 97744 198058 97753
rect 198002 97679 198058 97688
rect 197358 94616 197414 94625
rect 197358 94551 197414 94560
rect 197372 93906 197400 94551
rect 197360 93900 197412 93906
rect 197360 93842 197412 93848
rect 197358 92712 197414 92721
rect 197358 92647 197414 92656
rect 197372 92546 197400 92647
rect 197360 92540 197412 92546
rect 197360 92482 197412 92488
rect 197358 91488 197414 91497
rect 197358 91423 197414 91432
rect 197372 91118 197400 91423
rect 197360 91112 197412 91118
rect 197360 91054 197412 91060
rect 197358 90264 197414 90273
rect 197358 90199 197414 90208
rect 197372 89758 197400 90199
rect 197360 89752 197412 89758
rect 197360 89694 197412 89700
rect 197358 89040 197414 89049
rect 197358 88975 197414 88984
rect 197372 88398 197400 88975
rect 197360 88392 197412 88398
rect 197360 88334 197412 88340
rect 197358 87272 197414 87281
rect 197358 87207 197414 87216
rect 197372 87038 197400 87207
rect 197360 87032 197412 87038
rect 197360 86974 197412 86980
rect 197358 86592 197414 86601
rect 197358 86527 197414 86536
rect 197372 85610 197400 86527
rect 197360 85604 197412 85610
rect 197360 85546 197412 85552
rect 197358 85368 197414 85377
rect 197358 85303 197414 85312
rect 197372 84250 197400 85303
rect 197360 84244 197412 84250
rect 197360 84186 197412 84192
rect 197358 84144 197414 84153
rect 197358 84079 197414 84088
rect 197372 82890 197400 84079
rect 197360 82884 197412 82890
rect 197360 82826 197412 82832
rect 197450 82784 197506 82793
rect 197450 82719 197506 82728
rect 197358 81560 197414 81569
rect 197464 81530 197492 82719
rect 197358 81495 197414 81504
rect 197452 81524 197504 81530
rect 197372 81462 197400 81495
rect 197452 81466 197504 81472
rect 197360 81456 197412 81462
rect 197360 81398 197412 81404
rect 197358 80200 197414 80209
rect 197358 80135 197414 80144
rect 197372 80102 197400 80135
rect 197360 80096 197412 80102
rect 197360 80038 197412 80044
rect 197358 78840 197414 78849
rect 197358 78775 197414 78784
rect 197372 78742 197400 78775
rect 197360 78736 197412 78742
rect 197360 78678 197412 78684
rect 197358 77888 197414 77897
rect 197358 77823 197414 77832
rect 197372 77314 197400 77823
rect 197360 77308 197412 77314
rect 197360 77250 197412 77256
rect 197358 76664 197414 76673
rect 197358 76599 197414 76608
rect 197372 75954 197400 76599
rect 197360 75948 197412 75954
rect 197360 75890 197412 75896
rect 197358 75440 197414 75449
rect 197358 75375 197414 75384
rect 197372 74594 197400 75375
rect 197360 74588 197412 74594
rect 197360 74530 197412 74536
rect 197358 74216 197414 74225
rect 197358 74151 197414 74160
rect 197372 73234 197400 74151
rect 197360 73228 197412 73234
rect 197360 73170 197412 73176
rect 197358 72992 197414 73001
rect 197358 72927 197414 72936
rect 197372 71806 197400 72927
rect 197360 71800 197412 71806
rect 197360 71742 197412 71748
rect 197360 70440 197412 70446
rect 197358 70408 197360 70417
rect 197412 70408 197414 70417
rect 197358 70343 197414 70352
rect 197358 63880 197414 63889
rect 197358 63815 197414 63824
rect 197372 63578 197400 63815
rect 197360 63572 197412 63578
rect 197360 63514 197412 63520
rect 197910 63064 197966 63073
rect 197910 62999 197966 63008
rect 197358 61840 197414 61849
rect 197358 61775 197414 61784
rect 197372 60790 197400 61775
rect 197360 60784 197412 60790
rect 197360 60726 197412 60732
rect 197542 60616 197598 60625
rect 197542 60551 197598 60560
rect 197556 59430 197584 60551
rect 197544 59424 197596 59430
rect 197544 59366 197596 59372
rect 197924 28898 197952 62999
rect 198016 29442 198044 97679
rect 198094 95976 198150 95985
rect 198094 95911 198150 95920
rect 198108 29850 198136 95911
rect 559746 95840 559802 95849
rect 559746 95775 559802 95784
rect 559760 95266 559788 95775
rect 559748 95260 559800 95266
rect 559748 95202 559800 95208
rect 198186 93936 198242 93945
rect 198186 93871 198242 93880
rect 198200 29918 198228 93871
rect 560206 87952 560262 87961
rect 560206 87887 560262 87896
rect 560220 87038 560248 87887
rect 560208 87032 560260 87038
rect 560208 86974 560260 86980
rect 560956 86970 560984 111794
rect 566464 103828 566516 103834
rect 566464 103770 566516 103776
rect 565084 95260 565136 95266
rect 565084 95202 565136 95208
rect 560944 86964 560996 86970
rect 560944 86906 560996 86912
rect 560022 79928 560078 79937
rect 560022 79863 560078 79872
rect 560036 78742 560064 79863
rect 560024 78736 560076 78742
rect 560024 78678 560076 78684
rect 565096 73166 565124 95202
rect 565084 73160 565136 73166
rect 565084 73102 565136 73108
rect 559194 71904 559250 71913
rect 559194 71839 559196 71848
rect 559248 71839 559250 71848
rect 560944 71868 560996 71874
rect 559196 71810 559248 71816
rect 560944 71810 560996 71816
rect 198278 71088 198334 71097
rect 198278 71023 198334 71032
rect 198188 29912 198240 29918
rect 198188 29854 198240 29860
rect 198096 29844 198148 29850
rect 198096 29786 198148 29792
rect 198292 29646 198320 71023
rect 198370 69184 198426 69193
rect 198370 69119 198426 69128
rect 198384 29714 198412 69119
rect 198462 67960 198518 67969
rect 198462 67895 198518 67904
rect 198372 29708 198424 29714
rect 198372 29650 198424 29656
rect 198280 29640 198332 29646
rect 198280 29582 198332 29588
rect 198476 29510 198504 67895
rect 198554 66736 198610 66745
rect 198554 66671 198610 66680
rect 198568 29782 198596 66671
rect 198646 65512 198702 65521
rect 198646 65447 198702 65456
rect 198556 29776 198608 29782
rect 198556 29718 198608 29724
rect 198660 29578 198688 65447
rect 560206 64016 560262 64025
rect 560206 63951 560262 63960
rect 560220 63578 560248 63951
rect 560208 63572 560260 63578
rect 560208 63514 560260 63520
rect 200132 60030 200330 60058
rect 200408 60030 200974 60058
rect 201604 60030 201710 60058
rect 202064 60030 202446 60058
rect 198740 40792 198792 40798
rect 198740 40734 198792 40740
rect 198648 29572 198700 29578
rect 198648 29514 198700 29520
rect 198464 29504 198516 29510
rect 198464 29446 198516 29452
rect 198004 29436 198056 29442
rect 198004 29378 198056 29384
rect 197912 28892 197964 28898
rect 197912 28834 197964 28840
rect 196806 26344 196862 26353
rect 196806 26279 196862 26288
rect 197912 5364 197964 5370
rect 197912 5306 197964 5312
rect 196624 3596 196676 3602
rect 196624 3538 196676 3544
rect 196544 3454 196848 3482
rect 196820 480 196848 3454
rect 197924 480 197952 5306
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 40734
rect 200132 11762 200160 60030
rect 200408 55214 200436 60030
rect 201500 58064 201552 58070
rect 201500 58006 201552 58012
rect 200224 55186 200436 55214
rect 200120 11756 200172 11762
rect 200120 11698 200172 11704
rect 200224 4826 200252 55186
rect 200304 53100 200356 53106
rect 200304 53042 200356 53048
rect 200212 4820 200264 4826
rect 200212 4762 200264 4768
rect 200316 480 200344 53042
rect 201512 7614 201540 58006
rect 201604 22778 201632 60030
rect 202064 58070 202092 60030
rect 202052 58064 202104 58070
rect 202052 58006 202104 58012
rect 203168 57730 203196 60044
rect 203444 60030 203918 60058
rect 204272 60030 204654 60058
rect 204916 60030 205390 60058
rect 205836 60030 206034 60058
rect 203156 57724 203208 57730
rect 203156 57666 203208 57672
rect 203444 45554 203472 60030
rect 202984 45526 203472 45554
rect 201684 35284 201736 35290
rect 201684 35226 201736 35232
rect 201592 22772 201644 22778
rect 201592 22714 201644 22720
rect 201696 16574 201724 35226
rect 201696 16546 202736 16574
rect 201500 7608 201552 7614
rect 201500 7550 201552 7556
rect 201500 4820 201552 4826
rect 201500 4762 201552 4768
rect 201512 480 201540 4762
rect 202708 480 202736 16546
rect 202984 11830 203012 45526
rect 204272 15910 204300 60030
rect 204916 45554 204944 60030
rect 204364 45526 204944 45554
rect 204364 24138 204392 45526
rect 205732 39432 205784 39438
rect 205732 39374 205784 39380
rect 204904 29640 204956 29646
rect 204904 29582 204956 29588
rect 204444 26988 204496 26994
rect 204444 26930 204496 26936
rect 204352 24132 204404 24138
rect 204352 24074 204404 24080
rect 204456 16574 204484 26930
rect 204456 16546 204852 16574
rect 204260 15904 204312 15910
rect 204260 15846 204312 15852
rect 202972 11824 203024 11830
rect 202972 11766 203024 11772
rect 203892 3596 203944 3602
rect 203892 3538 203944 3544
rect 203904 480 203932 3538
rect 204824 3482 204852 16546
rect 204916 3602 204944 29582
rect 205744 6914 205772 39374
rect 205836 11898 205864 60030
rect 206756 57934 206784 60044
rect 207032 60030 207506 60058
rect 207768 60030 208242 60058
rect 208412 60030 208978 60058
rect 209332 60030 209714 60058
rect 209884 60030 210450 60058
rect 206744 57928 206796 57934
rect 206744 57870 206796 57876
rect 205824 11892 205876 11898
rect 205824 11834 205876 11840
rect 205744 6886 206232 6914
rect 204904 3596 204956 3602
rect 204904 3538 204956 3544
rect 204824 3454 205128 3482
rect 205100 480 205128 3454
rect 206204 480 206232 6886
rect 207032 4894 207060 60030
rect 207768 45554 207796 60030
rect 207124 45526 207796 45554
rect 207124 8974 207152 45526
rect 207204 33788 207256 33794
rect 207204 33730 207256 33736
rect 207112 8968 207164 8974
rect 207112 8910 207164 8916
rect 207020 4888 207072 4894
rect 207020 4830 207072 4836
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207216 354 207244 33730
rect 208412 7682 208440 60030
rect 209332 45554 209360 60030
rect 209780 51808 209832 51814
rect 209780 51750 209832 51756
rect 208504 45526 209360 45554
rect 208504 11966 208532 45526
rect 208584 31204 208636 31210
rect 208584 31146 208636 31152
rect 208492 11960 208544 11966
rect 208492 11902 208544 11908
rect 208400 7676 208452 7682
rect 208400 7618 208452 7624
rect 208596 480 208624 31146
rect 209792 9674 209820 51750
rect 209884 21418 209912 60030
rect 209964 36576 210016 36582
rect 209964 36518 210016 36524
rect 209872 21412 209924 21418
rect 209872 21354 209924 21360
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209976 6914 210004 36518
rect 211172 10334 211200 60044
rect 211816 57798 211844 60044
rect 212566 60030 212672 60058
rect 211804 57792 211856 57798
rect 211804 57734 211856 57740
rect 212644 33862 212672 60030
rect 212736 60030 213302 60058
rect 212632 33856 212684 33862
rect 212632 33798 212684 33804
rect 211252 29708 211304 29714
rect 211252 29650 211304 29656
rect 211264 16574 211292 29650
rect 211264 16546 211752 16574
rect 211160 10328 211212 10334
rect 211160 10270 211212 10276
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 210004 6914
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207216 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 212736 6186 212764 60030
rect 214024 19990 214052 60044
rect 214656 57792 214708 57798
rect 214656 57734 214708 57740
rect 214564 57724 214616 57730
rect 214564 57666 214616 57672
rect 214012 19984 214064 19990
rect 214012 19926 214064 19932
rect 214576 13598 214604 57666
rect 214668 20194 214696 57734
rect 214760 57594 214788 60044
rect 215312 60030 215510 60058
rect 215864 60030 216246 60058
rect 216876 60030 216982 60058
rect 214748 57588 214800 57594
rect 214748 57530 214800 57536
rect 214748 27056 214800 27062
rect 214748 26998 214800 27004
rect 214656 20188 214708 20194
rect 214656 20130 214708 20136
rect 214564 13592 214616 13598
rect 214564 13534 214616 13540
rect 212724 6180 212776 6186
rect 212724 6122 212776 6128
rect 214472 3596 214524 3602
rect 214472 3538 214524 3544
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213380 480 213408 3470
rect 214484 480 214512 3538
rect 214760 3534 214788 26998
rect 215312 14482 215340 60030
rect 215864 45554 215892 60030
rect 215404 45526 215892 45554
rect 215404 18630 215432 45526
rect 216772 43512 216824 43518
rect 216772 43454 216824 43460
rect 215392 18624 215444 18630
rect 215392 18566 215444 18572
rect 215300 14476 215352 14482
rect 215300 14418 215352 14424
rect 216784 6914 216812 43454
rect 216876 9042 216904 60030
rect 217612 57662 217640 60044
rect 218072 60030 218362 60058
rect 218716 60030 219098 60058
rect 219452 60030 219834 60058
rect 219912 60030 220570 60058
rect 220924 60030 221306 60058
rect 217600 57656 217652 57662
rect 217600 57598 217652 57604
rect 217324 33856 217376 33862
rect 217324 33798 217376 33804
rect 216864 9036 216916 9042
rect 216864 8978 216916 8984
rect 216784 6886 216904 6914
rect 214748 3528 214800 3534
rect 214748 3470 214800 3476
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 215680 480 215708 3470
rect 216876 480 216904 6886
rect 217336 3534 217364 33798
rect 218072 6254 218100 60030
rect 218716 55214 218744 60030
rect 218164 55186 218744 55214
rect 218164 9110 218192 55186
rect 218704 50380 218756 50386
rect 218704 50322 218756 50328
rect 218244 47592 218296 47598
rect 218244 47534 218296 47540
rect 218256 16574 218284 47534
rect 218256 16546 218652 16574
rect 218152 9104 218204 9110
rect 218152 9046 218204 9052
rect 218060 6248 218112 6254
rect 218060 6190 218112 6196
rect 217324 3528 217376 3534
rect 217324 3470 217376 3476
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 218624 3482 218652 16546
rect 218716 3602 218744 50322
rect 219452 12034 219480 60030
rect 219912 45554 219940 60030
rect 220820 47660 220872 47666
rect 220820 47602 220872 47608
rect 219544 45526 219940 45554
rect 219544 17270 219572 45526
rect 219532 17264 219584 17270
rect 219532 17206 219584 17212
rect 220832 16574 220860 47602
rect 220924 21486 220952 60030
rect 222028 57526 222056 60044
rect 222212 60030 222778 60058
rect 222856 60030 223422 60058
rect 222016 57520 222068 57526
rect 222016 57462 222068 57468
rect 220912 21480 220964 21486
rect 220912 21422 220964 21428
rect 220832 16546 221136 16574
rect 219440 12028 219492 12034
rect 219440 11970 219492 11976
rect 219992 11756 220044 11762
rect 219992 11698 220044 11704
rect 218704 3596 218756 3602
rect 218704 3538 218756 3544
rect 218072 480 218100 3470
rect 218624 3454 219296 3482
rect 219268 480 219296 3454
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 11698
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222212 10402 222240 60030
rect 222856 45554 222884 60030
rect 224144 57798 224172 60044
rect 224236 60030 224894 60058
rect 224972 60030 225630 60058
rect 226366 60030 226564 60058
rect 224132 57792 224184 57798
rect 224132 57734 224184 57740
rect 224236 57644 224264 60030
rect 222304 45526 222884 45554
rect 223684 57616 224264 57644
rect 222304 22846 222332 45526
rect 222292 22840 222344 22846
rect 222292 22782 222344 22788
rect 223684 15978 223712 57616
rect 224224 57520 224276 57526
rect 224224 57462 224276 57468
rect 224236 17406 224264 57462
rect 224316 28280 224368 28286
rect 224316 28222 224368 28228
rect 224224 17400 224276 17406
rect 224224 17342 224276 17348
rect 223672 15972 223724 15978
rect 223672 15914 223724 15920
rect 223580 11824 223632 11830
rect 223580 11766 223632 11772
rect 222200 10396 222252 10402
rect 222200 10338 222252 10344
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 222764 480 222792 3470
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 11766
rect 224328 3534 224356 28222
rect 224972 12102 225000 60030
rect 226432 53168 226484 53174
rect 226432 53110 226484 53116
rect 226444 16574 226472 53110
rect 226536 49026 226564 60030
rect 226628 60030 227102 60058
rect 226524 49020 226576 49026
rect 226524 48962 226576 48968
rect 226444 16546 226564 16574
rect 224960 12096 225012 12102
rect 224960 12038 225012 12044
rect 225144 3664 225196 3670
rect 225144 3606 225196 3612
rect 224316 3528 224368 3534
rect 224316 3470 224368 3476
rect 225156 480 225184 3606
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 226536 3482 226564 16546
rect 226628 6322 226656 60030
rect 227720 57656 227772 57662
rect 227720 57598 227772 57604
rect 226984 49088 227036 49094
rect 226984 49030 227036 49036
rect 226616 6316 226668 6322
rect 226616 6258 226668 6264
rect 226996 3602 227024 49030
rect 227732 14550 227760 57598
rect 227824 18698 227852 60044
rect 228192 60030 228574 60058
rect 228192 57662 228220 60030
rect 228180 57656 228232 57662
rect 228180 57598 228232 57604
rect 229100 57656 229152 57662
rect 229100 57598 229152 57604
rect 228364 32496 228416 32502
rect 228364 32438 228416 32444
rect 227812 18692 227864 18698
rect 227812 18634 227864 18640
rect 227720 14544 227772 14550
rect 227720 14486 227772 14492
rect 226984 3596 227036 3602
rect 226984 3538 227036 3544
rect 228376 3534 228404 32438
rect 229112 20058 229140 57598
rect 229204 24206 229232 60044
rect 229664 60030 229954 60058
rect 230492 60030 230690 60058
rect 230768 60030 231426 60058
rect 231964 60030 232162 60058
rect 229664 57662 229692 60030
rect 229652 57656 229704 57662
rect 229652 57598 229704 57604
rect 229192 24200 229244 24206
rect 229192 24142 229244 24148
rect 229100 20052 229152 20058
rect 229100 19994 229152 20000
rect 230492 12170 230520 60030
rect 230768 45554 230796 60030
rect 231124 56976 231176 56982
rect 231124 56918 231176 56924
rect 230584 45526 230796 45554
rect 230584 20126 230612 45526
rect 230572 20120 230624 20126
rect 230572 20062 230624 20068
rect 230480 12164 230532 12170
rect 230480 12106 230532 12112
rect 231032 11892 231084 11898
rect 231032 11834 231084 11840
rect 228732 3596 228784 3602
rect 228732 3538 228784 3544
rect 228364 3528 228416 3534
rect 226352 480 226380 3470
rect 226536 3454 227576 3482
rect 228364 3470 228416 3476
rect 227548 480 227576 3454
rect 228744 480 228772 3538
rect 229836 3324 229888 3330
rect 229836 3266 229888 3272
rect 229848 480 229876 3266
rect 231044 480 231072 11834
rect 231136 4962 231164 56918
rect 231216 37936 231268 37942
rect 231216 37878 231268 37884
rect 231124 4956 231176 4962
rect 231124 4898 231176 4904
rect 231228 3330 231256 37878
rect 231964 9178 231992 60030
rect 232884 56982 232912 60044
rect 233436 60030 233634 60058
rect 233896 60030 234278 60058
rect 234632 60030 235014 60058
rect 235276 60030 235750 60058
rect 236012 60030 236486 60058
rect 236564 60030 237222 60058
rect 237484 60030 237958 60058
rect 238312 60030 238694 60058
rect 233240 57656 233292 57662
rect 233240 57598 233292 57604
rect 232872 56976 232924 56982
rect 232872 56918 232924 56924
rect 233252 9246 233280 57598
rect 233332 49020 233384 49026
rect 233332 48962 233384 48968
rect 233344 16574 233372 48962
rect 233436 22914 233464 60030
rect 233896 57662 233924 60030
rect 233884 57656 233936 57662
rect 233884 57598 233936 57604
rect 233884 56636 233936 56642
rect 233884 56578 233936 56584
rect 233424 22908 233476 22914
rect 233424 22850 233476 22856
rect 233344 16546 233464 16574
rect 233240 9240 233292 9246
rect 233240 9182 233292 9188
rect 231952 9172 232004 9178
rect 231952 9114 232004 9120
rect 232228 3392 232280 3398
rect 232228 3334 232280 3340
rect 231216 3324 231268 3330
rect 231216 3266 231268 3272
rect 232240 480 232268 3334
rect 233436 480 233464 16546
rect 233896 10470 233924 56578
rect 234632 12238 234660 60030
rect 235276 45554 235304 60030
rect 234724 45526 235304 45554
rect 234724 21554 234752 45526
rect 234712 21548 234764 21554
rect 234712 21490 234764 21496
rect 234620 12232 234672 12238
rect 234620 12174 234672 12180
rect 234620 11960 234672 11966
rect 234620 11902 234672 11908
rect 233884 10464 233936 10470
rect 233884 10406 233936 10412
rect 234632 480 234660 11902
rect 236012 9314 236040 60030
rect 236564 45554 236592 60030
rect 237380 57656 237432 57662
rect 237380 57598 237432 57604
rect 236104 45526 236592 45554
rect 236104 25634 236132 45526
rect 236644 43580 236696 43586
rect 236644 43522 236696 43528
rect 236092 25628 236144 25634
rect 236092 25570 236144 25576
rect 236000 9308 236052 9314
rect 236000 9250 236052 9256
rect 236656 3534 236684 43522
rect 236736 35352 236788 35358
rect 236736 35294 236788 35300
rect 236748 3670 236776 35294
rect 237392 21622 237420 57598
rect 237484 25566 237512 60030
rect 238312 57662 238340 60030
rect 238300 57656 238352 57662
rect 238300 57598 238352 57604
rect 239416 56642 239444 60044
rect 239508 60030 240074 60058
rect 240152 60030 240810 60058
rect 239404 56636 239456 56642
rect 239404 56578 239456 56584
rect 238024 50448 238076 50454
rect 238024 50390 238076 50396
rect 237564 29776 237616 29782
rect 237564 29718 237616 29724
rect 237472 25560 237524 25566
rect 237472 25502 237524 25508
rect 237380 21616 237432 21622
rect 237380 21558 237432 21564
rect 237576 16574 237604 29718
rect 237576 16546 237696 16574
rect 236736 3664 236788 3670
rect 236736 3606 236788 3612
rect 235816 3528 235868 3534
rect 235816 3470 235868 3476
rect 236644 3528 236696 3534
rect 236644 3470 236696 3476
rect 235828 480 235856 3470
rect 237012 3392 237064 3398
rect 237012 3334 237064 3340
rect 237024 480 237052 3334
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 237668 354 237696 16546
rect 238036 3398 238064 50390
rect 239508 45554 239536 60030
rect 238864 45526 239536 45554
rect 238864 5030 238892 45526
rect 240152 9382 240180 60030
rect 241532 57526 241560 60044
rect 241624 60030 242282 60058
rect 241520 57520 241572 57526
rect 241520 57462 241572 57468
rect 240784 46300 240836 46306
rect 240784 46242 240836 46248
rect 240140 9376 240192 9382
rect 240140 9318 240192 9324
rect 240508 8968 240560 8974
rect 240508 8910 240560 8916
rect 238852 5024 238904 5030
rect 238852 4966 238904 4972
rect 238024 3392 238076 3398
rect 238024 3334 238076 3340
rect 239312 3324 239364 3330
rect 239312 3266 239364 3272
rect 239324 480 239352 3266
rect 240520 480 240548 8910
rect 240796 3602 240824 46242
rect 240876 39500 240928 39506
rect 240876 39442 240928 39448
rect 240784 3596 240836 3602
rect 240784 3538 240836 3544
rect 240888 3330 240916 39442
rect 241624 18766 241652 60030
rect 242900 57656 242952 57662
rect 242900 57598 242952 57604
rect 241612 18760 241664 18766
rect 241612 18702 241664 18708
rect 242912 6390 242940 57598
rect 243004 22982 243032 60044
rect 243464 60030 243754 60058
rect 244384 60030 244490 60058
rect 244936 60030 245226 60058
rect 243464 57662 243492 60030
rect 243452 57656 243504 57662
rect 243452 57598 243504 57604
rect 244280 57656 244332 57662
rect 244280 57598 244332 57604
rect 242992 22976 243044 22982
rect 242992 22918 243044 22924
rect 242900 6384 242952 6390
rect 242900 6326 242952 6332
rect 244292 5098 244320 57598
rect 244384 7750 244412 60030
rect 244936 57662 244964 60030
rect 244924 57656 244976 57662
rect 244924 57598 244976 57604
rect 245856 57458 245884 60044
rect 245948 60030 246606 60058
rect 247144 60030 247342 60058
rect 247696 60030 248078 60058
rect 248432 60030 248814 60058
rect 249076 60030 249550 60058
rect 245844 57452 245896 57458
rect 245844 57394 245896 57400
rect 244924 54596 244976 54602
rect 244924 54538 244976 54544
rect 244464 28348 244516 28354
rect 244464 28290 244516 28296
rect 244476 16574 244504 28290
rect 244476 16546 244872 16574
rect 244372 7744 244424 7750
rect 244372 7686 244424 7692
rect 244280 5092 244332 5098
rect 244280 5034 244332 5040
rect 241704 4072 241756 4078
rect 241704 4014 241756 4020
rect 240876 3324 240928 3330
rect 240876 3266 240928 3272
rect 241716 480 241744 4014
rect 244096 3596 244148 3602
rect 244096 3538 244148 3544
rect 242900 3256 242952 3262
rect 242900 3198 242952 3204
rect 242912 480 242940 3198
rect 244108 480 244136 3538
rect 244844 3482 244872 16546
rect 244936 3602 244964 54538
rect 245752 40860 245804 40866
rect 245752 40802 245804 40808
rect 245764 6914 245792 40802
rect 245948 16574 245976 60030
rect 247040 57656 247092 57662
rect 247040 57598 247092 57604
rect 246304 57452 246356 57458
rect 246304 57394 246356 57400
rect 246316 18834 246344 57394
rect 246304 18828 246356 18834
rect 246304 18770 246356 18776
rect 245948 16546 246068 16574
rect 245764 6886 245976 6914
rect 244924 3596 244976 3602
rect 244924 3538 244976 3544
rect 244844 3454 245240 3482
rect 245212 480 245240 3454
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 6886
rect 246040 6526 246068 16546
rect 247052 9450 247080 57598
rect 247144 13122 247172 60030
rect 247696 57662 247724 60030
rect 247684 57656 247736 57662
rect 247684 57598 247736 57604
rect 247684 57520 247736 57526
rect 247684 57462 247736 57468
rect 247696 17814 247724 57462
rect 247776 42220 247828 42226
rect 247776 42162 247828 42168
rect 247684 17808 247736 17814
rect 247684 17750 247736 17756
rect 247132 13116 247184 13122
rect 247132 13058 247184 13064
rect 247040 9444 247092 9450
rect 247040 9386 247092 9392
rect 247592 9036 247644 9042
rect 247592 8978 247644 8984
rect 246028 6520 246080 6526
rect 246028 6462 246080 6468
rect 247604 480 247632 8978
rect 247788 3262 247816 42162
rect 248432 6458 248460 60030
rect 249076 45554 249104 60030
rect 250272 57594 250300 60044
rect 250364 60030 251022 60058
rect 250260 57588 250312 57594
rect 250260 57530 250312 57536
rect 250364 45554 250392 60030
rect 250536 57656 250588 57662
rect 250536 57598 250588 57604
rect 248524 45526 249104 45554
rect 249904 45526 250392 45554
rect 248524 13190 248552 45526
rect 248512 13184 248564 13190
rect 248512 13126 248564 13132
rect 249904 6594 249932 45526
rect 250444 45076 250496 45082
rect 250444 45018 250496 45024
rect 249892 6588 249944 6594
rect 249892 6530 249944 6536
rect 248420 6452 248472 6458
rect 248420 6394 248472 6400
rect 250456 3602 250484 45018
rect 250548 16046 250576 57598
rect 251652 57458 251680 60044
rect 251836 60030 252402 60058
rect 251640 57452 251692 57458
rect 251640 57394 251692 57400
rect 251836 45554 251864 60030
rect 253124 57662 253152 60044
rect 253584 60030 253874 60058
rect 254320 60030 254610 60058
rect 253112 57656 253164 57662
rect 253112 57598 253164 57604
rect 253584 45554 253612 60030
rect 254320 57254 254348 60030
rect 255332 57662 255360 60044
rect 255424 60030 256082 60058
rect 256712 60030 256818 60058
rect 256896 60030 257462 60058
rect 254860 57656 254912 57662
rect 254860 57598 254912 57604
rect 255320 57656 255372 57662
rect 255320 57598 255372 57604
rect 254584 57588 254636 57594
rect 254584 57530 254636 57536
rect 254308 57248 254360 57254
rect 254308 57190 254360 57196
rect 251284 45526 251864 45554
rect 252664 45526 253612 45554
rect 250628 33924 250680 33930
rect 250628 33866 250680 33872
rect 250536 16040 250588 16046
rect 250536 15982 250588 15988
rect 250640 4078 250668 33866
rect 251284 24274 251312 45526
rect 251272 24268 251324 24274
rect 251272 24210 251324 24216
rect 252664 13258 252692 45526
rect 253940 19984 253992 19990
rect 253940 19926 253992 19932
rect 253952 16574 253980 19926
rect 253952 16546 254256 16574
rect 252652 13252 252704 13258
rect 252652 13194 252704 13200
rect 251180 9104 251232 9110
rect 251180 9046 251232 9052
rect 250628 4072 250680 4078
rect 250628 4014 250680 4020
rect 250444 3596 250496 3602
rect 250444 3538 250496 3544
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 247776 3256 247828 3262
rect 247776 3198 247828 3204
rect 248788 3120 248840 3126
rect 248788 3062 248840 3068
rect 248800 480 248828 3062
rect 249996 480 250024 3470
rect 251192 480 251220 9046
rect 252376 3664 252428 3670
rect 252376 3606 252428 3612
rect 252388 480 252416 3606
rect 253480 3324 253532 3330
rect 253480 3266 253532 3272
rect 253492 480 253520 3266
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 254596 16182 254624 57530
rect 254676 57452 254728 57458
rect 254676 57394 254728 57400
rect 254688 20534 254716 57394
rect 254768 36644 254820 36650
rect 254768 36586 254820 36592
rect 254676 20528 254728 20534
rect 254676 20470 254728 20476
rect 254584 16176 254636 16182
rect 254584 16118 254636 16124
rect 254780 3534 254808 36586
rect 254872 24342 254900 57598
rect 254860 24336 254912 24342
rect 254860 24278 254912 24284
rect 255424 13326 255452 60030
rect 256712 14618 256740 60030
rect 256896 17338 256924 60030
rect 257344 47728 257396 47734
rect 257344 47670 257396 47676
rect 256884 17332 256936 17338
rect 256884 17274 256936 17280
rect 256700 14612 256752 14618
rect 256700 14554 256752 14560
rect 255412 13320 255464 13326
rect 255412 13262 255464 13268
rect 257068 6180 257120 6186
rect 257068 6122 257120 6128
rect 255872 3596 255924 3602
rect 255872 3538 255924 3544
rect 254768 3528 254820 3534
rect 254768 3470 254820 3476
rect 255884 480 255912 3538
rect 257080 480 257108 6122
rect 257356 3126 257384 47670
rect 258184 13394 258212 60044
rect 258920 57322 258948 60044
rect 259564 60030 259670 60058
rect 260024 60030 260406 60058
rect 260944 60030 261142 60058
rect 261496 60030 261878 60058
rect 262324 60030 262614 60058
rect 259460 57656 259512 57662
rect 259460 57598 259512 57604
rect 258908 57316 258960 57322
rect 258908 57258 258960 57264
rect 258816 57248 258868 57254
rect 258816 57190 258868 57196
rect 258724 55956 258776 55962
rect 258724 55898 258776 55904
rect 258172 13388 258224 13394
rect 258172 13330 258224 13336
rect 258264 9172 258316 9178
rect 258264 9114 258316 9120
rect 257344 3120 257396 3126
rect 257344 3062 257396 3068
rect 258276 480 258304 9114
rect 258736 3330 258764 55898
rect 258828 21962 258856 57190
rect 258816 21956 258868 21962
rect 258816 21898 258868 21904
rect 259472 16574 259500 57598
rect 259564 20262 259592 60030
rect 260024 57662 260052 60030
rect 260012 57656 260064 57662
rect 260012 57598 260064 57604
rect 260840 57656 260892 57662
rect 260840 57598 260892 57604
rect 259644 38004 259696 38010
rect 259644 37946 259696 37952
rect 259552 20256 259604 20262
rect 259552 20198 259604 20204
rect 259472 16546 259592 16574
rect 259564 6662 259592 16546
rect 259552 6656 259604 6662
rect 259552 6598 259604 6604
rect 259656 3482 259684 37946
rect 260852 5166 260880 57598
rect 260944 14686 260972 60030
rect 261496 57662 261524 60030
rect 261484 57656 261536 57662
rect 261484 57598 261536 57604
rect 260932 14680 260984 14686
rect 260932 14622 260984 14628
rect 262324 13462 262352 60030
rect 263244 57594 263272 60044
rect 263612 60030 263994 60058
rect 264072 60030 264730 60058
rect 265084 60030 265466 60058
rect 263232 57588 263284 57594
rect 263232 57530 263284 57536
rect 262312 13456 262364 13462
rect 262312 13398 262364 13404
rect 263612 10538 263640 60030
rect 264072 45554 264100 60030
rect 264244 57112 264296 57118
rect 264244 57054 264296 57060
rect 263704 45526 264100 45554
rect 263704 25702 263732 45526
rect 263692 25696 263744 25702
rect 263692 25638 263744 25644
rect 264256 23050 264284 57054
rect 264336 32564 264388 32570
rect 264336 32506 264388 32512
rect 264244 23044 264296 23050
rect 264244 22986 264296 22992
rect 263600 10532 263652 10538
rect 263600 10474 263652 10480
rect 261760 9240 261812 9246
rect 261760 9182 261812 9188
rect 260840 5160 260892 5166
rect 260840 5102 260892 5108
rect 260656 3732 260708 3738
rect 260656 3674 260708 3680
rect 259472 3454 259684 3482
rect 258724 3324 258776 3330
rect 258724 3266 258776 3272
rect 259472 480 259500 3454
rect 260668 480 260696 3674
rect 261772 480 261800 9182
rect 264348 3602 264376 32506
rect 265084 14754 265112 60030
rect 266188 57118 266216 60044
rect 266464 60030 266938 60058
rect 267016 60030 267674 60058
rect 267752 60030 268318 60058
rect 268580 60030 269054 60058
rect 266176 57112 266228 57118
rect 266176 57054 266228 57060
rect 266360 51876 266412 51882
rect 266360 51818 266412 51824
rect 265072 14748 265124 14754
rect 265072 14690 265124 14696
rect 266372 6914 266400 51818
rect 266464 13530 266492 60030
rect 267016 57610 267044 60030
rect 266556 57582 267044 57610
rect 266556 14822 266584 57582
rect 267004 57316 267056 57322
rect 267004 57258 267056 57264
rect 266544 14816 266596 14822
rect 266544 14758 266596 14764
rect 266452 13524 266504 13530
rect 266452 13466 266504 13472
rect 266372 6886 266584 6914
rect 265348 4140 265400 4146
rect 265348 4082 265400 4088
rect 264336 3596 264388 3602
rect 264336 3538 264388 3544
rect 262956 3528 263008 3534
rect 262956 3470 263008 3476
rect 262968 480 262996 3470
rect 264152 2916 264204 2922
rect 264152 2858 264204 2864
rect 264164 480 264192 2858
rect 265360 480 265388 4082
rect 266556 480 266584 6886
rect 267016 5234 267044 57258
rect 267752 10606 267780 60030
rect 268580 55214 268608 60030
rect 269776 57390 269804 60044
rect 270526 60030 270632 60058
rect 269764 57384 269816 57390
rect 269764 57326 269816 57332
rect 269764 56024 269816 56030
rect 269764 55966 269816 55972
rect 267844 55186 268608 55214
rect 267844 24410 267872 55186
rect 268384 53236 268436 53242
rect 268384 53178 268436 53184
rect 267832 24404 267884 24410
rect 267832 24346 267884 24352
rect 267740 10600 267792 10606
rect 267740 10542 267792 10548
rect 267004 5228 267056 5234
rect 267004 5170 267056 5176
rect 267740 3392 267792 3398
rect 267740 3334 267792 3340
rect 267752 480 267780 3334
rect 268396 2922 268424 53178
rect 268844 4888 268896 4894
rect 268844 4830 268896 4836
rect 268384 2916 268436 2922
rect 268384 2858 268436 2864
rect 268856 480 268884 4830
rect 269776 4146 269804 55966
rect 270604 25770 270632 60030
rect 270696 60030 271262 60058
rect 270592 25764 270644 25770
rect 270592 25706 270644 25712
rect 270696 16114 270724 60030
rect 271144 57384 271196 57390
rect 271144 57326 271196 57332
rect 271156 26042 271184 57326
rect 271144 26036 271196 26042
rect 271144 25978 271196 25984
rect 271236 25560 271288 25566
rect 271236 25502 271288 25508
rect 270684 16108 270736 16114
rect 270684 16050 270736 16056
rect 270776 15904 270828 15910
rect 270776 15846 270828 15852
rect 269764 4140 269816 4146
rect 269764 4082 269816 4088
rect 270040 3596 270092 3602
rect 270040 3538 270092 3544
rect 270052 480 270080 3538
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 354 270816 15846
rect 271248 3398 271276 25502
rect 271984 14890 272012 60044
rect 272720 57322 272748 60044
rect 273456 57526 273484 60044
rect 273548 60030 274114 60058
rect 274652 60030 274850 60058
rect 275204 60030 275586 60058
rect 276124 60030 276322 60058
rect 276768 60030 277058 60058
rect 277504 60030 277794 60058
rect 278240 60030 278530 60058
rect 273444 57520 273496 57526
rect 273444 57462 273496 57468
rect 272708 57316 272760 57322
rect 272708 57258 272760 57264
rect 273352 18624 273404 18630
rect 273352 18566 273404 18572
rect 271972 14884 272024 14890
rect 271972 14826 272024 14832
rect 271236 3392 271288 3398
rect 271236 3334 271288 3340
rect 272432 3324 272484 3330
rect 272432 3266 272484 3272
rect 272444 480 272472 3266
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273364 354 273392 18566
rect 273548 14958 273576 60030
rect 273904 57316 273956 57322
rect 273904 57258 273956 57264
rect 273916 19174 273944 57258
rect 273904 19168 273956 19174
rect 273904 19110 273956 19116
rect 273536 14952 273588 14958
rect 273536 14894 273588 14900
rect 273904 14544 273956 14550
rect 273904 14486 273956 14492
rect 273916 3670 273944 14486
rect 274652 7818 274680 60030
rect 275204 45554 275232 60030
rect 276020 57656 276072 57662
rect 276020 57598 276072 57604
rect 274744 45526 275232 45554
rect 274744 7886 274772 45526
rect 276032 16250 276060 57598
rect 276124 31278 276152 60030
rect 276768 57662 276796 60030
rect 276756 57656 276808 57662
rect 276756 57598 276808 57604
rect 277400 56840 277452 56846
rect 277400 56782 277452 56788
rect 276664 54664 276716 54670
rect 276664 54606 276716 54612
rect 276112 31272 276164 31278
rect 276112 31214 276164 31220
rect 276020 16244 276072 16250
rect 276020 16186 276072 16192
rect 274732 7880 274784 7886
rect 274732 7822 274784 7828
rect 274640 7812 274692 7818
rect 274640 7754 274692 7760
rect 274824 6248 274876 6254
rect 274824 6190 274876 6196
rect 273904 3664 273956 3670
rect 273904 3606 273956 3612
rect 274836 480 274864 6190
rect 276020 3868 276072 3874
rect 276020 3810 276072 3816
rect 276032 480 276060 3810
rect 276676 3738 276704 54606
rect 276756 46368 276808 46374
rect 276756 46310 276808 46316
rect 276664 3732 276716 3738
rect 276664 3674 276716 3680
rect 276768 3330 276796 46310
rect 277412 18902 277440 56782
rect 277504 21758 277532 60030
rect 278044 57656 278096 57662
rect 278044 57598 278096 57604
rect 278056 25838 278084 57598
rect 278240 56846 278268 60030
rect 279252 57662 279280 60044
rect 279436 60030 279910 60058
rect 280264 60030 280646 60058
rect 280724 60030 281382 60058
rect 281552 60030 282118 60058
rect 282380 60030 282854 60058
rect 282932 60030 283590 60058
rect 279240 57656 279292 57662
rect 279240 57598 279292 57604
rect 278228 56840 278280 56846
rect 278228 56782 278280 56788
rect 279436 45554 279464 60030
rect 278884 45526 279464 45554
rect 278044 25832 278096 25838
rect 278044 25774 278096 25780
rect 277492 21752 277544 21758
rect 277492 21694 277544 21700
rect 278044 21412 278096 21418
rect 278044 21354 278096 21360
rect 277400 18896 277452 18902
rect 277400 18838 277452 18844
rect 277952 14476 278004 14482
rect 277952 14418 278004 14424
rect 277124 3664 277176 3670
rect 277124 3606 277176 3612
rect 276756 3324 276808 3330
rect 276756 3266 276808 3272
rect 277136 480 277164 3606
rect 277964 3482 277992 14418
rect 278056 3874 278084 21354
rect 278884 7954 278912 45526
rect 280160 45008 280212 45014
rect 280160 44950 280212 44956
rect 280172 16574 280200 44950
rect 280264 17474 280292 60030
rect 280724 45554 280752 60030
rect 280356 45526 280752 45554
rect 280356 21826 280384 45526
rect 280344 21820 280396 21826
rect 280344 21762 280396 21768
rect 280252 17468 280304 17474
rect 280252 17410 280304 17416
rect 280804 17264 280856 17270
rect 280804 17206 280856 17212
rect 280172 16546 280752 16574
rect 278872 7948 278924 7954
rect 278872 7890 278924 7896
rect 278044 3868 278096 3874
rect 278044 3810 278096 3816
rect 277964 3454 278360 3482
rect 278332 480 278360 3454
rect 279516 3052 279568 3058
rect 279516 2994 279568 3000
rect 279528 480 279556 2994
rect 280724 480 280752 16546
rect 280816 3058 280844 17206
rect 281552 8022 281580 60030
rect 282380 45554 282408 60030
rect 281644 45526 282408 45554
rect 281644 16318 281672 45526
rect 282932 19038 282960 60030
rect 283012 31272 283064 31278
rect 283012 31214 283064 31220
rect 282920 19032 282972 19038
rect 282920 18974 282972 18980
rect 283024 16574 283052 31214
rect 284312 17542 284340 60044
rect 284680 60030 285062 60058
rect 284680 57458 284708 60030
rect 284668 57452 284720 57458
rect 284668 57394 284720 57400
rect 284944 57452 284996 57458
rect 284944 57394 284996 57400
rect 284300 17536 284352 17542
rect 284300 17478 284352 17484
rect 283024 16546 283144 16574
rect 281632 16312 281684 16318
rect 281632 16254 281684 16260
rect 281540 8016 281592 8022
rect 281540 7958 281592 7964
rect 281908 3392 281960 3398
rect 281908 3334 281960 3340
rect 280804 3052 280856 3058
rect 280804 2994 280856 3000
rect 281920 480 281948 3334
rect 283116 480 283144 16546
rect 284956 5302 284984 57394
rect 285036 51944 285088 51950
rect 285036 51886 285088 51892
rect 284944 5296 284996 5302
rect 284944 5238 284996 5244
rect 284300 3800 284352 3806
rect 284300 3742 284352 3748
rect 284312 480 284340 3742
rect 285048 3398 285076 51886
rect 285692 23118 285720 60044
rect 285784 60030 286442 60058
rect 285784 24478 285812 60030
rect 287164 57390 287192 60044
rect 287256 60030 287914 60058
rect 288544 60030 288650 60058
rect 287152 57384 287204 57390
rect 287152 57326 287204 57332
rect 287152 42288 287204 42294
rect 287152 42230 287204 42236
rect 285772 24472 285824 24478
rect 285772 24414 285824 24420
rect 285680 23112 285732 23118
rect 285680 23054 285732 23060
rect 286324 22772 286376 22778
rect 286324 22714 286376 22720
rect 285404 6316 285456 6322
rect 285404 6258 285456 6264
rect 285036 3392 285088 3398
rect 285036 3334 285088 3340
rect 285416 480 285444 6258
rect 286336 3670 286364 22714
rect 287164 16574 287192 42230
rect 287256 17610 287284 60030
rect 287704 57384 287756 57390
rect 287704 57326 287756 57332
rect 287244 17604 287296 17610
rect 287244 17546 287296 17552
rect 287164 16546 287376 16574
rect 286600 9308 286652 9314
rect 286600 9250 286652 9256
rect 286324 3664 286376 3670
rect 286324 3606 286376 3612
rect 286612 480 286640 9250
rect 273598 354 273710 480
rect 273364 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 287716 8090 287744 57326
rect 288544 16386 288572 60030
rect 289372 57390 289400 60044
rect 290016 60030 290122 60058
rect 290568 60030 290858 60058
rect 289820 57656 289872 57662
rect 289820 57598 289872 57604
rect 289360 57384 289412 57390
rect 289360 57326 289412 57332
rect 289832 20330 289860 57598
rect 289912 36712 289964 36718
rect 289912 36654 289964 36660
rect 289820 20324 289872 20330
rect 289820 20266 289872 20272
rect 288532 16380 288584 16386
rect 288532 16322 288584 16328
rect 287704 8084 287756 8090
rect 287704 8026 287756 8032
rect 288992 6384 289044 6390
rect 288992 6326 289044 6332
rect 289004 480 289032 6326
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289924 354 289952 36654
rect 290016 24546 290044 60030
rect 290568 57662 290596 60030
rect 290556 57656 290608 57662
rect 290556 57598 290608 57604
rect 291488 57254 291516 60044
rect 291764 60030 292238 60058
rect 292684 60030 292974 60058
rect 291476 57248 291528 57254
rect 291476 57190 291528 57196
rect 291764 45554 291792 60030
rect 291304 45526 291792 45554
rect 290004 24540 290056 24546
rect 290004 24482 290056 24488
rect 290464 24132 290516 24138
rect 290464 24074 290516 24080
rect 290476 3534 290504 24074
rect 291304 20398 291332 45526
rect 291292 20392 291344 20398
rect 291292 20334 291344 20340
rect 292684 8158 292712 60030
rect 293696 57322 293724 60044
rect 293972 60030 294446 60058
rect 294524 60030 295182 60058
rect 293684 57316 293736 57322
rect 293684 57258 293736 57264
rect 293972 16454 294000 60030
rect 294524 45554 294552 60030
rect 295904 57458 295932 60044
rect 296088 60030 296654 60058
rect 296824 60030 297298 60058
rect 297744 60030 298034 60058
rect 298112 60030 298770 60058
rect 295892 57452 295944 57458
rect 295892 57394 295944 57400
rect 296088 45554 296116 60030
rect 296720 57656 296772 57662
rect 296720 57598 296772 57604
rect 294064 45526 294552 45554
rect 295444 45526 296116 45554
rect 294064 25906 294092 45526
rect 295444 25974 295472 45526
rect 295432 25968 295484 25974
rect 295432 25910 295484 25916
rect 294052 25900 294104 25906
rect 294052 25842 294104 25848
rect 294604 25628 294656 25634
rect 294604 25570 294656 25576
rect 293960 16448 294012 16454
rect 293960 16390 294012 16396
rect 294512 15972 294564 15978
rect 294512 15914 294564 15920
rect 292672 8152 292724 8158
rect 292672 8094 292724 8100
rect 293684 7608 293736 7614
rect 293684 7550 293736 7556
rect 292580 3596 292632 3602
rect 292580 3538 292632 3544
rect 290464 3528 290516 3534
rect 290464 3470 290516 3476
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 291396 480 291424 3470
rect 292592 480 292620 3538
rect 293696 480 293724 7550
rect 294524 3482 294552 15914
rect 294616 3670 294644 25570
rect 296732 17746 296760 57598
rect 296824 21894 296852 60030
rect 297744 57662 297772 60030
rect 297732 57656 297784 57662
rect 297732 57598 297784 57604
rect 297364 38072 297416 38078
rect 297364 38014 297416 38020
rect 296812 21888 296864 21894
rect 296812 21830 296864 21836
rect 296720 17740 296772 17746
rect 296720 17682 296772 17688
rect 294696 13116 294748 13122
rect 294696 13058 294748 13064
rect 294604 3664 294656 3670
rect 294604 3606 294656 3612
rect 294708 3602 294736 13058
rect 297376 4146 297404 38014
rect 298112 17678 298140 60030
rect 298744 53304 298796 53310
rect 298744 53246 298796 53252
rect 298100 17672 298152 17678
rect 298100 17614 298152 17620
rect 297456 13184 297508 13190
rect 297456 13126 297508 13132
rect 296076 4140 296128 4146
rect 296076 4082 296128 4088
rect 297364 4140 297416 4146
rect 297364 4082 297416 4088
rect 294696 3596 294748 3602
rect 294696 3538 294748 3544
rect 294524 3454 294920 3482
rect 294892 480 294920 3454
rect 296088 480 296116 4082
rect 297468 3806 297496 13126
rect 297456 3800 297508 3806
rect 297456 3742 297508 3748
rect 298468 3732 298520 3738
rect 298468 3674 298520 3680
rect 297272 3528 297324 3534
rect 297272 3470 297324 3476
rect 297284 480 297312 3470
rect 298480 480 298508 3674
rect 298756 3534 298784 53246
rect 299492 19106 299520 60044
rect 299584 60030 300242 60058
rect 300872 60030 300978 60058
rect 301056 60030 301714 60058
rect 299584 24614 299612 60030
rect 299572 24608 299624 24614
rect 299572 24550 299624 24556
rect 300872 23186 300900 60030
rect 301056 23322 301084 60030
rect 302240 57656 302292 57662
rect 302240 57598 302292 57604
rect 301044 23316 301096 23322
rect 301044 23258 301096 23264
rect 300860 23180 300912 23186
rect 300860 23122 300912 23128
rect 299480 19100 299532 19106
rect 299480 19042 299532 19048
rect 299480 17332 299532 17338
rect 299480 17274 299532 17280
rect 299492 16574 299520 17274
rect 299492 16546 299704 16574
rect 298744 3528 298796 3534
rect 298744 3470 298796 3476
rect 299676 480 299704 16546
rect 300768 7676 300820 7682
rect 300768 7618 300820 7624
rect 300780 480 300808 7618
rect 301964 3528 302016 3534
rect 301964 3470 302016 3476
rect 301976 480 302004 3470
rect 302252 3466 302280 57598
rect 302344 23254 302372 60044
rect 302712 60030 303094 60058
rect 303724 60030 303830 60058
rect 304184 60030 304566 60058
rect 302712 57662 302740 60030
rect 302700 57656 302752 57662
rect 302700 57598 302752 57604
rect 303620 57656 303672 57662
rect 303620 57598 303672 57604
rect 302332 23248 302384 23254
rect 302332 23190 302384 23196
rect 302332 18692 302384 18698
rect 302332 18634 302384 18640
rect 302344 16574 302372 18634
rect 302344 16546 303200 16574
rect 302240 3460 302292 3466
rect 302240 3402 302292 3408
rect 303172 480 303200 16546
rect 303632 10674 303660 57598
rect 303724 31074 303752 60030
rect 304184 57662 304212 60030
rect 304172 57656 304224 57662
rect 304172 57598 304224 57604
rect 305288 55894 305316 60044
rect 305564 60030 306038 60058
rect 306392 60030 306774 60058
rect 307036 60030 307510 60058
rect 307864 60030 308154 60058
rect 308600 60030 308890 60058
rect 309152 60030 309626 60058
rect 309888 60030 310362 60058
rect 310532 60030 311098 60058
rect 311268 60030 311834 60058
rect 311912 60030 312570 60058
rect 305276 55888 305328 55894
rect 305276 55830 305328 55836
rect 305564 45554 305592 60030
rect 305012 45526 305592 45554
rect 305012 44878 305040 45526
rect 305000 44872 305052 44878
rect 305000 44814 305052 44820
rect 304264 40928 304316 40934
rect 304264 40870 304316 40876
rect 303712 31068 303764 31074
rect 303712 31010 303764 31016
rect 303620 10668 303672 10674
rect 303620 10610 303672 10616
rect 304276 3602 304304 40870
rect 306392 10742 306420 60030
rect 307036 45554 307064 60030
rect 307760 57656 307812 57662
rect 307760 57598 307812 57604
rect 306484 45526 307064 45554
rect 306484 18970 306512 45526
rect 306564 22840 306616 22846
rect 306564 22782 306616 22788
rect 306472 18964 306524 18970
rect 306472 18906 306524 18912
rect 306380 10736 306432 10742
rect 306380 10678 306432 10684
rect 304356 7744 304408 7750
rect 304356 7686 304408 7692
rect 304264 3596 304316 3602
rect 304264 3538 304316 3544
rect 304368 480 304396 7686
rect 305552 3596 305604 3602
rect 305552 3538 305604 3544
rect 305564 480 305592 3538
rect 290158 354 290270 480
rect 289924 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306576 354 306604 22782
rect 307772 10810 307800 57598
rect 307864 42090 307892 60030
rect 308600 57662 308628 60030
rect 308588 57656 308640 57662
rect 308588 57598 308640 57604
rect 308404 55888 308456 55894
rect 308404 55830 308456 55836
rect 307852 42084 307904 42090
rect 307852 42026 307904 42032
rect 307760 10804 307812 10810
rect 307760 10746 307812 10752
rect 307944 7880 307996 7886
rect 307944 7822 307996 7828
rect 307956 480 307984 7822
rect 308416 3738 308444 55830
rect 309152 54534 309180 60030
rect 309140 54528 309192 54534
rect 309140 54470 309192 54476
rect 309140 50516 309192 50522
rect 309140 50458 309192 50464
rect 309152 16574 309180 50458
rect 309888 46238 309916 60030
rect 309876 46232 309928 46238
rect 309876 46174 309928 46180
rect 309152 16546 309824 16574
rect 308404 3732 308456 3738
rect 308404 3674 308456 3680
rect 309048 3460 309100 3466
rect 309048 3402 309100 3408
rect 309060 480 309088 3402
rect 306718 354 306830 480
rect 306576 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 310532 10878 310560 60030
rect 311268 55214 311296 60030
rect 310624 55186 311296 55214
rect 310624 20466 310652 55186
rect 311164 54528 311216 54534
rect 311164 54470 311216 54476
rect 310612 20460 310664 20466
rect 310612 20402 310664 20408
rect 310520 10872 310572 10878
rect 310520 10814 310572 10820
rect 311176 3466 311204 54470
rect 311912 40730 311940 60030
rect 313292 51746 313320 60044
rect 313384 60030 313950 60058
rect 314686 60030 314792 60058
rect 313280 51740 313332 51746
rect 313280 51682 313332 51688
rect 313280 49156 313332 49162
rect 313280 49098 313332 49104
rect 311900 40724 311952 40730
rect 311900 40666 311952 40672
rect 313292 16574 313320 49098
rect 313384 21690 313412 60030
rect 314764 39370 314792 60030
rect 314856 60030 315422 60058
rect 316052 60030 316158 60058
rect 316236 60030 316894 60058
rect 317432 60030 317630 60058
rect 317984 60030 318366 60058
rect 318904 60030 319102 60058
rect 319456 60030 319746 60058
rect 320284 60030 320482 60058
rect 320928 60030 321218 60058
rect 321572 60030 321954 60058
rect 322032 60030 322690 60058
rect 322952 60030 323426 60058
rect 323780 60030 324162 60058
rect 324424 60030 324898 60058
rect 325160 60030 325542 60058
rect 325804 60030 326278 60058
rect 326632 60030 327014 60058
rect 327092 60030 327750 60058
rect 314752 39364 314804 39370
rect 314752 39306 314804 39312
rect 313372 21684 313424 21690
rect 313372 21626 313424 21632
rect 313292 16546 313872 16574
rect 311440 7812 311492 7818
rect 311440 7754 311492 7760
rect 311164 3460 311216 3466
rect 311164 3402 311216 3408
rect 311452 480 311480 7754
rect 312636 3460 312688 3466
rect 312636 3402 312688 3408
rect 312648 480 312676 3402
rect 313844 480 313872 16546
rect 314856 10946 314884 60030
rect 316052 31142 316080 60030
rect 316236 35222 316264 60030
rect 317432 44946 317460 60030
rect 317984 45554 318012 60030
rect 318800 57656 318852 57662
rect 318800 57598 318852 57604
rect 317524 45526 318012 45554
rect 317420 44940 317472 44946
rect 317420 44882 317472 44888
rect 317420 43648 317472 43654
rect 317420 43590 317472 43596
rect 316684 35420 316736 35426
rect 316684 35362 316736 35368
rect 316224 35216 316276 35222
rect 316224 35158 316276 35164
rect 316040 31136 316092 31142
rect 316040 31078 316092 31084
rect 316040 21480 316092 21486
rect 316040 21422 316092 21428
rect 314844 10940 314896 10946
rect 314844 10882 314896 10888
rect 314752 10328 314804 10334
rect 314752 10270 314804 10276
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314764 354 314792 10270
rect 316052 1018 316080 21422
rect 316224 3732 316276 3738
rect 316224 3674 316276 3680
rect 316040 1012 316092 1018
rect 316040 954 316092 960
rect 316236 480 316264 3674
rect 316696 3534 316724 35362
rect 317432 6914 317460 43590
rect 317524 26926 317552 45526
rect 318812 42158 318840 57598
rect 318904 43450 318932 60030
rect 319456 57662 319484 60030
rect 319444 57656 319496 57662
rect 319444 57598 319496 57604
rect 320180 57656 320232 57662
rect 320180 57598 320232 57604
rect 318892 43444 318944 43450
rect 318892 43386 318944 43392
rect 318800 42152 318852 42158
rect 318800 42094 318852 42100
rect 318064 31068 318116 31074
rect 318064 31010 318116 31016
rect 317512 26920 317564 26926
rect 317512 26862 317564 26868
rect 318076 16574 318104 31010
rect 318076 16546 318196 16574
rect 317432 6886 318104 6914
rect 316684 3528 316736 3534
rect 316684 3470 316736 3476
rect 317328 1012 317380 1018
rect 317328 954 317380 960
rect 317340 480 317368 954
rect 314998 354 315110 480
rect 314764 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 6886
rect 318168 3602 318196 16546
rect 320192 5370 320220 57598
rect 320284 32434 320312 60030
rect 320928 57662 320956 60030
rect 320916 57656 320968 57662
rect 320916 57598 320968 57604
rect 321572 40798 321600 60030
rect 322032 53106 322060 60030
rect 322020 53100 322072 53106
rect 322020 53042 322072 53048
rect 321560 40792 321612 40798
rect 321560 40734 321612 40740
rect 320364 32632 320416 32638
rect 320364 32574 320416 32580
rect 320272 32428 320324 32434
rect 320272 32370 320324 32376
rect 320376 16574 320404 32574
rect 320376 16546 320496 16574
rect 320180 5364 320232 5370
rect 320180 5306 320232 5312
rect 319720 3664 319772 3670
rect 319720 3606 319772 3612
rect 318156 3596 318208 3602
rect 318156 3538 318208 3544
rect 319732 480 319760 3606
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322112 7948 322164 7954
rect 322112 7890 322164 7896
rect 322124 480 322152 7890
rect 322952 4826 322980 60030
rect 323780 45554 323808 60030
rect 324320 57656 324372 57662
rect 324320 57598 324372 57604
rect 323044 45526 323808 45554
rect 323044 35290 323072 45526
rect 323032 35284 323084 35290
rect 323032 35226 323084 35232
rect 324332 26994 324360 57598
rect 324424 29646 324452 60030
rect 325160 57662 325188 60030
rect 325148 57656 325200 57662
rect 325148 57598 325200 57604
rect 325700 57656 325752 57662
rect 325700 57598 325752 57604
rect 325712 33794 325740 57598
rect 325804 39438 325832 60030
rect 326632 57662 326660 60030
rect 326620 57656 326672 57662
rect 326620 57598 326672 57604
rect 325792 39432 325844 39438
rect 325792 39374 325844 39380
rect 325700 33788 325752 33794
rect 325700 33730 325752 33736
rect 327092 31210 327120 60030
rect 327724 39432 327776 39438
rect 327724 39374 327776 39380
rect 327080 31204 327132 31210
rect 327080 31146 327132 31152
rect 324412 29640 324464 29646
rect 324412 29582 324464 29588
rect 324320 26988 324372 26994
rect 324320 26930 324372 26936
rect 324964 26988 325016 26994
rect 324964 26930 325016 26936
rect 324320 20052 324372 20058
rect 324320 19994 324372 20000
rect 324332 16574 324360 19994
rect 324332 16546 324452 16574
rect 322940 4820 322992 4826
rect 322940 4762 322992 4768
rect 323308 3528 323360 3534
rect 323308 3470 323360 3476
rect 323320 480 323348 3470
rect 324424 480 324452 16546
rect 324976 3466 325004 26930
rect 327080 26920 327132 26926
rect 327080 26862 327132 26868
rect 327092 16574 327120 26862
rect 327092 16546 327672 16574
rect 325608 8016 325660 8022
rect 325608 7958 325660 7964
rect 324964 3460 325016 3466
rect 324964 3402 325016 3408
rect 325620 480 325648 7958
rect 327644 3482 327672 16546
rect 327736 3738 327764 39374
rect 328472 36582 328500 60044
rect 328564 60030 329222 60058
rect 328564 51814 328592 60030
rect 329840 57656 329892 57662
rect 329840 57598 329892 57604
rect 328552 51808 328604 51814
rect 328552 51750 328604 51756
rect 328460 36576 328512 36582
rect 328460 36518 328512 36524
rect 328460 33788 328512 33794
rect 328460 33730 328512 33736
rect 328472 16574 328500 33730
rect 329852 27062 329880 57598
rect 329944 29714 329972 60044
rect 330312 60030 330602 60058
rect 330312 57662 330340 60030
rect 330300 57656 330352 57662
rect 330300 57598 330352 57604
rect 331220 57656 331272 57662
rect 331220 57598 331272 57604
rect 330484 49224 330536 49230
rect 330484 49166 330536 49172
rect 329932 29708 329984 29714
rect 329932 29650 329984 29656
rect 329840 27056 329892 27062
rect 329840 26998 329892 27004
rect 328472 16546 328776 16574
rect 327724 3732 327776 3738
rect 327724 3674 327776 3680
rect 327644 3454 328040 3482
rect 326804 3392 326856 3398
rect 326804 3334 326856 3340
rect 326816 480 326844 3334
rect 328012 480 328040 3454
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330496 3670 330524 49166
rect 331232 33862 331260 57598
rect 331324 50386 331352 60044
rect 331784 60030 332074 60058
rect 332612 60030 332810 60058
rect 333164 60030 333546 60058
rect 334084 60030 334282 60058
rect 334728 60030 335018 60058
rect 335372 60030 335754 60058
rect 335832 60030 336398 60058
rect 336752 60030 337134 60058
rect 337396 60030 337870 60058
rect 338132 60030 338606 60058
rect 338684 60030 339342 60058
rect 339512 60030 340078 60058
rect 340340 60030 340814 60058
rect 340892 60030 341550 60058
rect 341628 60030 342194 60058
rect 342272 60030 342930 60058
rect 343666 60030 343772 60058
rect 331784 57662 331812 60030
rect 331772 57656 331824 57662
rect 331772 57598 331824 57604
rect 331312 50380 331364 50386
rect 331312 50322 331364 50328
rect 332612 43518 332640 60030
rect 333164 49094 333192 60030
rect 333980 57656 334032 57662
rect 333980 57598 334032 57604
rect 333152 49088 333204 49094
rect 333152 49030 333204 49036
rect 332600 43512 332652 43518
rect 332600 43454 332652 43460
rect 332600 35216 332652 35222
rect 332600 35158 332652 35164
rect 331220 33856 331272 33862
rect 331220 33798 331272 33804
rect 331220 29640 331272 29646
rect 331220 29582 331272 29588
rect 330484 3664 330536 3670
rect 330484 3606 330536 3612
rect 330392 3596 330444 3602
rect 330392 3538 330444 3544
rect 330404 480 330432 3538
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 29582
rect 332612 16574 332640 35158
rect 332612 16546 332732 16574
rect 332704 480 332732 16546
rect 333992 11762 334020 57598
rect 334084 47598 334112 60030
rect 334728 57662 334756 60030
rect 334716 57656 334768 57662
rect 334716 57598 334768 57604
rect 334624 47796 334676 47802
rect 334624 47738 334676 47744
rect 334072 47592 334124 47598
rect 334072 47534 334124 47540
rect 334636 16574 334664 47738
rect 335372 47666 335400 60030
rect 335360 47660 335412 47666
rect 335360 47602 335412 47608
rect 335832 45554 335860 60030
rect 335464 45526 335860 45554
rect 335360 39364 335412 39370
rect 335360 39306 335412 39312
rect 335372 16574 335400 39306
rect 335464 28286 335492 45526
rect 335452 28280 335504 28286
rect 335452 28222 335504 28228
rect 334636 16546 334756 16574
rect 335372 16546 336320 16574
rect 334624 16040 334676 16046
rect 334624 15982 334676 15988
rect 333980 11756 334032 11762
rect 333980 11698 334032 11704
rect 333888 3460 333940 3466
rect 333888 3402 333940 3408
rect 333900 480 333928 3402
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 15982
rect 334728 3398 334756 16546
rect 334716 3392 334768 3398
rect 334716 3334 334768 3340
rect 336292 480 336320 16546
rect 336752 11830 336780 60030
rect 337396 45554 337424 60030
rect 336844 45526 337424 45554
rect 336844 35358 336872 45526
rect 336832 35352 336884 35358
rect 336832 35294 336884 35300
rect 338132 32502 338160 60030
rect 338684 53174 338712 60030
rect 338764 57248 338816 57254
rect 338764 57190 338816 57196
rect 338672 53168 338724 53174
rect 338672 53110 338724 53116
rect 338120 32496 338172 32502
rect 338120 32438 338172 32444
rect 338672 14612 338724 14618
rect 338672 14554 338724 14560
rect 336740 11824 336792 11830
rect 336740 11766 336792 11772
rect 337384 11824 337436 11830
rect 337384 11766 337436 11772
rect 337396 3534 337424 11766
rect 337384 3528 337436 3534
rect 337384 3470 337436 3476
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 337488 480 337516 3470
rect 338684 480 338712 14554
rect 338776 3534 338804 57190
rect 339512 46306 339540 60030
rect 340340 55214 340368 60030
rect 339604 55186 340368 55214
rect 339500 46300 339552 46306
rect 339500 46242 339552 46248
rect 339604 37942 339632 55186
rect 339684 47592 339736 47598
rect 339684 47534 339736 47540
rect 339592 37936 339644 37942
rect 339592 37878 339644 37884
rect 338764 3528 338816 3534
rect 338764 3470 338816 3476
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339696 354 339724 47534
rect 340892 11898 340920 60030
rect 341628 45554 341656 60030
rect 342272 49026 342300 60030
rect 343640 57316 343692 57322
rect 343640 57258 343692 57264
rect 342260 49020 342312 49026
rect 342260 48962 342312 48968
rect 340984 45526 341656 45554
rect 340984 45082 341012 45526
rect 340972 45076 341024 45082
rect 340972 45018 341024 45024
rect 340972 44872 341024 44878
rect 340972 44814 341024 44820
rect 340880 11892 340932 11898
rect 340880 11834 340932 11840
rect 340984 3534 341012 44814
rect 342260 40724 342312 40730
rect 342260 40666 342312 40672
rect 342272 16574 342300 40666
rect 342272 16546 342944 16574
rect 341064 3664 341116 3670
rect 341064 3606 341116 3612
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 341076 1850 341104 3606
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 340984 1822 341104 1850
rect 340984 480 341012 1822
rect 342180 480 342208 3470
rect 339838 354 339950 480
rect 339696 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 343652 6914 343680 57258
rect 343744 11966 343772 60030
rect 343836 60030 344402 60058
rect 343836 43586 343864 60030
rect 345020 57656 345072 57662
rect 345020 57598 345072 57604
rect 343824 43580 343876 43586
rect 343824 43522 343876 43528
rect 345032 29782 345060 57598
rect 345124 50454 345152 60044
rect 345584 60030 345874 60058
rect 345584 57662 345612 60030
rect 345572 57656 345624 57662
rect 345572 57598 345624 57604
rect 346492 57656 346544 57662
rect 346492 57598 346544 57604
rect 346400 54732 346452 54738
rect 346400 54674 346452 54680
rect 345112 50448 345164 50454
rect 345112 50390 345164 50396
rect 345020 29776 345072 29782
rect 345020 29718 345072 29724
rect 343732 11960 343784 11966
rect 343732 11902 343784 11908
rect 345296 11756 345348 11762
rect 345296 11698 345348 11704
rect 343652 6886 344600 6914
rect 344572 480 344600 6886
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 11698
rect 346412 6914 346440 54674
rect 346504 8974 346532 57598
rect 346596 39506 346624 60044
rect 347056 60030 347346 60058
rect 347792 60030 347990 60058
rect 348160 60030 348726 60058
rect 349264 60030 349462 60058
rect 349816 60030 350198 60058
rect 350736 60030 350934 60058
rect 351288 60030 351670 60058
rect 351932 60030 352406 60058
rect 352484 60030 353142 60058
rect 353312 60030 353786 60058
rect 354048 60030 354522 60058
rect 347056 57662 347084 60030
rect 347044 57656 347096 57662
rect 347044 57598 347096 57604
rect 346584 39500 346636 39506
rect 346584 39442 346636 39448
rect 347792 33930 347820 60030
rect 348160 45554 348188 60030
rect 349160 57656 349212 57662
rect 349160 57598 349212 57604
rect 347884 45526 348188 45554
rect 347884 42226 347912 45526
rect 348424 43444 348476 43450
rect 348424 43386 348476 43392
rect 347872 42220 347924 42226
rect 347872 42162 347924 42168
rect 347780 33924 347832 33930
rect 347780 33866 347832 33872
rect 346492 8968 346544 8974
rect 346492 8910 346544 8916
rect 346412 6886 346992 6914
rect 346964 480 346992 6886
rect 348056 3596 348108 3602
rect 348056 3538 348108 3544
rect 348068 480 348096 3538
rect 348436 3534 348464 43386
rect 349172 28354 349200 57598
rect 349264 54602 349292 60030
rect 349816 57662 349844 60030
rect 349804 57656 349856 57662
rect 349804 57598 349856 57604
rect 350632 57656 350684 57662
rect 350632 57598 350684 57604
rect 350540 57384 350592 57390
rect 350540 57326 350592 57332
rect 349252 54596 349304 54602
rect 349252 54538 349304 54544
rect 349160 28348 349212 28354
rect 349160 28290 349212 28296
rect 349160 13252 349212 13258
rect 349160 13194 349212 13200
rect 348424 3528 348476 3534
rect 348424 3470 348476 3476
rect 349172 3346 349200 13194
rect 349252 10396 349304 10402
rect 349252 10338 349304 10344
rect 349264 3534 349292 10338
rect 350552 6914 350580 57326
rect 350644 9042 350672 57598
rect 350736 40866 350764 60030
rect 351288 57662 351316 60030
rect 351276 57656 351328 57662
rect 351276 57598 351328 57604
rect 351932 47734 351960 60030
rect 351920 47728 351972 47734
rect 351920 47670 351972 47676
rect 352484 45554 352512 60030
rect 352024 45526 352512 45554
rect 351920 42084 351972 42090
rect 351920 42026 351972 42032
rect 350724 40860 350776 40866
rect 350724 40802 350776 40808
rect 351932 16574 351960 42026
rect 352024 36650 352052 45526
rect 352012 36644 352064 36650
rect 352012 36586 352064 36592
rect 351932 16546 352880 16574
rect 350632 9036 350684 9042
rect 350632 8978 350684 8984
rect 350552 6886 351224 6914
rect 349252 3528 349304 3534
rect 349252 3470 349304 3476
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 349172 3318 349292 3346
rect 349264 480 349292 3318
rect 350460 480 350488 3470
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 6886
rect 352852 480 352880 16546
rect 353312 9110 353340 60030
rect 353392 46232 353444 46238
rect 353392 46174 353444 46180
rect 353300 9104 353352 9110
rect 353300 9046 353352 9052
rect 353404 6914 353432 46174
rect 354048 45554 354076 60030
rect 355244 55962 355272 60044
rect 355428 60030 355994 60058
rect 356072 60030 356730 60058
rect 355232 55956 355284 55962
rect 355232 55898 355284 55904
rect 355428 45554 355456 60030
rect 353496 45526 354076 45554
rect 354692 45526 355456 45554
rect 353496 14550 353524 45526
rect 354692 19990 354720 45526
rect 356072 32570 356100 60030
rect 356704 37936 356756 37942
rect 356704 37878 356756 37884
rect 356060 32564 356112 32570
rect 356060 32506 356112 32512
rect 354680 19984 354732 19990
rect 354680 19926 354732 19932
rect 353484 14544 353536 14550
rect 353484 14486 353536 14492
rect 353404 6886 353616 6914
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 6886
rect 356336 4820 356388 4826
rect 356336 4762 356388 4768
rect 355232 3596 355284 3602
rect 355232 3538 355284 3544
rect 355244 480 355272 3538
rect 356348 480 356376 4762
rect 356716 3670 356744 37878
rect 357452 6914 357480 60044
rect 357544 60030 358202 60058
rect 358832 60030 358938 60058
rect 359016 60030 359582 60058
rect 357544 9178 357572 60030
rect 358832 38010 358860 60030
rect 359016 54670 359044 60030
rect 359004 54664 359056 54670
rect 359004 54606 359056 54612
rect 360200 51740 360252 51746
rect 360200 51682 360252 51688
rect 358820 38004 358872 38010
rect 358820 37946 358872 37952
rect 357624 18760 357676 18766
rect 357624 18702 357676 18708
rect 357532 9172 357584 9178
rect 357532 9114 357584 9120
rect 357452 6886 357572 6914
rect 357544 6186 357572 6886
rect 357532 6180 357584 6186
rect 357532 6122 357584 6128
rect 356704 3664 356756 3670
rect 356704 3606 356756 3612
rect 357636 3482 357664 18702
rect 359924 8968 359976 8974
rect 359924 8910 359976 8916
rect 358728 3596 358780 3602
rect 358728 3538 358780 3544
rect 357544 3454 357664 3482
rect 357544 480 357572 3454
rect 358740 480 358768 3538
rect 359936 480 359964 8910
rect 360212 6914 360240 51682
rect 360304 9246 360332 60044
rect 360396 60030 361054 60058
rect 361592 60030 361790 60058
rect 360396 24138 360424 60030
rect 361592 53242 361620 60030
rect 362512 56030 362540 60044
rect 363064 60030 363262 60058
rect 363616 60030 363998 60058
rect 364444 60030 364642 60058
rect 364996 60030 365378 60058
rect 365732 60030 366114 60058
rect 366192 60030 366850 60058
rect 367296 60030 367586 60058
rect 368032 60030 368322 60058
rect 368492 60030 369058 60058
rect 369228 60030 369794 60058
rect 369872 60030 370438 60058
rect 370700 60030 371174 60058
rect 371252 60030 371910 60058
rect 372646 60030 372752 60058
rect 362960 57656 363012 57662
rect 362960 57598 363012 57604
rect 362500 56024 362552 56030
rect 362500 55966 362552 55972
rect 361580 53236 361632 53242
rect 361580 53178 361632 53184
rect 362972 25566 363000 57598
rect 363064 51882 363092 60030
rect 363616 57662 363644 60030
rect 363604 57656 363656 57662
rect 363604 57598 363656 57604
rect 364340 55956 364392 55962
rect 364340 55898 364392 55904
rect 363052 51876 363104 51882
rect 363052 51818 363104 51824
rect 362960 25560 363012 25566
rect 362960 25502 363012 25508
rect 363052 25560 363104 25566
rect 363052 25502 363104 25508
rect 360384 24132 360436 24138
rect 360384 24074 360436 24080
rect 360844 21548 360896 21554
rect 360844 21490 360896 21496
rect 360292 9240 360344 9246
rect 360292 9182 360344 9188
rect 360212 6886 360792 6914
rect 360764 3482 360792 6886
rect 360856 3602 360884 21490
rect 363064 16574 363092 25502
rect 363064 16546 363552 16574
rect 362316 3664 362368 3670
rect 362316 3606 362368 3612
rect 360844 3596 360896 3602
rect 360844 3538 360896 3544
rect 360764 3454 361160 3482
rect 361132 480 361160 3454
rect 362328 480 362356 3606
rect 363524 480 363552 16546
rect 364352 3482 364380 55898
rect 364444 4894 364472 60030
rect 364996 45554 365024 60030
rect 364536 45526 365024 45554
rect 364536 25634 364564 45526
rect 364524 25628 364576 25634
rect 364524 25570 364576 25576
rect 365732 15910 365760 60030
rect 366192 46374 366220 60030
rect 367100 57656 367152 57662
rect 367100 57598 367152 57604
rect 366180 46368 366232 46374
rect 366180 46310 366232 46316
rect 365812 33856 365864 33862
rect 365812 33798 365864 33804
rect 365720 15904 365772 15910
rect 365720 15846 365772 15852
rect 364432 4888 364484 4894
rect 364432 4830 364484 4836
rect 364352 3454 364656 3482
rect 364628 480 364656 3454
rect 365824 480 365852 33798
rect 367112 6254 367140 57598
rect 367192 53100 367244 53106
rect 367192 53042 367244 53048
rect 367204 16574 367232 53042
rect 367296 18630 367324 60030
rect 368032 57662 368060 60030
rect 368020 57656 368072 57662
rect 368020 57598 368072 57604
rect 368492 21418 368520 60030
rect 369228 45554 369256 60030
rect 368584 45526 369256 45554
rect 368584 22778 368612 45526
rect 368572 22772 368624 22778
rect 368572 22714 368624 22720
rect 368480 21412 368532 21418
rect 368480 21354 368532 21360
rect 367284 18624 367336 18630
rect 367284 18566 367336 18572
rect 367204 16546 367784 16574
rect 367100 6248 367152 6254
rect 367100 6190 367152 6196
rect 367008 6180 367060 6186
rect 367008 6122 367060 6128
rect 367020 480 367048 6122
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369872 14482 369900 60030
rect 370700 45554 370728 60030
rect 369964 45526 370728 45554
rect 369964 17270 369992 45526
rect 371252 45014 371280 60030
rect 372724 51950 372752 60030
rect 372816 60030 373382 60058
rect 374118 60030 374224 60058
rect 372712 51944 372764 51950
rect 372712 51886 372764 51892
rect 371240 45008 371292 45014
rect 371240 44950 371292 44956
rect 372816 31278 372844 60030
rect 374000 57656 374052 57662
rect 374000 57598 374052 57604
rect 372804 31272 372856 31278
rect 372804 31214 372856 31220
rect 370504 29708 370556 29714
rect 370504 29650 370556 29656
rect 369952 17264 370004 17270
rect 369952 17206 370004 17212
rect 369860 14476 369912 14482
rect 369860 14418 369912 14424
rect 370516 3194 370544 29650
rect 371240 17264 371292 17270
rect 371240 17206 371292 17212
rect 370596 4888 370648 4894
rect 370596 4830 370648 4836
rect 369400 3188 369452 3194
rect 369400 3130 369452 3136
rect 370504 3188 370556 3194
rect 370504 3130 370556 3136
rect 369412 480 369440 3130
rect 370608 480 370636 4830
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 17206
rect 374012 6322 374040 57598
rect 374092 50380 374144 50386
rect 374092 50322 374144 50328
rect 374104 7546 374132 50322
rect 374196 13190 374224 60030
rect 374472 60030 374854 60058
rect 375392 60030 375590 60058
rect 375760 60030 376234 60058
rect 376772 60030 376970 60058
rect 377324 60030 377706 60058
rect 378244 60030 378442 60058
rect 378888 60030 379178 60058
rect 379532 60030 379914 60058
rect 379992 60030 380650 60058
rect 380912 60030 381386 60058
rect 381556 60030 382030 60058
rect 374472 57662 374500 60030
rect 374460 57656 374512 57662
rect 374460 57598 374512 57604
rect 374184 13184 374236 13190
rect 374184 13126 374236 13132
rect 375392 9314 375420 60030
rect 375760 45554 375788 60030
rect 375484 45526 375788 45554
rect 375484 42294 375512 45526
rect 375472 42288 375524 42294
rect 375472 42230 375524 42236
rect 375380 9308 375432 9314
rect 375380 9250 375432 9256
rect 374092 7540 374144 7546
rect 374092 7482 374144 7488
rect 375288 7540 375340 7546
rect 375288 7482 375340 7488
rect 374000 6316 374052 6322
rect 374000 6258 374052 6264
rect 374184 4956 374236 4962
rect 374184 4898 374236 4904
rect 372896 3732 372948 3738
rect 372896 3674 372948 3680
rect 372908 480 372936 3674
rect 374196 2530 374224 4898
rect 374104 2502 374224 2530
rect 374104 480 374132 2502
rect 375300 480 375328 7482
rect 376772 6390 376800 60030
rect 377324 45554 377352 60030
rect 378140 57656 378192 57662
rect 378140 57598 378192 57604
rect 377404 57452 377456 57458
rect 377404 57394 377456 57400
rect 376864 45526 377352 45554
rect 376864 36718 376892 45526
rect 376852 36712 376904 36718
rect 376852 36654 376904 36660
rect 376760 6384 376812 6390
rect 376760 6326 376812 6332
rect 377416 4146 377444 57394
rect 378152 13122 378180 57598
rect 378244 40934 378272 60030
rect 378888 57662 378916 60030
rect 378876 57656 378928 57662
rect 378876 57598 378928 57604
rect 378232 40928 378284 40934
rect 378232 40870 378284 40876
rect 378232 36576 378284 36582
rect 378232 36518 378284 36524
rect 378244 16574 378272 36518
rect 378244 16546 378456 16574
rect 378140 13116 378192 13122
rect 378140 13058 378192 13064
rect 377680 6248 377732 6254
rect 377680 6190 377732 6196
rect 376484 4140 376536 4146
rect 376484 4082 376536 4088
rect 377404 4140 377456 4146
rect 377404 4082 377456 4088
rect 376496 480 376524 4082
rect 377692 480 377720 6190
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379532 7614 379560 60030
rect 379612 51808 379664 51814
rect 379612 51750 379664 51756
rect 379520 7608 379572 7614
rect 379520 7550 379572 7556
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379624 354 379652 51750
rect 379992 45554 380020 60030
rect 379716 45526 380020 45554
rect 379716 15978 379744 45526
rect 380912 38078 380940 60030
rect 381556 53310 381584 60030
rect 382752 55894 382780 60044
rect 383028 60030 383502 60058
rect 383764 60030 384238 60058
rect 384500 60030 384974 60058
rect 385052 60030 385710 60058
rect 386446 60030 386552 60058
rect 382740 55888 382792 55894
rect 382740 55830 382792 55836
rect 381544 53304 381596 53310
rect 381544 53246 381596 53252
rect 383028 45554 383056 60030
rect 383660 55888 383712 55894
rect 383660 55830 383712 55836
rect 382292 45526 383056 45554
rect 380900 38072 380952 38078
rect 380900 38014 380952 38020
rect 382292 17338 382320 45526
rect 382372 31136 382424 31142
rect 382372 31078 382424 31084
rect 382280 17332 382332 17338
rect 382280 17274 382332 17280
rect 379704 15972 379756 15978
rect 379704 15914 379756 15920
rect 381176 6316 381228 6322
rect 381176 6258 381228 6264
rect 381188 480 381216 6258
rect 382384 480 382412 31078
rect 383672 6914 383700 55830
rect 383764 7682 383792 60030
rect 384500 45554 384528 60030
rect 383856 45526 384528 45554
rect 383856 35426 383884 45526
rect 383844 35420 383896 35426
rect 383844 35362 383896 35368
rect 384304 35284 384356 35290
rect 384304 35226 384356 35232
rect 383752 7676 383804 7682
rect 383752 7618 383804 7624
rect 383672 6886 384252 6914
rect 383568 4140 383620 4146
rect 383568 4082 383620 4088
rect 383580 480 383608 4082
rect 384224 490 384252 6886
rect 384316 4146 384344 35226
rect 385052 18698 385080 60030
rect 386420 57520 386472 57526
rect 386420 57462 386472 57468
rect 385132 22772 385184 22778
rect 385132 22714 385184 22720
rect 385040 18692 385092 18698
rect 385040 18634 385092 18640
rect 385144 16574 385172 22714
rect 385144 16546 386000 16574
rect 384304 4140 384356 4146
rect 384304 4082 384356 4088
rect 379950 354 380062 480
rect 379624 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384224 462 384344 490
rect 385972 480 386000 16546
rect 386432 6914 386460 57462
rect 386524 7750 386552 60030
rect 386616 60030 387182 60058
rect 387826 60030 387932 60058
rect 386616 31074 386644 60030
rect 386604 31068 386656 31074
rect 386604 31010 386656 31016
rect 387904 22846 387932 60030
rect 387996 60030 388562 60058
rect 387892 22840 387944 22846
rect 387892 22782 387944 22788
rect 387996 7886 388024 60030
rect 389180 57656 389232 57662
rect 389180 57598 389232 57604
rect 389192 50522 389220 57598
rect 389284 54534 389312 60044
rect 389744 60030 390034 60058
rect 390572 60030 390770 60058
rect 391124 60030 391506 60058
rect 392044 60030 392242 60058
rect 392688 60030 392978 60058
rect 393516 60030 393622 60058
rect 393976 60030 394358 60058
rect 394804 60030 395094 60058
rect 395448 60030 395830 60058
rect 396184 60030 396566 60058
rect 396920 60030 397302 60058
rect 397472 60030 398038 60058
rect 398208 60030 398682 60058
rect 398852 60030 399418 60058
rect 399496 60030 400154 60058
rect 400324 60030 400890 60058
rect 389744 57662 389772 60030
rect 389732 57656 389784 57662
rect 389732 57598 389784 57604
rect 389272 54528 389324 54534
rect 389272 54470 389324 54476
rect 389180 50516 389232 50522
rect 389180 50458 389232 50464
rect 389180 28280 389232 28286
rect 389180 28222 389232 28228
rect 389192 16574 389220 28222
rect 389192 16546 389496 16574
rect 387984 7880 388036 7886
rect 387984 7822 388036 7828
rect 386512 7744 386564 7750
rect 386512 7686 386564 7692
rect 386432 6886 386736 6914
rect 384316 354 384344 462
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 6886
rect 388260 5024 388312 5030
rect 388260 4966 388312 4972
rect 388272 480 388300 4966
rect 389468 480 389496 16546
rect 390572 7818 390600 60030
rect 391124 45554 391152 60030
rect 391940 57656 391992 57662
rect 391940 57598 391992 57604
rect 390664 45526 391152 45554
rect 390664 26994 390692 45526
rect 390652 26988 390704 26994
rect 390652 26930 390704 26936
rect 391952 10334 391980 57598
rect 392044 49162 392072 60030
rect 392688 57662 392716 60030
rect 392676 57656 392728 57662
rect 392676 57598 392728 57604
rect 393412 57656 393464 57662
rect 393412 57598 393464 57604
rect 393320 57588 393372 57594
rect 393320 57530 393372 57536
rect 392032 49156 392084 49162
rect 392032 49098 392084 49104
rect 392032 24132 392084 24138
rect 392032 24074 392084 24080
rect 392044 16574 392072 24074
rect 393332 16574 393360 57530
rect 393424 21486 393452 57598
rect 393516 39438 393544 60030
rect 393976 57662 394004 60030
rect 393964 57656 394016 57662
rect 393964 57598 394016 57604
rect 394700 57656 394752 57662
rect 394700 57598 394752 57604
rect 394712 49230 394740 57598
rect 394700 49224 394752 49230
rect 394700 49166 394752 49172
rect 394700 49020 394752 49026
rect 394700 48962 394752 48968
rect 393504 39432 393556 39438
rect 393504 39374 393556 39380
rect 393412 21480 393464 21486
rect 393412 21422 393464 21428
rect 394712 16574 394740 48962
rect 394804 43654 394832 60030
rect 395448 57662 395476 60030
rect 395436 57656 395488 57662
rect 395436 57598 395488 57604
rect 396080 57656 396132 57662
rect 396080 57598 396132 57604
rect 394792 43648 394844 43654
rect 394792 43590 394844 43596
rect 392044 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 391940 10328 391992 10334
rect 391940 10270 391992 10276
rect 390560 7812 390612 7818
rect 390560 7754 390612 7760
rect 391848 5092 391900 5098
rect 391848 5034 391900 5040
rect 390652 3800 390704 3806
rect 390652 3742 390704 3748
rect 390664 480 390692 3742
rect 391860 480 391888 5034
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 396092 7954 396120 57598
rect 396184 32638 396212 60030
rect 396920 57662 396948 60030
rect 396908 57656 396960 57662
rect 396908 57598 396960 57604
rect 396172 32632 396224 32638
rect 396172 32574 396224 32580
rect 396172 32428 396224 32434
rect 396172 32370 396224 32376
rect 396080 7948 396132 7954
rect 396080 7890 396132 7896
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396184 354 396212 32370
rect 397472 11830 397500 60030
rect 398208 45554 398236 60030
rect 397564 45526 398236 45554
rect 397564 20058 397592 45526
rect 397644 39432 397696 39438
rect 397644 39374 397696 39380
rect 397552 20052 397604 20058
rect 397552 19994 397604 20000
rect 397656 16574 397684 39374
rect 397656 16546 397776 16574
rect 397460 11824 397512 11830
rect 397460 11766 397512 11772
rect 397748 480 397776 16546
rect 398852 8022 398880 60030
rect 399496 47802 399524 60030
rect 400220 57656 400272 57662
rect 400220 57598 400272 57604
rect 399484 47796 399536 47802
rect 399484 47738 399536 47744
rect 400232 16574 400260 57598
rect 400324 26926 400352 60030
rect 401612 33794 401640 60044
rect 401704 60030 402362 60058
rect 402992 60030 403098 60058
rect 403176 60030 403834 60058
rect 404372 60030 404478 60058
rect 404556 60030 405214 60058
rect 405844 60030 405950 60058
rect 401704 43450 401732 60030
rect 401692 43444 401744 43450
rect 401692 43386 401744 43392
rect 401600 33788 401652 33794
rect 401600 33730 401652 33736
rect 402992 29646 403020 60030
rect 403176 35222 403204 60030
rect 403164 35216 403216 35222
rect 403164 35158 403216 35164
rect 402980 29640 403032 29646
rect 402980 29582 403032 29588
rect 400312 26920 400364 26926
rect 400312 26862 400364 26868
rect 402980 19984 403032 19990
rect 402980 19926 403032 19932
rect 402992 16574 403020 19926
rect 400232 16546 400904 16574
rect 402992 16546 403664 16574
rect 398932 15904 398984 15910
rect 398932 15846 398984 15852
rect 398840 8016 398892 8022
rect 398840 7958 398892 7964
rect 398944 3398 398972 15846
rect 399024 5160 399076 5166
rect 399024 5102 399076 5108
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 399036 2666 399064 5102
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398944 2638 399064 2666
rect 398944 480 398972 2638
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396184 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402520 7608 402572 7614
rect 402520 7550 402572 7556
rect 402532 480 402560 7550
rect 403636 480 403664 16546
rect 404372 3466 404400 60030
rect 404556 16046 404584 60030
rect 405740 54528 405792 54534
rect 405740 54470 405792 54476
rect 405752 16574 405780 54470
rect 405844 39370 405872 60030
rect 406672 57254 406700 60044
rect 407316 60030 407422 60058
rect 407776 60030 408158 60058
rect 408512 60030 408894 60058
rect 409156 60030 409630 60058
rect 409984 60030 410274 60058
rect 407212 57724 407264 57730
rect 407212 57666 407264 57672
rect 406660 57248 406712 57254
rect 406660 57190 406712 57196
rect 407120 57248 407172 57254
rect 407120 57190 407172 57196
rect 405832 39364 405884 39370
rect 405832 39306 405884 39312
rect 405752 16546 406056 16574
rect 404544 16040 404596 16046
rect 404544 15982 404596 15988
rect 404360 3460 404412 3466
rect 404360 3402 404412 3408
rect 404820 3460 404872 3466
rect 404820 3402 404872 3408
rect 404832 480 404860 3402
rect 406028 480 406056 16546
rect 407132 3534 407160 57190
rect 407224 47598 407252 57666
rect 407212 47592 407264 47598
rect 407212 47534 407264 47540
rect 407316 14618 407344 60030
rect 407776 57730 407804 60030
rect 407764 57724 407816 57730
rect 407764 57666 407816 57672
rect 407396 47728 407448 47734
rect 407396 47670 407448 47676
rect 407304 14612 407356 14618
rect 407304 14554 407356 14560
rect 407408 6914 407436 47670
rect 408512 37942 408540 60030
rect 409156 45554 409184 60030
rect 408604 45526 409184 45554
rect 408604 44878 408632 45526
rect 408592 44872 408644 44878
rect 408592 44814 408644 44820
rect 409880 44872 409932 44878
rect 409880 44814 409932 44820
rect 408500 37936 408552 37942
rect 408500 37878 408552 37884
rect 409892 16574 409920 44814
rect 409984 40730 410012 60030
rect 410996 57322 411024 60044
rect 411272 60030 411746 60058
rect 411916 60030 412482 60058
rect 410984 57316 411036 57322
rect 410984 57258 411036 57264
rect 410524 56636 410576 56642
rect 410524 56578 410576 56584
rect 409972 40724 410024 40730
rect 409972 40666 410024 40672
rect 409892 16546 410472 16574
rect 409144 10328 409196 10334
rect 409144 10270 409196 10276
rect 407224 6886 407436 6914
rect 407120 3528 407172 3534
rect 407120 3470 407172 3476
rect 407224 480 407252 6886
rect 408408 3528 408460 3534
rect 408408 3470 408460 3476
rect 408420 480 408448 3470
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 10270
rect 409880 3868 409932 3874
rect 409880 3810 409932 3816
rect 409892 3398 409920 3810
rect 410444 3482 410472 16546
rect 410536 3874 410564 56578
rect 411272 11762 411300 60030
rect 411916 54738 411944 60030
rect 413204 56642 413232 60044
rect 413388 60030 413954 60058
rect 414032 60030 414690 60058
rect 413192 56636 413244 56642
rect 413192 56578 413244 56584
rect 411904 54732 411956 54738
rect 411904 54674 411956 54680
rect 412640 53168 412692 53174
rect 412640 53110 412692 53116
rect 411260 11756 411312 11762
rect 411260 11698 411312 11704
rect 410524 3868 410576 3874
rect 410524 3810 410576 3816
rect 411904 3528 411956 3534
rect 410444 3454 410840 3482
rect 411904 3470 411956 3476
rect 409880 3392 409932 3398
rect 409880 3334 409932 3340
rect 410812 480 410840 3454
rect 411916 480 411944 3470
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 53110
rect 413388 45554 413416 60030
rect 412744 45526 413416 45554
rect 412744 13258 412772 45526
rect 412732 13252 412784 13258
rect 412732 13194 412784 13200
rect 414032 10402 414060 60030
rect 415412 57390 415440 60044
rect 415504 60030 416070 60058
rect 416806 60030 416912 60058
rect 415400 57384 415452 57390
rect 415400 57326 415452 57332
rect 414112 43444 414164 43450
rect 414112 43386 414164 43392
rect 414124 16574 414152 43386
rect 415504 42090 415532 60030
rect 416884 46238 416912 60030
rect 417068 60030 417542 60058
rect 418172 60030 418278 60058
rect 418448 60030 419014 60058
rect 419644 60030 419750 60058
rect 420104 60030 420486 60058
rect 421024 60030 421222 60058
rect 421576 60030 421866 60058
rect 422312 60030 422602 60058
rect 416964 46368 417016 46374
rect 416964 46310 417016 46316
rect 416872 46232 416924 46238
rect 416872 46174 416924 46180
rect 415492 42084 415544 42090
rect 415492 42026 415544 42032
rect 415400 21412 415452 21418
rect 415400 21354 415452 21360
rect 415412 16574 415440 21354
rect 414124 16546 414336 16574
rect 415412 16546 415532 16574
rect 414020 10396 414072 10402
rect 414020 10338 414072 10344
rect 414308 480 414336 16546
rect 415504 480 415532 16546
rect 416688 9036 416740 9042
rect 416688 8978 416740 8984
rect 416700 480 416728 8978
rect 416976 490 417004 46310
rect 417068 3602 417096 60030
rect 418172 4826 418200 60030
rect 418344 26920 418396 26926
rect 418344 26862 418396 26868
rect 418356 16574 418384 26862
rect 418448 18766 418476 60030
rect 419540 57724 419592 57730
rect 419540 57666 419592 57672
rect 418436 18760 418488 18766
rect 418436 18702 418488 18708
rect 418356 16546 418568 16574
rect 418160 4820 418212 4826
rect 418160 4762 418212 4768
rect 417056 3596 417108 3602
rect 417056 3538 417108 3544
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 416976 462 417464 490
rect 417436 354 417464 462
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 419552 8974 419580 57666
rect 419644 21554 419672 60030
rect 420104 57730 420132 60030
rect 420092 57724 420144 57730
rect 420092 57666 420144 57672
rect 420920 57724 420972 57730
rect 420920 57666 420972 57672
rect 419632 21548 419684 21554
rect 419632 21490 419684 21496
rect 420184 14476 420236 14482
rect 420184 14418 420236 14424
rect 419540 8968 419592 8974
rect 419540 8910 419592 8916
rect 420196 480 420224 14418
rect 420932 3670 420960 57666
rect 421024 51746 421052 60030
rect 421576 57730 421604 60030
rect 421564 57724 421616 57730
rect 421564 57666 421616 57672
rect 421012 51740 421064 51746
rect 421012 51682 421064 51688
rect 422312 25566 422340 60030
rect 423324 55962 423352 60044
rect 423784 60030 424074 60058
rect 424520 60030 424810 60058
rect 425164 60030 425546 60058
rect 425992 60030 426282 60058
rect 426544 60030 427018 60058
rect 427188 60030 427662 60058
rect 427832 60030 428398 60058
rect 428660 60030 429134 60058
rect 429212 60030 429870 60058
rect 423680 57724 423732 57730
rect 423680 57666 423732 57672
rect 423312 55956 423364 55962
rect 423312 55898 423364 55904
rect 422300 25560 422352 25566
rect 422300 25502 422352 25508
rect 422300 17332 422352 17338
rect 422300 17274 422352 17280
rect 422312 16574 422340 17274
rect 422312 16546 422616 16574
rect 421012 13116 421064 13122
rect 421012 13058 421064 13064
rect 420920 3664 420972 3670
rect 420920 3606 420972 3612
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 421024 354 421052 13058
rect 422588 480 422616 16546
rect 423692 6186 423720 57666
rect 423784 33862 423812 60030
rect 424520 57730 424548 60030
rect 424508 57724 424560 57730
rect 424508 57666 424560 57672
rect 425060 57724 425112 57730
rect 425060 57666 425112 57672
rect 423772 33856 423824 33862
rect 423772 33798 423824 33804
rect 425072 29714 425100 57666
rect 425164 53106 425192 60030
rect 425992 57730 426020 60030
rect 425980 57724 426032 57730
rect 425980 57666 426032 57672
rect 426440 55956 426492 55962
rect 426440 55898 426492 55904
rect 425152 53100 425204 53106
rect 425152 53042 425204 53048
rect 425060 29708 425112 29714
rect 425060 29650 425112 29656
rect 423772 18624 423824 18630
rect 423772 18566 423824 18572
rect 423680 6180 423732 6186
rect 423680 6122 423732 6128
rect 423784 3602 423812 18566
rect 423864 11756 423916 11762
rect 423864 11698 423916 11704
rect 423772 3596 423824 3602
rect 423772 3538 423824 3544
rect 423876 3482 423904 11698
rect 424968 3596 425020 3602
rect 424968 3538 425020 3544
rect 426164 3596 426216 3602
rect 426164 3538 426216 3544
rect 423784 3454 423904 3482
rect 423784 480 423812 3454
rect 424980 480 425008 3538
rect 426176 480 426204 3538
rect 426452 490 426480 55898
rect 426544 4894 426572 60030
rect 427188 45554 427216 60030
rect 426636 45526 427216 45554
rect 426636 17270 426664 45526
rect 426624 17264 426676 17270
rect 426624 17206 426676 17212
rect 426532 4888 426584 4894
rect 426532 4830 426584 4836
rect 427832 3738 427860 60030
rect 428660 45554 428688 60030
rect 429212 50386 429240 60030
rect 430592 57458 430620 60044
rect 430776 60030 431342 60058
rect 431972 60030 432078 60058
rect 432156 60030 432722 60058
rect 433352 60030 433458 60058
rect 433536 60030 434194 60058
rect 434732 60030 434930 60058
rect 430580 57452 430632 57458
rect 430580 57394 430632 57400
rect 430672 51740 430724 51746
rect 430672 51682 430724 51688
rect 429200 50380 429252 50386
rect 429200 50322 429252 50328
rect 427924 45526 428688 45554
rect 427924 4962 427952 45526
rect 428004 42084 428056 42090
rect 428004 42026 428056 42032
rect 428016 16574 428044 42026
rect 429200 29640 429252 29646
rect 429200 29582 429252 29588
rect 428016 16546 428504 16574
rect 427912 4956 427964 4962
rect 427912 4898 427964 4904
rect 427820 3732 427872 3738
rect 427820 3674 427872 3680
rect 421350 354 421462 480
rect 421024 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426452 462 426848 490
rect 428476 480 428504 16546
rect 426820 354 426848 462
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 29582
rect 430684 3482 430712 51682
rect 430776 6254 430804 60030
rect 431972 36582 432000 60030
rect 432156 51814 432184 60030
rect 432144 51808 432196 51814
rect 432144 51750 432196 51756
rect 431960 36576 432012 36582
rect 431960 36518 432012 36524
rect 431960 25560 432012 25566
rect 431960 25502 432012 25508
rect 431972 16574 432000 25502
rect 431972 16546 432092 16574
rect 430764 6248 430816 6254
rect 430764 6190 430816 6196
rect 430684 3454 430896 3482
rect 430868 480 430896 3454
rect 432064 480 432092 16546
rect 433352 6322 433380 60030
rect 433432 50380 433484 50386
rect 433432 50322 433484 50328
rect 433444 6914 433472 50322
rect 433536 31142 433564 60030
rect 434732 35290 434760 60030
rect 435652 55894 435680 60044
rect 436204 60030 436402 60058
rect 436100 57316 436152 57322
rect 436100 57258 436152 57264
rect 435640 55888 435692 55894
rect 435640 55830 435692 55836
rect 434720 35284 434772 35290
rect 434720 35226 434772 35232
rect 433524 31136 433576 31142
rect 433524 31078 433576 31084
rect 433984 31068 434036 31074
rect 433984 31010 434036 31016
rect 433996 16574 434024 31010
rect 436112 16574 436140 57258
rect 436204 22778 436232 60030
rect 437124 57526 437152 60044
rect 437492 60030 437874 60058
rect 437952 60030 438518 60058
rect 437112 57520 437164 57526
rect 437112 57462 437164 57468
rect 436192 22772 436244 22778
rect 436192 22714 436244 22720
rect 433996 16546 434116 16574
rect 436112 16546 436784 16574
rect 433444 6886 434024 6914
rect 433340 6316 433392 6322
rect 433340 6258 433392 6264
rect 433248 2984 433300 2990
rect 433248 2926 433300 2932
rect 433260 480 433288 2926
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 6886
rect 434088 2990 434116 16546
rect 435548 7676 435600 7682
rect 435548 7618 435600 7624
rect 434076 2984 434128 2990
rect 434076 2926 434128 2932
rect 435560 480 435588 7618
rect 436756 480 436784 16546
rect 437492 5030 437520 60030
rect 437952 45554 437980 60030
rect 439240 57730 439268 60044
rect 439516 60030 439990 60058
rect 440344 60030 440726 60058
rect 438124 57724 438176 57730
rect 438124 57666 438176 57672
rect 439228 57724 439280 57730
rect 439228 57666 439280 57672
rect 437584 45526 437980 45554
rect 437584 28286 437612 45526
rect 437572 28280 437624 28286
rect 437572 28222 437624 28228
rect 437940 6180 437992 6186
rect 437940 6122 437992 6128
rect 437480 5024 437532 5030
rect 437480 4966 437532 4972
rect 437952 480 437980 6122
rect 438136 3806 438164 57666
rect 439516 45554 439544 60030
rect 440240 54596 440292 54602
rect 440240 54538 440292 54544
rect 438964 45526 439544 45554
rect 438964 5098 438992 45526
rect 438952 5092 439004 5098
rect 438952 5034 439004 5040
rect 438124 3800 438176 3806
rect 438124 3742 438176 3748
rect 439136 3664 439188 3670
rect 439136 3606 439188 3612
rect 439148 480 439176 3606
rect 440252 3398 440280 54538
rect 440344 24138 440372 60030
rect 441448 57594 441476 60044
rect 441724 60030 442198 60058
rect 442552 60030 442934 60058
rect 443104 60030 443670 60058
rect 444024 60030 444314 60058
rect 444484 60030 445050 60058
rect 441436 57588 441488 57594
rect 441436 57530 441488 57536
rect 441620 57588 441672 57594
rect 441620 57530 441672 57536
rect 440884 57384 440936 57390
rect 440884 57326 440936 57332
rect 440332 24132 440384 24138
rect 440332 24074 440384 24080
rect 440332 22772 440384 22778
rect 440332 22714 440384 22720
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 22714
rect 440896 3670 440924 57326
rect 441632 32434 441660 57530
rect 441724 49026 441752 60030
rect 442552 57594 442580 60030
rect 442540 57588 442592 57594
rect 442540 57530 442592 57536
rect 443000 56636 443052 56642
rect 443000 56578 443052 56584
rect 441712 49020 441764 49026
rect 441712 48962 441764 48968
rect 441620 32428 441672 32434
rect 441620 32370 441672 32376
rect 442632 10396 442684 10402
rect 442632 10338 442684 10344
rect 440884 3664 440936 3670
rect 440884 3606 440936 3612
rect 441620 3596 441672 3602
rect 441620 3538 441672 3544
rect 441632 3398 441660 3538
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441620 3392 441672 3398
rect 441620 3334 441672 3340
rect 441540 480 441568 3334
rect 442644 480 442672 10338
rect 443012 5166 443040 56578
rect 443104 39438 443132 60030
rect 444024 56642 444052 60030
rect 444012 56636 444064 56642
rect 444012 56578 444064 56584
rect 444380 53100 444432 53106
rect 444380 53042 444432 53048
rect 443092 39432 443144 39438
rect 443092 39374 443144 39380
rect 444392 6914 444420 53042
rect 444484 15910 444512 60030
rect 445772 57662 445800 60044
rect 445864 60030 446522 60058
rect 445760 57656 445812 57662
rect 445760 57598 445812 57604
rect 444472 15904 444524 15910
rect 444472 15846 444524 15852
rect 445864 7614 445892 60030
rect 446404 57656 446456 57662
rect 446404 57598 446456 57604
rect 445852 7608 445904 7614
rect 445852 7550 445904 7556
rect 444392 6886 445064 6914
rect 443000 5160 443052 5166
rect 443000 5102 443052 5108
rect 443828 3732 443880 3738
rect 443828 3674 443880 3680
rect 443840 480 443868 3674
rect 445036 480 445064 6886
rect 446220 3528 446272 3534
rect 446220 3470 446272 3476
rect 446232 480 446260 3470
rect 446416 3466 446444 57598
rect 447244 19990 447272 60044
rect 447980 57662 448008 60044
rect 448532 60030 448730 60058
rect 448808 60030 449466 60058
rect 447968 57656 448020 57662
rect 447968 57598 448020 57604
rect 447784 56636 447836 56642
rect 447784 56578 447836 56584
rect 447232 19984 447284 19990
rect 447232 19926 447284 19932
rect 447796 3602 447824 56578
rect 448532 54534 448560 60030
rect 448808 57610 448836 60030
rect 448624 57582 448836 57610
rect 448520 54528 448572 54534
rect 448520 54470 448572 54476
rect 448624 47734 448652 57582
rect 450096 57254 450124 60044
rect 450280 60030 450846 60058
rect 451384 60030 451582 60058
rect 450084 57248 450136 57254
rect 450084 57190 450136 57196
rect 448704 55888 448756 55894
rect 448704 55830 448756 55836
rect 448612 47728 448664 47734
rect 448612 47670 448664 47676
rect 447876 47592 447928 47598
rect 447876 47534 447928 47540
rect 447784 3596 447836 3602
rect 447784 3538 447836 3544
rect 447888 3534 447916 47534
rect 448716 6914 448744 55830
rect 450280 45554 450308 60030
rect 450004 45526 450308 45554
rect 450004 10334 450032 45526
rect 450544 44940 450596 44946
rect 450544 44882 450596 44888
rect 449992 10328 450044 10334
rect 449992 10270 450044 10276
rect 448624 6886 448744 6914
rect 447876 3528 447928 3534
rect 447876 3470 447928 3476
rect 446404 3460 446456 3466
rect 446404 3402 446456 3408
rect 447416 3188 447468 3194
rect 447416 3130 447468 3136
rect 447428 480 447456 3130
rect 448624 480 448652 6886
rect 449808 3664 449860 3670
rect 449808 3606 449860 3612
rect 449820 480 449848 3606
rect 450556 3194 450584 44882
rect 451384 44878 451412 60030
rect 452304 56642 452332 60044
rect 452764 60030 453054 60058
rect 453408 60030 453790 60058
rect 454144 60030 454526 60058
rect 454880 60030 455262 60058
rect 455524 60030 455906 60058
rect 452660 57656 452712 57662
rect 452660 57598 452712 57604
rect 452292 56636 452344 56642
rect 452292 56578 452344 56584
rect 451372 44872 451424 44878
rect 451372 44814 451424 44820
rect 452672 43450 452700 57598
rect 452764 53174 452792 60030
rect 453408 57662 453436 60030
rect 453396 57656 453448 57662
rect 453396 57598 453448 57604
rect 454040 55412 454092 55418
rect 454040 55354 454092 55360
rect 452752 53168 452804 53174
rect 452752 53110 452804 53116
rect 452660 43444 452712 43450
rect 452660 43386 452712 43392
rect 454052 9042 454080 55354
rect 454144 21418 454172 60030
rect 454684 57248 454736 57254
rect 454684 57190 454736 57196
rect 454696 26926 454724 57190
rect 454880 55418 454908 60030
rect 454868 55412 454920 55418
rect 454868 55354 454920 55360
rect 455420 49020 455472 49026
rect 455420 48962 455472 48968
rect 454684 26920 454736 26926
rect 454684 26862 454736 26868
rect 454224 24132 454276 24138
rect 454224 24074 454276 24080
rect 454132 21412 454184 21418
rect 454132 21354 454184 21360
rect 454040 9036 454092 9042
rect 454040 8978 454092 8984
rect 452108 4820 452160 4826
rect 452108 4762 452160 4768
rect 450912 3460 450964 3466
rect 450912 3402 450964 3408
rect 450544 3188 450596 3194
rect 450544 3130 450596 3136
rect 450924 480 450952 3402
rect 452120 480 452148 4762
rect 453304 3392 453356 3398
rect 453304 3334 453356 3340
rect 453316 480 453344 3334
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 434414 -960 434526 326
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454236 354 454264 24074
rect 455432 16574 455460 48962
rect 455524 46374 455552 60030
rect 456628 57254 456656 60044
rect 456996 60030 457378 60058
rect 457824 60030 458114 60058
rect 458192 60030 458850 60058
rect 459586 60030 459692 60058
rect 456616 57248 456668 57254
rect 456616 57190 456668 57196
rect 456800 57248 456852 57254
rect 456800 57190 456852 57196
rect 455512 46368 455564 46374
rect 455512 46310 455564 46316
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3534 456840 57190
rect 456892 55480 456944 55486
rect 456892 55422 456944 55428
rect 456904 13122 456932 55422
rect 456996 14482 457024 60030
rect 457824 55486 457852 60030
rect 457812 55480 457864 55486
rect 457812 55422 457864 55428
rect 458192 17338 458220 60030
rect 458916 57656 458968 57662
rect 458916 57598 458968 57604
rect 458824 57588 458876 57594
rect 458824 57530 458876 57536
rect 458180 17332 458232 17338
rect 458180 17274 458232 17280
rect 456984 14476 457036 14482
rect 456984 14418 457036 14424
rect 456892 13116 456944 13122
rect 456892 13058 456944 13064
rect 456892 3800 456944 3806
rect 456892 3742 456944 3748
rect 456800 3528 456852 3534
rect 456800 3470 456852 3476
rect 456904 480 456932 3742
rect 458836 3738 458864 57530
rect 458928 18630 458956 57598
rect 459560 57452 459612 57458
rect 459560 57394 459612 57400
rect 458916 18624 458968 18630
rect 458916 18566 458968 18572
rect 459192 8968 459244 8974
rect 459192 8910 459244 8916
rect 458824 3732 458876 3738
rect 458824 3674 458876 3680
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 458100 480 458128 3470
rect 459204 480 459232 8910
rect 459572 6914 459600 57394
rect 459664 11762 459692 60030
rect 460308 57662 460336 60044
rect 460296 57656 460348 57662
rect 460296 57598 460348 57604
rect 459652 11756 459704 11762
rect 459652 11698 459704 11704
rect 459572 6886 459968 6914
rect 454470 354 454582 480
rect 454236 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 6886
rect 460952 3602 460980 60044
rect 461688 55962 461716 60044
rect 462320 57656 462372 57662
rect 462320 57598 462372 57604
rect 461676 55956 461728 55962
rect 461676 55898 461728 55904
rect 462332 29646 462360 57598
rect 462424 42090 462452 60044
rect 462792 60030 463174 60058
rect 463804 60030 463910 60058
rect 464264 60030 464646 60058
rect 465092 60030 465382 60058
rect 465552 60030 466118 60058
rect 466564 60030 466762 60058
rect 462792 57662 462820 60030
rect 462780 57656 462832 57662
rect 462780 57598 462832 57604
rect 463700 57656 463752 57662
rect 463700 57598 463752 57604
rect 462412 42084 462464 42090
rect 462412 42026 462464 42032
rect 462320 29640 462372 29646
rect 462320 29582 462372 29588
rect 463712 25566 463740 57598
rect 463804 51746 463832 60030
rect 464264 57662 464292 60030
rect 464252 57656 464304 57662
rect 464252 57598 464304 57604
rect 464344 57656 464396 57662
rect 464344 57598 464396 57604
rect 463792 51740 463844 51746
rect 463792 51682 463844 51688
rect 463700 25560 463752 25566
rect 463700 25502 463752 25508
rect 462780 7608 462832 7614
rect 462780 7550 462832 7556
rect 460940 3596 460992 3602
rect 460940 3538 460992 3544
rect 461584 3596 461636 3602
rect 461584 3538 461636 3544
rect 461596 480 461624 3538
rect 462792 480 462820 7550
rect 464356 3806 464384 57598
rect 465092 31074 465120 60030
rect 465552 50386 465580 60030
rect 465540 50380 465592 50386
rect 465540 50322 465592 50328
rect 465080 31068 465132 31074
rect 465080 31010 465132 31016
rect 466564 7682 466592 60030
rect 467104 57724 467156 57730
rect 467104 57666 467156 57672
rect 466552 7676 466604 7682
rect 466552 7618 466604 7624
rect 466276 6248 466328 6254
rect 466276 6190 466328 6196
rect 464344 3800 464396 3806
rect 464344 3742 464396 3748
rect 465172 3732 465224 3738
rect 465172 3674 465224 3680
rect 463976 3256 464028 3262
rect 463976 3198 464028 3204
rect 463988 480 464016 3198
rect 465184 480 465212 3674
rect 466288 480 466316 6190
rect 467116 3670 467144 57666
rect 467196 57520 467248 57526
rect 467196 57462 467248 57468
rect 467104 3664 467156 3670
rect 467104 3606 467156 3612
rect 467208 3262 467236 57462
rect 467484 57322 467512 60044
rect 467944 60030 468234 60058
rect 467472 57316 467524 57322
rect 467472 57258 467524 57264
rect 467944 6186 467972 60030
rect 468484 57384 468536 57390
rect 468484 57326 468536 57332
rect 467932 6180 467984 6186
rect 467932 6122 467984 6128
rect 468496 3602 468524 57326
rect 468956 57322 468984 60044
rect 469232 60030 469706 60058
rect 469968 60030 470442 60058
rect 470704 60030 471178 60058
rect 468944 57316 468996 57322
rect 468944 57258 468996 57264
rect 469232 22778 469260 60030
rect 469968 54602 469996 60030
rect 470600 57316 470652 57322
rect 470600 57258 470652 57264
rect 469956 54596 470008 54602
rect 469956 54538 470008 54544
rect 469220 22772 469272 22778
rect 469220 22714 469272 22720
rect 469864 4888 469916 4894
rect 469864 4830 469916 4836
rect 468668 3664 468720 3670
rect 468668 3606 468720 3612
rect 467472 3596 467524 3602
rect 467472 3538 467524 3544
rect 468484 3596 468536 3602
rect 468484 3538 468536 3544
rect 467196 3256 467248 3262
rect 467196 3198 467248 3204
rect 467484 480 467512 3538
rect 468680 480 468708 3606
rect 469876 480 469904 4830
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 57258
rect 470704 10402 470732 60030
rect 471244 57792 471296 57798
rect 471244 57734 471296 57740
rect 470692 10396 470744 10402
rect 470692 10338 470744 10344
rect 471256 3534 471284 57734
rect 471900 57594 471928 60044
rect 472084 60030 472558 60058
rect 472912 60030 473294 60058
rect 473464 60030 474030 60058
rect 471888 57588 471940 57594
rect 471888 57530 471940 57536
rect 471980 55616 472032 55622
rect 471980 55558 472032 55564
rect 471992 47598 472020 55558
rect 472084 53106 472112 60030
rect 472912 55622 472940 60030
rect 472900 55616 472952 55622
rect 472900 55558 472952 55564
rect 472072 53100 472124 53106
rect 472072 53042 472124 53048
rect 473360 53100 473412 53106
rect 473360 53042 473412 53048
rect 471980 47592 472032 47598
rect 471980 47534 472032 47540
rect 473372 16574 473400 53042
rect 473464 44946 473492 60030
rect 474004 57656 474056 57662
rect 474004 57598 474056 57604
rect 473452 44940 473504 44946
rect 473452 44882 473504 44888
rect 473372 16546 473492 16574
rect 472256 3596 472308 3602
rect 472256 3538 472308 3544
rect 471244 3528 471296 3534
rect 471244 3470 471296 3476
rect 472268 480 472296 3538
rect 473464 480 473492 16546
rect 473912 10328 473964 10334
rect 473912 10270 473964 10276
rect 473924 490 473952 10270
rect 474016 3466 474044 57598
rect 474752 55894 474780 60044
rect 475488 57730 475516 60044
rect 475476 57724 475528 57730
rect 475476 57666 475528 57672
rect 476224 57662 476252 60044
rect 476316 60030 476974 60058
rect 476212 57656 476264 57662
rect 476212 57598 476264 57604
rect 474740 55888 474792 55894
rect 474740 55830 474792 55836
rect 476212 54528 476264 54534
rect 476212 54470 476264 54476
rect 475752 14476 475804 14482
rect 475752 14418 475804 14424
rect 474004 3460 474056 3466
rect 474004 3402 474056 3408
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 473924 462 474136 490
rect 475764 480 475792 14418
rect 476224 490 476252 54470
rect 476316 4826 476344 60030
rect 477696 57798 477724 60044
rect 478064 60030 478354 60058
rect 478984 60030 479090 60058
rect 477684 57792 477736 57798
rect 477684 57734 477736 57740
rect 477500 57588 477552 57594
rect 477500 57530 477552 57536
rect 476764 56636 476816 56642
rect 476764 56578 476816 56584
rect 476304 4820 476356 4826
rect 476304 4762 476356 4768
rect 476776 3534 476804 56578
rect 477512 6914 477540 57530
rect 478064 45554 478092 60030
rect 478144 57724 478196 57730
rect 478144 57666 478196 57672
rect 477604 45526 478092 45554
rect 477604 24138 477632 45526
rect 477592 24132 477644 24138
rect 477592 24074 477644 24080
rect 478156 16574 478184 57666
rect 478984 49026 479012 60030
rect 479812 57662 479840 60044
rect 479800 57656 479852 57662
rect 479800 57598 479852 57604
rect 480548 57254 480576 60044
rect 480824 60030 481298 60058
rect 480536 57248 480588 57254
rect 480536 57190 480588 57196
rect 478972 49020 479024 49026
rect 478972 48962 479024 48968
rect 480824 45554 480852 60030
rect 480904 57792 480956 57798
rect 480904 57734 480956 57740
rect 480456 45526 480852 45554
rect 478156 16546 478276 16574
rect 477512 6886 478184 6914
rect 476764 3528 476816 3534
rect 476764 3470 476816 3476
rect 474108 354 474136 462
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476224 462 476528 490
rect 478156 480 478184 6886
rect 478248 3738 478276 16546
rect 480456 8974 480484 45526
rect 480536 9036 480588 9042
rect 480536 8978 480588 8984
rect 480444 8968 480496 8974
rect 480444 8910 480496 8916
rect 479340 4140 479392 4146
rect 479340 4082 479392 4088
rect 478236 3732 478288 3738
rect 478236 3674 478288 3680
rect 479352 480 479380 4082
rect 480548 480 480576 8978
rect 480916 3670 480944 57734
rect 482020 57458 482048 60044
rect 482008 57452 482060 57458
rect 482008 57394 482060 57400
rect 482284 57384 482336 57390
rect 482284 57326 482336 57332
rect 482296 4146 482324 57326
rect 482756 56642 482784 60044
rect 483124 60030 483506 60058
rect 482744 56636 482796 56642
rect 482744 56578 482796 56584
rect 483020 55888 483072 55894
rect 483020 55830 483072 55836
rect 483032 6914 483060 55830
rect 483124 7614 483152 60030
rect 484136 57526 484164 60044
rect 484872 57730 484900 60044
rect 484964 60030 485622 60058
rect 484860 57724 484912 57730
rect 484860 57666 484912 57672
rect 484124 57520 484176 57526
rect 484124 57462 484176 57468
rect 484400 57248 484452 57254
rect 484400 57190 484452 57196
rect 483112 7608 483164 7614
rect 483112 7550 483164 7556
rect 483032 6886 484072 6914
rect 482284 4140 482336 4146
rect 482284 4082 482336 4088
rect 480904 3664 480956 3670
rect 480904 3606 480956 3612
rect 481732 3528 481784 3534
rect 481732 3470 481784 3476
rect 481744 480 481772 3470
rect 482836 3392 482888 3398
rect 482836 3334 482888 3340
rect 482848 480 482876 3334
rect 484044 480 484072 6886
rect 484412 490 484440 57190
rect 484964 45554 484992 60030
rect 485044 57452 485096 57458
rect 485044 57394 485096 57400
rect 484504 45526 484992 45554
rect 484504 6254 484532 45526
rect 484492 6248 484544 6254
rect 484492 6190 484544 6196
rect 485056 3534 485084 57394
rect 486344 57322 486372 60044
rect 487080 57798 487108 60044
rect 487172 60030 487830 60058
rect 488566 60030 488672 60058
rect 487068 57792 487120 57798
rect 487068 57734 487120 57740
rect 486424 57656 486476 57662
rect 486424 57598 486476 57604
rect 486332 57316 486384 57322
rect 486332 57258 486384 57264
rect 486436 3602 486464 57598
rect 487172 4894 487200 60030
rect 487804 57724 487856 57730
rect 487804 57666 487856 57672
rect 487252 54596 487304 54602
rect 487252 54538 487304 54544
rect 487160 4888 487212 4894
rect 487160 4830 487212 4836
rect 486424 3596 486476 3602
rect 486424 3538 486476 3544
rect 485044 3528 485096 3534
rect 485044 3470 485096 3476
rect 486424 3460 486476 3466
rect 486424 3402 486476 3408
rect 476500 354 476528 462
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484412 462 484808 490
rect 486436 480 486464 3402
rect 484780 354 484808 462
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487264 354 487292 54538
rect 487816 3398 487844 57666
rect 488540 57520 488592 57526
rect 488540 57462 488592 57468
rect 488552 16574 488580 57462
rect 488644 57186 488672 60030
rect 489288 57662 489316 60044
rect 489276 57656 489328 57662
rect 489276 57598 489328 57604
rect 489368 57656 489420 57662
rect 489368 57598 489420 57604
rect 489380 57458 489408 57598
rect 489368 57452 489420 57458
rect 489368 57394 489420 57400
rect 488632 57180 488684 57186
rect 488632 57122 488684 57128
rect 489932 53106 489960 60044
rect 490024 60030 490682 60058
rect 491312 60030 491418 60058
rect 491496 60030 492154 60058
rect 489920 53100 489972 53106
rect 489920 53042 489972 53048
rect 488552 16546 488856 16574
rect 487804 3392 487856 3398
rect 487804 3334 487856 3340
rect 488828 480 488856 16546
rect 490024 10334 490052 60030
rect 490196 57316 490248 57322
rect 490196 57258 490248 57264
rect 490208 16574 490236 57258
rect 490208 16546 490696 16574
rect 490012 10328 490064 10334
rect 490012 10270 490064 10276
rect 490104 10328 490156 10334
rect 490104 10270 490156 10276
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 354 490002 480
rect 490116 354 490144 10270
rect 489890 326 490144 354
rect 490668 354 490696 16546
rect 491312 14482 491340 60030
rect 491496 54534 491524 60030
rect 492876 57594 492904 60044
rect 492864 57588 492916 57594
rect 492864 57530 492916 57536
rect 493612 57390 493640 60044
rect 494164 60030 494362 60058
rect 494060 57452 494112 57458
rect 494060 57394 494112 57400
rect 493600 57384 493652 57390
rect 493600 57326 493652 57332
rect 491484 54528 491536 54534
rect 491484 54470 491536 54476
rect 491300 14476 491352 14482
rect 491300 14418 491352 14424
rect 494072 6914 494100 57394
rect 494164 9042 494192 60030
rect 494992 57662 495020 60044
rect 495728 57730 495756 60044
rect 495716 57724 495768 57730
rect 495716 57666 495768 57672
rect 494980 57656 495032 57662
rect 494980 57598 495032 57604
rect 496464 55894 496492 60044
rect 496832 60030 497214 60058
rect 497292 60030 497950 60058
rect 498396 60030 498686 60058
rect 496832 57254 496860 60030
rect 497292 57610 497320 60030
rect 496924 57582 497320 57610
rect 496820 57248 496872 57254
rect 496820 57190 496872 57196
rect 496452 55888 496504 55894
rect 496452 55830 496504 55836
rect 494152 9036 494204 9042
rect 494152 8978 494204 8984
rect 494072 6886 494744 6914
rect 492312 4820 492364 4826
rect 492312 4762 492364 4768
rect 492324 480 492352 4762
rect 493508 3596 493560 3602
rect 493508 3538 493560 3544
rect 493520 480 493548 3538
rect 494716 480 494744 6886
rect 495900 6180 495952 6186
rect 495900 6122 495952 6128
rect 495912 480 495940 6122
rect 496924 3466 496952 57582
rect 497004 57520 497056 57526
rect 497004 57462 497056 57468
rect 498292 57520 498344 57526
rect 498292 57462 498344 57468
rect 497016 16574 497044 57462
rect 498200 57248 498252 57254
rect 498200 57190 498252 57196
rect 497016 16546 497136 16574
rect 496912 3460 496964 3466
rect 496912 3402 496964 3408
rect 497108 480 497136 16546
rect 498212 480 498240 57190
rect 498304 16574 498332 57462
rect 498396 54602 498424 60030
rect 499408 57662 499436 60044
rect 499684 60030 500158 60058
rect 499396 57656 499448 57662
rect 499396 57598 499448 57604
rect 498384 54596 498436 54602
rect 498384 54538 498436 54544
rect 498304 16546 498976 16574
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 489890 -960 490002 326
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 499684 10334 499712 60030
rect 500224 57384 500276 57390
rect 500224 57326 500276 57332
rect 499764 56772 499816 56778
rect 499764 56714 499816 56720
rect 499776 16574 499804 56714
rect 499776 16546 500172 16574
rect 499672 10328 499724 10334
rect 499672 10270 499724 10276
rect 500144 3482 500172 16546
rect 500236 3602 500264 57326
rect 500788 57322 500816 60044
rect 501064 60030 501538 60058
rect 500776 57316 500828 57322
rect 500776 57258 500828 57264
rect 501064 4826 501092 60030
rect 502260 57390 502288 60044
rect 502432 57792 502484 57798
rect 502432 57734 502484 57740
rect 502248 57384 502300 57390
rect 502248 57326 502300 57332
rect 502444 16574 502472 57734
rect 502996 57458 503024 60044
rect 503746 60030 503852 60058
rect 503720 57724 503772 57730
rect 503720 57666 503772 57672
rect 502984 57452 503036 57458
rect 502984 57394 503036 57400
rect 502444 16546 503024 16574
rect 501052 4820 501104 4826
rect 501052 4762 501104 4768
rect 500224 3596 500276 3602
rect 500224 3538 500276 3544
rect 501788 3596 501840 3602
rect 501788 3538 501840 3544
rect 500144 3454 500632 3482
rect 500604 480 500632 3454
rect 501800 480 501828 3538
rect 502996 480 503024 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 57666
rect 503824 6186 503852 60030
rect 504468 57594 504496 60044
rect 504456 57588 504508 57594
rect 504456 57530 504508 57536
rect 505204 57254 505232 60044
rect 505284 57656 505336 57662
rect 505284 57598 505336 57604
rect 505192 57248 505244 57254
rect 505192 57190 505244 57196
rect 505296 45554 505324 57598
rect 505940 57526 505968 60044
rect 505928 57520 505980 57526
rect 505928 57462 505980 57468
rect 506584 56778 506612 60044
rect 506768 60030 507334 60058
rect 506572 56772 506624 56778
rect 506572 56714 506624 56720
rect 506480 56704 506532 56710
rect 506480 56646 506532 56652
rect 505112 45526 505324 45554
rect 505112 16574 505140 45526
rect 506492 16574 506520 56646
rect 505112 16546 505416 16574
rect 506492 16546 506704 16574
rect 503812 6180 503864 6186
rect 503812 6122 503864 6128
rect 505388 480 505416 16546
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506492 480 506520 3470
rect 506676 490 506704 16546
rect 506768 3602 506796 60030
rect 508056 57798 508084 60044
rect 508044 57792 508096 57798
rect 508044 57734 508096 57740
rect 508792 57730 508820 60044
rect 508780 57724 508832 57730
rect 508780 57666 508832 57672
rect 509528 57662 509556 60044
rect 509516 57656 509568 57662
rect 509516 57598 509568 57604
rect 509332 57588 509384 57594
rect 509332 57530 509384 57536
rect 508504 56636 508556 56642
rect 508504 56578 508556 56584
rect 506756 3596 506808 3602
rect 506756 3538 506808 3544
rect 508516 3534 508544 56578
rect 509344 45554 509372 57530
rect 510264 56642 510292 60044
rect 510632 60030 511014 60058
rect 511092 60030 511750 60058
rect 510632 56710 510660 60030
rect 511092 57610 511120 60030
rect 510724 57582 511120 57610
rect 512380 57594 512408 60044
rect 512368 57588 512420 57594
rect 510620 56704 510672 56710
rect 510620 56646 510672 56652
rect 510252 56636 510304 56642
rect 510252 56578 510304 56584
rect 509252 45526 509372 45554
rect 509252 16574 509280 45526
rect 509252 16546 509648 16574
rect 508872 3596 508924 3602
rect 508872 3538 508924 3544
rect 508504 3528 508556 3534
rect 508504 3470 508556 3476
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 506676 462 507256 490
rect 508884 480 508912 3538
rect 507228 354 507256 462
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 510724 3602 510752 57582
rect 512368 57530 512420 57536
rect 513116 57526 513144 60044
rect 513484 60030 513866 60058
rect 514312 60030 514602 60058
rect 514864 60030 515338 60058
rect 515784 60030 516074 60058
rect 516152 60030 516810 60058
rect 513380 57656 513432 57662
rect 513380 57598 513432 57604
rect 510804 57520 510856 57526
rect 510804 57462 510856 57468
rect 513104 57520 513156 57526
rect 513104 57462 513156 57468
rect 510816 16574 510844 57462
rect 510816 16546 511304 16574
rect 510712 3596 510764 3602
rect 510712 3538 510764 3544
rect 511276 480 511304 16546
rect 512460 3188 512512 3194
rect 512460 3130 512512 3136
rect 512472 480 512500 3130
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 57598
rect 513484 3194 513512 60030
rect 514312 57662 514340 60030
rect 514300 57656 514352 57662
rect 514300 57598 514352 57604
rect 514760 57656 514812 57662
rect 514760 57598 514812 57604
rect 514772 3534 514800 57598
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 60030
rect 515784 57662 515812 60030
rect 515772 57656 515824 57662
rect 515772 57598 515824 57604
rect 516152 16574 516180 60030
rect 516152 16546 517192 16574
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 513472 3188 513524 3194
rect 513472 3130 513524 3136
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 16546
rect 517532 490 517560 60044
rect 517624 60030 518190 60058
rect 517624 3262 517652 60030
rect 518912 57118 518940 60044
rect 519004 60030 519662 60058
rect 518900 57112 518952 57118
rect 518900 57054 518952 57060
rect 519004 3534 519032 60030
rect 520280 57112 520332 57118
rect 520280 57054 520332 57060
rect 518992 3528 519044 3534
rect 518992 3470 519044 3476
rect 517612 3256 517664 3262
rect 517612 3198 517664 3204
rect 519544 3256 519596 3262
rect 519544 3198 519596 3204
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517532 462 517928 490
rect 519556 480 519584 3198
rect 517900 354 517928 462
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 57054
rect 520384 3194 520412 60044
rect 520476 60030 521134 60058
rect 521672 60030 521870 60058
rect 520476 3262 520504 60030
rect 521672 3466 521700 60030
rect 522592 57730 522620 60044
rect 522580 57724 522632 57730
rect 522580 57666 522632 57672
rect 523328 56846 523356 60044
rect 523512 60030 523986 60058
rect 524524 60030 524722 60058
rect 525168 60030 525458 60058
rect 525812 60030 526194 60058
rect 526364 60030 526930 60058
rect 527376 60030 527666 60058
rect 528112 60030 528402 60058
rect 523316 56840 523368 56846
rect 523316 56782 523368 56788
rect 523512 45554 523540 60030
rect 524420 57656 524472 57662
rect 524420 57598 524472 57604
rect 523052 45526 523540 45554
rect 523052 4078 523080 45526
rect 523040 4072 523092 4078
rect 523040 4014 523092 4020
rect 524432 3534 524460 57598
rect 521844 3528 521896 3534
rect 521844 3470 521896 3476
rect 524420 3528 524472 3534
rect 524420 3470 524472 3476
rect 521660 3460 521712 3466
rect 521660 3402 521712 3408
rect 520464 3256 520516 3262
rect 520464 3198 520516 3204
rect 520372 3188 520424 3194
rect 520372 3130 520424 3136
rect 521856 480 521884 3470
rect 524236 3256 524288 3262
rect 524236 3198 524288 3204
rect 523040 3188 523092 3194
rect 523040 3130 523092 3136
rect 523052 480 523080 3130
rect 524248 480 524276 3198
rect 524524 3194 524552 60030
rect 525168 57662 525196 60030
rect 525156 57656 525208 57662
rect 525156 57598 525208 57604
rect 525812 3874 525840 60030
rect 525892 57724 525944 57730
rect 525892 57666 525944 57672
rect 525800 3868 525852 3874
rect 525800 3810 525852 3816
rect 525432 3460 525484 3466
rect 525432 3402 525484 3408
rect 524512 3188 524564 3194
rect 524512 3130 524564 3136
rect 525444 480 525472 3402
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 525904 354 525932 57666
rect 526364 45554 526392 60030
rect 527180 56840 527232 56846
rect 527180 56782 527232 56788
rect 525996 45526 526392 45554
rect 525996 3670 526024 45526
rect 525984 3664 526036 3670
rect 525984 3606 526036 3612
rect 527192 3482 527220 56782
rect 527272 56296 527324 56302
rect 527272 56238 527324 56244
rect 527284 4146 527312 56238
rect 527272 4140 527324 4146
rect 527272 4082 527324 4088
rect 527376 3738 527404 60030
rect 528112 56302 528140 60030
rect 529032 57390 529060 60044
rect 529768 57594 529796 60044
rect 529952 60030 530518 60058
rect 530596 60030 531254 60058
rect 529756 57588 529808 57594
rect 529756 57530 529808 57536
rect 529020 57384 529072 57390
rect 529020 57326 529072 57332
rect 528100 56296 528152 56302
rect 528100 56238 528152 56244
rect 527916 4140 527968 4146
rect 527916 4082 527968 4088
rect 527364 3732 527416 3738
rect 527364 3674 527416 3680
rect 527192 3454 527864 3482
rect 527928 3466 527956 4082
rect 529020 4072 529072 4078
rect 529020 4014 529072 4020
rect 527836 480 527864 3454
rect 527916 3460 527968 3466
rect 527916 3402 527968 3408
rect 529032 480 529060 4014
rect 529952 3806 529980 60030
rect 530596 57644 530624 60030
rect 530044 57616 530624 57644
rect 530044 18630 530072 57616
rect 530584 57384 530636 57390
rect 530584 57326 530636 57332
rect 530032 18624 530084 18630
rect 530032 18566 530084 18572
rect 529940 3800 529992 3806
rect 529940 3742 529992 3748
rect 530124 3188 530176 3194
rect 530124 3130 530176 3136
rect 530136 480 530164 3130
rect 530596 3058 530624 57326
rect 531976 57118 532004 60044
rect 531964 57112 532016 57118
rect 531964 57054 532016 57060
rect 532712 8974 532740 60044
rect 533448 55894 533476 60044
rect 534080 57656 534132 57662
rect 534080 57598 534132 57604
rect 533436 55888 533488 55894
rect 533436 55830 533488 55836
rect 532700 8968 532752 8974
rect 532700 8910 532752 8916
rect 532516 3868 532568 3874
rect 532516 3810 532568 3816
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 530584 3052 530636 3058
rect 530584 2994 530636 3000
rect 531332 480 531360 3470
rect 532528 480 532556 3810
rect 533712 3664 533764 3670
rect 533712 3606 533764 3612
rect 533724 480 533752 3606
rect 534092 3534 534120 57598
rect 534184 3602 534212 60044
rect 534552 60030 534842 60058
rect 534552 57662 534580 60030
rect 534540 57656 534592 57662
rect 534540 57598 534592 57604
rect 534724 57588 534776 57594
rect 534724 57530 534776 57536
rect 534736 3942 534764 57530
rect 535564 57458 535592 60044
rect 536300 57662 536328 60044
rect 536852 60030 537050 60058
rect 537128 60030 537786 60058
rect 538324 60030 538522 60058
rect 538968 60030 539258 60058
rect 539704 60030 539994 60058
rect 540256 60030 540638 60058
rect 536288 57656 536340 57662
rect 536288 57598 536340 57604
rect 535552 57452 535604 57458
rect 535552 57394 535604 57400
rect 536852 4078 536880 60030
rect 537128 45554 537156 60030
rect 537484 57656 537536 57662
rect 537484 57598 537536 57604
rect 538220 57656 538272 57662
rect 538220 57598 538272 57604
rect 536944 45526 537156 45554
rect 536944 6254 536972 45526
rect 536932 6248 536984 6254
rect 536932 6190 536984 6196
rect 537496 4146 537524 57598
rect 537484 4140 537536 4146
rect 537484 4082 537536 4088
rect 536840 4072 536892 4078
rect 536840 4014 536892 4020
rect 538232 4010 538260 57598
rect 538220 4004 538272 4010
rect 538220 3946 538272 3952
rect 534724 3936 534776 3942
rect 534724 3878 534776 3884
rect 534908 3732 534960 3738
rect 534908 3674 534960 3680
rect 534172 3596 534224 3602
rect 534172 3538 534224 3544
rect 534080 3528 534132 3534
rect 534080 3470 534132 3476
rect 534920 480 534948 3674
rect 536104 3460 536156 3466
rect 536104 3402 536156 3408
rect 536116 480 536144 3402
rect 538324 3398 538352 60030
rect 538968 57662 538996 60030
rect 538956 57656 539008 57662
rect 538956 57598 539008 57604
rect 539600 57656 539652 57662
rect 539600 57598 539652 57604
rect 538864 57112 538916 57118
rect 538864 57054 538916 57060
rect 538404 3936 538456 3942
rect 538404 3878 538456 3884
rect 538312 3392 538364 3398
rect 538312 3334 538364 3340
rect 537208 3052 537260 3058
rect 537208 2994 537260 3000
rect 537220 480 537248 2994
rect 538416 480 538444 3878
rect 538876 3534 538904 57054
rect 539612 3942 539640 57598
rect 539704 4826 539732 60030
rect 540256 57662 540284 60030
rect 541360 57730 541388 60044
rect 541544 60030 542110 60058
rect 541348 57724 541400 57730
rect 541348 57666 541400 57672
rect 540244 57656 540296 57662
rect 540244 57598 540296 57604
rect 541544 45554 541572 60030
rect 542832 57526 542860 60044
rect 542820 57520 542872 57526
rect 542820 57462 542872 57468
rect 543568 57390 543596 60044
rect 543936 60030 544318 60058
rect 544672 60030 545054 60058
rect 543740 57656 543792 57662
rect 543740 57598 543792 57604
rect 543556 57384 543608 57390
rect 543556 57326 543608 57332
rect 540992 45526 541572 45554
rect 539784 18624 539836 18630
rect 539784 18566 539836 18572
rect 539796 16574 539824 18566
rect 539796 16546 540376 16574
rect 539692 4820 539744 4826
rect 539692 4762 539744 4768
rect 539600 3936 539652 3942
rect 539600 3878 539652 3884
rect 539600 3664 539652 3670
rect 539600 3606 539652 3612
rect 538864 3528 538916 3534
rect 538864 3470 538916 3476
rect 539612 480 539640 3606
rect 526598 354 526710 480
rect 525904 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 540992 7614 541020 45526
rect 543188 8968 543240 8974
rect 543188 8910 543240 8916
rect 540980 7608 541032 7614
rect 540980 7550 541032 7556
rect 541992 3528 542044 3534
rect 541992 3470 542044 3476
rect 542004 480 542032 3470
rect 543200 480 543228 8910
rect 543752 3806 543780 57598
rect 543832 55888 543884 55894
rect 543832 55830 543884 55836
rect 543844 6914 543872 55830
rect 543936 14482 543964 60030
rect 544672 57662 544700 60030
rect 544660 57656 544712 57662
rect 544660 57598 544712 57604
rect 545776 57322 545804 60044
rect 545764 57316 545816 57322
rect 545764 57258 545816 57264
rect 546420 55894 546448 60044
rect 546512 60030 547170 60058
rect 546408 55888 546460 55894
rect 546408 55830 546460 55836
rect 543924 14476 543976 14482
rect 543924 14418 543976 14424
rect 543844 6886 544424 6914
rect 543740 3800 543792 3806
rect 543740 3742 543792 3748
rect 544396 480 544424 6886
rect 546512 3874 546540 60030
rect 547144 57452 547196 57458
rect 547144 57394 547196 57400
rect 547156 4894 547184 57394
rect 547892 5250 547920 60044
rect 547984 60030 548642 60058
rect 547984 6186 548012 60030
rect 549364 57458 549392 60044
rect 549732 60030 550114 60058
rect 550744 60030 550850 60058
rect 551296 60030 551586 60058
rect 549352 57452 549404 57458
rect 549352 57394 549404 57400
rect 549732 45554 549760 60030
rect 550640 57656 550692 57662
rect 550640 57598 550692 57604
rect 549272 45526 549760 45554
rect 547972 6180 548024 6186
rect 547972 6122 548024 6128
rect 547892 5222 548012 5250
rect 547144 4888 547196 4894
rect 547144 4830 547196 4836
rect 547880 4888 547932 4894
rect 547880 4830 547932 4836
rect 546500 3868 546552 3874
rect 546500 3810 546552 3816
rect 545488 3596 545540 3602
rect 545488 3538 545540 3544
rect 545500 480 545528 3538
rect 546684 3460 546736 3466
rect 546684 3402 546736 3408
rect 546696 480 546724 3402
rect 547892 480 547920 4830
rect 547984 3738 548012 5222
rect 549076 4140 549128 4146
rect 549076 4082 549128 4088
rect 547972 3732 548024 3738
rect 547972 3674 548024 3680
rect 549088 480 549116 4082
rect 549272 3602 549300 45526
rect 550272 4072 550324 4078
rect 550272 4014 550324 4020
rect 549260 3596 549312 3602
rect 549260 3538 549312 3544
rect 550284 480 550312 4014
rect 550652 3670 550680 57598
rect 550744 8974 550772 60030
rect 551296 57662 551324 60030
rect 551284 57656 551336 57662
rect 551284 57598 551336 57604
rect 552216 57594 552244 60044
rect 552492 60030 552966 60058
rect 553412 60030 553702 60058
rect 553964 60030 554438 60058
rect 554884 60030 555174 60058
rect 555528 60030 555910 60058
rect 552204 57588 552256 57594
rect 552204 57530 552256 57536
rect 552492 54534 552520 60030
rect 552480 54528 552532 54534
rect 552480 54470 552532 54476
rect 550732 8968 550784 8974
rect 550732 8910 550784 8916
rect 551468 6248 551520 6254
rect 551468 6190 551520 6196
rect 550640 3664 550692 3670
rect 550640 3606 550692 3612
rect 551480 480 551508 6190
rect 553412 3534 553440 60030
rect 553964 45554 553992 60030
rect 554780 57656 554832 57662
rect 554780 57598 554832 57604
rect 554792 51746 554820 57598
rect 554884 53106 554912 60030
rect 555528 57662 555556 60030
rect 556344 57724 556396 57730
rect 556344 57666 556396 57672
rect 555516 57656 555568 57662
rect 555516 57598 555568 57604
rect 554872 53100 554924 53106
rect 554872 53042 554924 53048
rect 554780 51740 554832 51746
rect 554780 51682 554832 51688
rect 553504 45526 553992 45554
rect 553400 3528 553452 3534
rect 553400 3470 553452 3476
rect 553504 3466 553532 45526
rect 556356 16574 556384 57666
rect 556632 57254 556660 60044
rect 560956 58682 560984 71810
rect 566476 60722 566504 103770
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 574836 87032 574888 87038
rect 574836 86974 574888 86980
rect 570604 63572 570656 63578
rect 570604 63514 570656 63520
rect 566464 60716 566516 60722
rect 566464 60658 566516 60664
rect 560944 58676 560996 58682
rect 560944 58618 560996 58624
rect 567844 57588 567896 57594
rect 567844 57530 567896 57536
rect 558184 57520 558236 57526
rect 558184 57462 558236 57468
rect 556620 57248 556672 57254
rect 556620 57190 556672 57196
rect 556356 16546 556936 16574
rect 554964 4820 555016 4826
rect 554964 4762 555016 4768
rect 553768 4004 553820 4010
rect 553768 3946 553820 3952
rect 553492 3460 553544 3466
rect 553492 3402 553544 3408
rect 552664 3392 552716 3398
rect 552664 3334 552716 3340
rect 552676 480 552704 3334
rect 553780 480 553808 3946
rect 554976 480 555004 4762
rect 556160 3936 556212 3942
rect 556160 3878 556212 3884
rect 556172 480 556200 3878
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558196 3330 558224 57462
rect 566464 57452 566516 57458
rect 566464 57394 566516 57400
rect 560300 57384 560352 57390
rect 560300 57326 560352 57332
rect 560312 16574 560340 57326
rect 564440 57316 564492 57322
rect 564440 57258 564492 57264
rect 560312 16546 560432 16574
rect 558552 7608 558604 7614
rect 558552 7550 558604 7556
rect 558184 3324 558236 3330
rect 558184 3266 558236 3272
rect 558564 480 558592 7550
rect 559748 3324 559800 3330
rect 559748 3266 559800 3272
rect 559760 480 559788 3266
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 354 560432 16546
rect 562048 14476 562100 14482
rect 562048 14418 562100 14424
rect 562060 480 562088 14418
rect 563244 3800 563296 3806
rect 563244 3742 563296 3748
rect 563256 480 563284 3742
rect 564452 480 564480 57258
rect 564532 55888 564584 55894
rect 564532 55830 564584 55836
rect 564544 16574 564572 55830
rect 564544 16546 565216 16574
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566476 3806 566504 57394
rect 566832 3868 566884 3874
rect 566832 3810 566884 3816
rect 566464 3800 566516 3806
rect 566464 3742 566516 3748
rect 566844 480 566872 3810
rect 567856 2990 567884 57530
rect 570616 6866 570644 63514
rect 574744 54528 574796 54534
rect 574744 54470 574796 54476
rect 572720 8968 572772 8974
rect 572720 8910 572772 8916
rect 570604 6860 570656 6866
rect 570604 6802 570656 6808
rect 569132 6180 569184 6186
rect 569132 6122 569184 6128
rect 568028 3732 568080 3738
rect 568028 3674 568080 3680
rect 567844 2984 567896 2990
rect 567844 2926 567896 2932
rect 568040 480 568068 3674
rect 569144 480 569172 6122
rect 570328 3800 570380 3806
rect 570328 3742 570380 3748
rect 570340 480 570368 3742
rect 571524 3596 571576 3602
rect 571524 3538 571576 3544
rect 571536 480 571564 3538
rect 572732 480 572760 8910
rect 573916 3664 573968 3670
rect 573916 3606 573968 3612
rect 573928 480 573956 3606
rect 574756 3602 574784 54470
rect 574848 46918 574876 86974
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 577504 78736 577556 78742
rect 577504 78678 577556 78684
rect 574836 46912 574888 46918
rect 574836 46854 574888 46860
rect 577516 20670 577544 78678
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580356 58676 580408 58682
rect 580356 58618 580408 58624
rect 578884 53100 578936 53106
rect 578884 53042 578936 53048
rect 577504 20664 577556 20670
rect 577504 20606 577556 20612
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 576308 3596 576360 3602
rect 576308 3538 576360 3544
rect 575112 2984 575164 2990
rect 575112 2926 575164 2932
rect 575124 480 575152 2926
rect 576320 480 576348 3538
rect 578896 3534 578924 53042
rect 580264 51740 580316 51746
rect 580264 51682 580316 51688
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579620 20664 579672 20670
rect 579620 20606 579672 20612
rect 579632 19825 579660 20606
rect 579618 19816 579674 19825
rect 579618 19751 579674 19760
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 577412 3528 577464 3534
rect 577412 3470 577464 3476
rect 578884 3528 578936 3534
rect 578884 3470 578936 3476
rect 577424 480 577452 3470
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 578620 480 578648 3402
rect 580276 3330 580304 51682
rect 580368 33153 580396 58618
rect 582380 57248 582432 57254
rect 582380 57190 582432 57196
rect 580354 33144 580410 33153
rect 580354 33079 580410 33088
rect 582392 16574 582420 57190
rect 582392 16546 583432 16574
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 580264 3324 580316 3330
rect 580264 3266 580316 3272
rect 581012 480 581040 3470
rect 582196 3324 582248 3330
rect 582196 3266 582248 3272
rect 582208 480 582236 3266
rect 583404 480 583432 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 2962 619112 3018 619168
rect 3146 579944 3202 580000
rect 3514 658144 3570 658200
rect 3606 632032 3662 632088
rect 3698 606056 3754 606112
rect 3514 571920 3570 571976
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3054 501744 3110 501800
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 475632 3570 475688
rect 3514 462576 3570 462632
rect 3422 450880 3478 450936
rect 21362 450608 21418 450664
rect 89166 700440 89222 700496
rect 40498 700304 40554 700360
rect 154118 700576 154174 700632
rect 28170 669160 28226 669216
rect 27434 609320 27490 609376
rect 27342 607688 27398 607744
rect 27158 604832 27214 604888
rect 27066 494264 27122 494320
rect 23478 450472 23534 450528
rect 3330 449520 3386 449576
rect 3514 423544 3570 423600
rect 3422 410488 3478 410544
rect 3238 397432 3294 397488
rect 27250 603608 27306 603664
rect 27158 493992 27214 494048
rect 27526 606328 27582 606384
rect 27434 497256 27490 497312
rect 27342 495624 27398 495680
rect 27250 491544 27306 491600
rect 27158 386280 27214 386336
rect 27158 385328 27214 385384
rect 27066 382336 27122 382392
rect 27066 379752 27122 379808
rect 3422 371320 3478 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3238 241032 3294 241088
rect 3330 136720 3386 136776
rect 3698 340040 3754 340096
rect 4066 319232 4122 319288
rect 3974 306176 4030 306232
rect 3882 293120 3938 293176
rect 27526 494264 27582 494320
rect 27526 493992 27582 494048
rect 27526 492768 27582 492824
rect 27434 386280 27490 386336
rect 27342 383696 27398 383752
rect 27250 379616 27306 379672
rect 27158 273264 27214 273320
rect 27066 269048 27122 269104
rect 3790 267144 3846 267200
rect 3698 254088 3754 254144
rect 27434 382336 27490 382392
rect 27342 271632 27398 271688
rect 27250 269048 27306 269104
rect 27158 252592 27214 252648
rect 26974 252456 27030 252512
rect 26974 251504 27030 251560
rect 3606 201864 3662 201920
rect 3974 227024 4030 227080
rect 3790 226888 3846 226944
rect 3974 214920 4030 214976
rect 3882 188808 3938 188864
rect 3790 162832 3846 162888
rect 26974 158344 27030 158400
rect 27526 380840 27582 380896
rect 27526 379752 27582 379808
rect 27526 379616 27582 379672
rect 27434 270272 27490 270328
rect 27342 253816 27398 253872
rect 27158 161336 27214 161392
rect 27158 160112 27214 160168
rect 27526 267552 27582 267608
rect 27434 252456 27490 252512
rect 27434 160112 27490 160168
rect 27342 159704 27398 159760
rect 27250 158344 27306 158400
rect 27066 156848 27122 156904
rect 3698 149776 3754 149832
rect 3514 58520 3570 58576
rect 4066 110608 4122 110664
rect 3882 97552 3938 97608
rect 3790 84632 3846 84688
rect 3698 71576 3754 71632
rect 3606 45464 3662 45520
rect 27158 155624 27214 155680
rect 27066 44920 27122 44976
rect 34518 674908 34520 674928
rect 34520 674908 34572 674928
rect 34572 674908 34574 674928
rect 34518 674872 34574 674908
rect 46202 674908 46204 674928
rect 46204 674908 46256 674928
rect 46256 674908 46258 674928
rect 46202 674872 46258 674908
rect 46938 674892 46994 674928
rect 46938 674872 46940 674892
rect 46940 674872 46992 674892
rect 46992 674872 46994 674892
rect 169022 626864 169078 626920
rect 168562 618160 168618 618216
rect 43074 587832 43130 587888
rect 43534 587832 43590 587888
rect 60646 587832 60702 587888
rect 62946 587832 63002 587888
rect 68926 587832 68982 587888
rect 74446 587832 74502 587888
rect 83830 587832 83886 587888
rect 86406 587832 86462 587888
rect 88246 587832 88302 587888
rect 95238 587832 95294 587888
rect 99194 587832 99250 587888
rect 100574 587832 100630 587888
rect 103150 587832 103206 587888
rect 105082 587832 105138 587888
rect 106278 587832 106334 587888
rect 107750 587832 107806 587888
rect 109498 587832 109554 587888
rect 110510 587832 110566 587888
rect 111614 587832 111670 587888
rect 112534 587832 112590 587888
rect 113086 587832 113142 587888
rect 113822 587832 113878 587888
rect 114834 587832 114890 587888
rect 117134 587832 117190 587888
rect 119802 587832 119858 587888
rect 120262 587832 120318 587888
rect 120538 587832 120594 587888
rect 122654 587832 122710 587888
rect 122838 587832 122894 587888
rect 125046 587832 125102 587888
rect 126886 587832 126942 587888
rect 129370 587832 129426 587888
rect 129646 587832 129702 587888
rect 130566 587832 130622 587888
rect 131118 587832 131174 587888
rect 132590 587832 132646 587888
rect 133142 587832 133198 587888
rect 136454 587832 136510 587888
rect 137926 587832 137982 587888
rect 139306 587832 139362 587888
rect 140134 587832 140190 587888
rect 142710 587832 142766 587888
rect 143446 587832 143502 587888
rect 147678 587832 147734 587888
rect 149518 587832 149574 587888
rect 150714 587832 150770 587888
rect 35714 563100 35770 563136
rect 35714 563080 35716 563100
rect 35716 563080 35768 563100
rect 35768 563080 35770 563100
rect 46754 563100 46810 563136
rect 46754 563080 46756 563100
rect 46756 563080 46808 563100
rect 46808 563080 46810 563100
rect 28814 557096 28870 557152
rect 28262 450744 28318 450800
rect 28722 445168 28778 445224
rect 27526 155624 27582 155680
rect 28538 333104 28594 333160
rect 28630 252320 28686 252376
rect 28446 221176 28502 221232
rect 64878 586472 64934 586528
rect 71686 586336 71742 586392
rect 75826 586336 75882 586392
rect 78586 586336 78642 586392
rect 81346 586336 81402 586392
rect 91006 586336 91062 586392
rect 93766 586336 93822 586392
rect 108946 586336 109002 586392
rect 107750 581712 107806 581768
rect 106278 581576 106334 581632
rect 111614 584432 111670 584488
rect 112534 584296 112590 584352
rect 114374 587696 114430 587752
rect 114558 587696 114614 587752
rect 114374 584568 114430 584624
rect 118606 586336 118662 586392
rect 120170 587696 120226 587752
rect 119802 584704 119858 584760
rect 120262 584840 120318 584896
rect 125506 586336 125562 586392
rect 128266 586336 128322 586392
rect 131026 587696 131082 587752
rect 136546 587016 136602 587072
rect 139030 587036 139086 587072
rect 139030 587016 139032 587036
rect 139032 587016 139084 587036
rect 139084 587016 139086 587036
rect 142066 586336 142122 586392
rect 48042 561720 48098 561776
rect 115478 477808 115534 477864
rect 122654 477808 122710 477864
rect 63406 476040 63462 476096
rect 66166 476040 66222 476096
rect 84106 476040 84162 476096
rect 86866 476040 86922 476096
rect 96526 476040 96582 476096
rect 106186 476040 106242 476096
rect 112994 476040 113050 476096
rect 42798 475516 42854 475552
rect 42798 475496 42800 475516
rect 42800 475496 42852 475516
rect 42852 475496 42854 475516
rect 42798 475380 42854 475416
rect 42798 475360 42800 475380
rect 42800 475360 42852 475380
rect 42852 475360 42854 475380
rect 60646 474836 60702 474872
rect 60646 474816 60648 474836
rect 60648 474816 60700 474836
rect 60700 474816 60702 474836
rect 34518 452512 34574 452568
rect 68926 474816 68982 474872
rect 71686 474816 71742 474872
rect 74446 474816 74502 474872
rect 75826 474816 75882 474872
rect 78586 474816 78642 474872
rect 81346 474816 81402 474872
rect 88246 474816 88302 474872
rect 91006 474816 91062 474872
rect 93766 474816 93822 474872
rect 99286 474816 99342 474872
rect 100666 474816 100722 474872
rect 103426 474816 103482 474872
rect 108854 474952 108910 475008
rect 110326 474972 110382 475008
rect 110326 474952 110328 474972
rect 110328 474952 110380 474972
rect 110380 474952 110382 474972
rect 107566 474816 107622 474872
rect 111614 474952 111670 475008
rect 108946 474816 109002 474872
rect 107566 456184 107622 456240
rect 111706 474816 111762 474872
rect 121182 475496 121238 475552
rect 114374 474952 114430 475008
rect 118606 474952 118662 475008
rect 113086 474816 113142 474872
rect 111706 456048 111762 456104
rect 114466 474816 114522 474872
rect 115754 474816 115810 474872
rect 117226 474816 117282 474872
rect 118514 474816 118570 474872
rect 108946 454688 109002 454744
rect 121366 474952 121422 475008
rect 119986 474816 120042 474872
rect 121274 474816 121330 474872
rect 165434 476176 165490 476232
rect 129554 476040 129610 476096
rect 132406 476040 132462 476096
rect 133786 476040 133842 476096
rect 143354 476040 143410 476096
rect 148322 476040 148378 476096
rect 124034 475768 124090 475824
rect 126886 475244 126942 475280
rect 126886 475224 126888 475244
rect 126888 475224 126940 475244
rect 126940 475224 126942 475244
rect 128266 475108 128322 475144
rect 128266 475088 128268 475108
rect 128268 475088 128320 475108
rect 128320 475088 128322 475108
rect 129646 475360 129702 475416
rect 131026 475224 131082 475280
rect 124126 474816 124182 474872
rect 125506 474816 125562 474872
rect 128266 474816 128322 474872
rect 131026 474816 131082 474872
rect 133694 475088 133750 475144
rect 141790 475768 141846 475824
rect 139306 475224 139362 475280
rect 136454 474952 136510 475008
rect 135166 474816 135222 474872
rect 136362 474816 136418 474872
rect 136546 474816 136602 474872
rect 137926 474816 137982 474872
rect 139214 474816 139270 474872
rect 140686 474816 140742 474872
rect 143446 474816 143502 474872
rect 151358 475496 151414 475552
rect 150346 474816 150402 474872
rect 45650 451868 45652 451888
rect 45652 451868 45704 451888
rect 45704 451868 45706 451888
rect 45650 451832 45706 451868
rect 48042 451288 48098 451344
rect 165434 449928 165490 449984
rect 42890 364248 42946 364304
rect 112994 364248 113050 364304
rect 115754 364248 115810 364304
rect 132958 364248 133014 364304
rect 136546 364248 136602 364304
rect 42798 364112 42854 364168
rect 63406 364112 63462 364168
rect 66166 364112 66222 364168
rect 73158 364112 73214 364168
rect 75826 364112 75882 364168
rect 84106 364112 84162 364168
rect 85670 364112 85726 364168
rect 93766 364112 93822 364168
rect 95606 364112 95662 364168
rect 103150 364112 103206 364168
rect 106186 364112 106242 364168
rect 109590 364112 109646 364168
rect 60646 363024 60702 363080
rect 27434 49408 27490 49464
rect 27342 47776 27398 47832
rect 27250 46416 27306 46472
rect 27158 43696 27214 43752
rect 3422 32408 3478 32464
rect 46938 340720 46994 340776
rect 46202 340212 46204 340232
rect 46204 340212 46256 340232
rect 46256 340212 46258 340232
rect 46202 340176 46258 340212
rect 35162 339532 35164 339552
rect 35164 339532 35216 339552
rect 35216 339532 35218 339552
rect 35162 339496 35218 339532
rect 68926 363024 68982 363080
rect 71686 363024 71742 363080
rect 78586 363024 78642 363080
rect 81346 363024 81402 363080
rect 88246 363024 88302 363080
rect 91006 363024 91062 363080
rect 99286 363024 99342 363080
rect 100666 363024 100722 363080
rect 108854 363296 108910 363352
rect 107566 363024 107622 363080
rect 108946 363024 109002 363080
rect 107566 353232 107622 353288
rect 111614 363160 111670 363216
rect 111706 363024 111762 363080
rect 113086 364112 113142 364168
rect 114466 364112 114522 364168
rect 114374 363024 114430 363080
rect 111706 343576 111762 343632
rect 115846 364112 115902 364168
rect 124034 364112 124090 364168
rect 125966 364112 126022 364168
rect 129554 364112 129610 364168
rect 132038 364112 132094 364168
rect 122746 363840 122802 363896
rect 119986 363296 120042 363352
rect 118514 363160 118570 363216
rect 117226 363024 117282 363080
rect 118606 363024 118662 363080
rect 121274 363160 121330 363216
rect 121182 363024 121238 363080
rect 124126 363432 124182 363488
rect 125506 363160 125562 363216
rect 125414 363024 125470 363080
rect 127622 363976 127678 364032
rect 128266 363704 128322 363760
rect 128174 363024 128230 363080
rect 130934 363160 130990 363216
rect 129646 363024 129702 363080
rect 131026 363024 131082 363080
rect 133142 364112 133198 364168
rect 135902 364112 135958 364168
rect 135166 363704 135222 363760
rect 135166 363024 135222 363080
rect 136546 363840 136602 363896
rect 138294 363432 138350 363488
rect 137926 363024 137982 363080
rect 143354 364248 143410 364304
rect 139214 363024 139270 363080
rect 140318 363024 140374 363080
rect 142066 363024 142122 363080
rect 143446 364112 143502 364168
rect 150346 364112 150402 364168
rect 148966 363024 149022 363080
rect 151174 363568 151230 363624
rect 167274 451868 167276 451888
rect 167276 451868 167328 451888
rect 167328 451868 167330 451888
rect 167274 451832 167330 451868
rect 168378 514936 168434 514992
rect 167734 382336 167790 382392
rect 167182 364148 167184 364168
rect 167184 364148 167236 364168
rect 167236 364148 167238 364168
rect 167182 364112 167238 364148
rect 168194 423544 168250 423600
rect 60646 253680 60702 253736
rect 65706 253680 65762 253736
rect 70674 253680 70730 253736
rect 75550 253680 75606 253736
rect 98274 253680 98330 253736
rect 115662 253716 115664 253736
rect 115664 253716 115716 253736
rect 115716 253716 115718 253736
rect 115662 253680 115718 253716
rect 118330 253680 118386 253736
rect 123022 253680 123078 253736
rect 125506 253700 125562 253736
rect 125506 253680 125508 253700
rect 125508 253680 125560 253700
rect 125560 253680 125562 253700
rect 43350 253544 43406 253600
rect 128082 253680 128138 253736
rect 130566 253544 130622 253600
rect 136454 253544 136510 253600
rect 132958 253408 133014 253464
rect 63406 252456 63462 252512
rect 68190 252456 68246 252512
rect 73158 252456 73214 252512
rect 78126 252456 78182 252512
rect 81254 252456 81310 252512
rect 83554 252456 83610 252512
rect 85670 252456 85726 252512
rect 88246 252456 88302 252512
rect 90822 252456 90878 252512
rect 93214 252456 93270 252512
rect 95606 252456 95662 252512
rect 100574 252456 100630 252512
rect 103150 252456 103206 252512
rect 106094 252456 106150 252512
rect 108486 252456 108542 252512
rect 110510 252456 110566 252512
rect 113086 252456 113142 252512
rect 115846 252456 115902 252512
rect 120906 252456 120962 252512
rect 135994 252456 136050 252512
rect 43350 251368 43406 251424
rect 107566 251232 107622 251288
rect 50342 250416 50398 250472
rect 110326 252320 110382 252376
rect 108946 251232 109002 251288
rect 111706 252320 111762 252376
rect 112994 252320 113050 252376
rect 114466 252320 114522 252376
rect 114374 251912 114430 251968
rect 126886 252320 126942 252376
rect 129554 252320 129610 252376
rect 132038 252320 132094 252376
rect 133786 252320 133842 252376
rect 121182 251640 121238 251696
rect 117226 251232 117282 251288
rect 118606 251232 118662 251288
rect 119986 251232 120042 251288
rect 121274 251232 121330 251288
rect 122746 251232 122802 251288
rect 124126 251232 124182 251288
rect 125506 251232 125562 251288
rect 128266 251232 128322 251288
rect 129646 251232 129702 251288
rect 131026 251232 131082 251288
rect 35162 227740 35164 227760
rect 35164 227740 35216 227760
rect 35216 227740 35218 227760
rect 35162 227704 35218 227740
rect 46754 227704 46810 227760
rect 47582 227704 47638 227760
rect 136362 251640 136418 251696
rect 135166 251232 135222 251288
rect 143354 252456 143410 252512
rect 148322 252456 148378 252512
rect 151082 252456 151138 252512
rect 138294 252320 138350 252376
rect 137926 251232 137982 251288
rect 142066 251912 142122 251968
rect 139214 251232 139270 251288
rect 140686 251232 140742 251288
rect 143446 252320 143502 252376
rect 166998 252592 167054 252648
rect 168470 511808 168526 511864
rect 168378 402872 168434 402928
rect 168378 401648 168434 401704
rect 168930 599936 168986 599992
rect 168746 598032 168802 598088
rect 168654 511944 168710 512000
rect 168654 510720 168710 510776
rect 168562 506096 168618 506152
rect 168562 456184 168618 456240
rect 168562 455504 168618 455560
rect 168470 399744 168526 399800
rect 169114 625912 169170 625968
rect 169206 623736 169262 623792
rect 169298 622784 169354 622840
rect 169482 621016 169538 621072
rect 169390 619928 169446 619984
rect 169022 514936 169078 514992
rect 169114 513848 169170 513904
rect 169298 511944 169354 512000
rect 169206 511808 169262 511864
rect 169666 598304 169722 598360
rect 169574 513848 169630 513904
rect 169482 508952 169538 509008
rect 169022 507864 169078 507920
rect 168930 487872 168986 487928
rect 168930 487192 168986 487248
rect 168838 486104 168894 486160
rect 168746 455776 168802 455832
rect 169114 506096 169170 506152
rect 168838 448568 168894 448624
rect 168746 399744 168802 399800
rect 168654 398792 168710 398848
rect 168654 397024 168710 397080
rect 168378 375264 168434 375320
rect 168378 374312 168434 374368
rect 167090 252048 167146 252104
rect 168562 374040 168618 374096
rect 168378 262248 168434 262304
rect 167642 245656 167698 245712
rect 122746 141752 122802 141808
rect 133142 141752 133198 141808
rect 108486 141616 108542 141672
rect 112166 141616 112222 141672
rect 109590 140664 109646 140720
rect 113270 140664 113326 140720
rect 116766 140664 116822 140720
rect 118974 140664 119030 140720
rect 43074 140120 43130 140176
rect 63222 140120 63278 140176
rect 65798 140120 65854 140176
rect 43442 139304 43498 139360
rect 60646 139304 60702 139360
rect 115478 140120 115534 140176
rect 115846 140120 115902 140176
rect 107382 139304 107438 139360
rect 110878 139304 110934 139360
rect 114374 139304 114430 139360
rect 68926 138624 68982 138680
rect 71042 138080 71098 138136
rect 74446 138080 74502 138136
rect 75826 138080 75882 138136
rect 78586 138080 78642 138136
rect 81346 138080 81402 138136
rect 84106 138080 84162 138136
rect 86866 138080 86922 138136
rect 88246 138080 88302 138136
rect 91006 138080 91062 138136
rect 93766 138080 93822 138136
rect 96526 138080 96582 138136
rect 99286 138080 99342 138136
rect 100666 138080 100722 138136
rect 103426 138080 103482 138136
rect 106186 138080 106242 138136
rect 108946 138080 109002 138136
rect 111706 138080 111762 138136
rect 113086 138080 113142 138136
rect 35806 117136 35862 117192
rect 45834 117000 45890 117056
rect 46938 116728 46994 116784
rect 117870 139304 117926 139360
rect 120354 139340 120356 139360
rect 120356 139340 120408 139360
rect 120408 139340 120410 139360
rect 120354 139304 120410 139340
rect 121366 139304 121422 139360
rect 122654 139304 122710 139360
rect 123758 141616 123814 141672
rect 128542 141616 128598 141672
rect 134246 141616 134302 141672
rect 136546 141616 136602 141672
rect 140042 141616 140098 141672
rect 142342 141616 142398 141672
rect 125966 140664 126022 140720
rect 132038 140664 132094 140720
rect 135350 140684 135406 140720
rect 135350 140664 135352 140684
rect 135352 140664 135404 140684
rect 135404 140664 135406 140684
rect 137926 140700 137928 140720
rect 137928 140700 137980 140720
rect 137980 140700 137982 140720
rect 137926 140664 137982 140700
rect 139030 140664 139086 140720
rect 141238 140664 141294 140720
rect 143446 140664 143502 140720
rect 149518 140664 149574 140720
rect 129646 140120 129702 140176
rect 125230 139304 125286 139360
rect 127714 139304 127770 139360
rect 122746 138624 122802 138680
rect 124126 138624 124182 138680
rect 130750 139304 130806 139360
rect 148414 139304 148470 139360
rect 151082 139304 151138 139360
rect 136454 139032 136510 139088
rect 118422 138080 118478 138136
rect 121366 138080 121422 138136
rect 125414 138080 125470 138136
rect 128266 138080 128322 138136
rect 131026 138080 131082 138136
rect 133786 138080 133842 138136
rect 139306 138080 139362 138136
rect 28906 109248 28962 109304
rect 128358 29824 128414 29880
rect 75550 29552 75606 29608
rect 88062 29552 88118 29608
rect 90730 29552 90786 29608
rect 122746 29552 122802 29608
rect 60646 28872 60702 28928
rect 68190 28872 68246 28928
rect 78126 28872 78182 28928
rect 80702 28872 80758 28928
rect 83094 28872 83150 28928
rect 103150 28872 103206 28928
rect 63222 28192 63278 28248
rect 112166 28192 112222 28248
rect 115662 28192 115718 28248
rect 42798 27548 42800 27568
rect 42800 27548 42852 27568
rect 42852 27548 42854 27568
rect 42798 27512 42854 27548
rect 43626 27532 43682 27568
rect 43626 27512 43628 27532
rect 43628 27512 43680 27532
rect 43680 27512 43682 27532
rect 64878 27512 64934 27568
rect 71594 27512 71650 27568
rect 73986 27512 74042 27568
rect 86590 27512 86646 27568
rect 92754 27512 92810 27568
rect 95238 27512 95294 27568
rect 98274 27512 98330 27568
rect 100206 27512 100262 27568
rect 105542 27512 105598 27568
rect 106278 27512 106334 27568
rect 108026 27512 108082 27568
rect 108762 27512 108818 27568
rect 110326 27512 110382 27568
rect 110970 27512 111026 27568
rect 3422 19352 3478 19408
rect 111522 27376 111578 27432
rect 112902 27512 112958 27568
rect 122746 27648 122802 27704
rect 117134 27512 117190 27568
rect 118238 27512 118294 27568
rect 118422 27512 118478 27568
rect 120078 27376 120134 27432
rect 120814 27512 120870 27568
rect 120630 27240 120686 27296
rect 130566 29552 130622 29608
rect 128542 28872 128598 28928
rect 134246 28908 134248 28928
rect 134248 28908 134300 28928
rect 134300 28908 134302 28928
rect 134246 28872 134302 28908
rect 129646 28192 129702 28248
rect 132038 28192 132094 28248
rect 124126 27512 124182 27568
rect 126334 27512 126390 27568
rect 128174 27512 128230 27568
rect 123758 27124 123814 27160
rect 123758 27104 123760 27124
rect 123760 27104 123812 27124
rect 123812 27104 123814 27124
rect 132774 27548 132776 27568
rect 132776 27548 132828 27568
rect 132828 27548 132830 27568
rect 132774 27512 132830 27548
rect 135350 27512 135406 27568
rect 138938 29552 138994 29608
rect 135902 28872 135958 28928
rect 138294 28872 138350 28928
rect 137190 27512 137246 27568
rect 140134 27512 140190 27568
rect 141238 27512 141294 27568
rect 149058 28328 149114 28384
rect 143446 28192 143502 28248
rect 143354 28056 143410 28112
rect 147678 27512 147734 27568
rect 143446 26560 143502 26616
rect 137190 24792 137246 24848
rect 150070 27512 150126 27568
rect 150622 27548 150624 27568
rect 150624 27548 150676 27568
rect 150676 27548 150678 27568
rect 150622 27512 150678 27548
rect 168930 401648 168986 401704
rect 168838 395936 168894 395992
rect 168746 288360 168802 288416
rect 168746 285640 168802 285696
rect 168654 284960 168710 285016
rect 168562 261976 168618 262032
rect 168194 238584 168250 238640
rect 168562 228928 168618 228984
rect 169206 455504 169262 455560
rect 169022 395936 169078 395992
rect 168930 290808 168986 290864
rect 168838 283872 168894 283928
rect 169022 288360 169078 288416
rect 169022 287680 169078 287736
rect 168930 178880 168986 178936
rect 169390 487192 169446 487248
rect 169206 379480 169262 379536
rect 173162 587424 173218 587480
rect 169666 486240 169722 486296
rect 169850 454688 169906 454744
rect 169850 454008 169906 454064
rect 170310 451188 170312 451208
rect 170312 451188 170364 451208
rect 170364 451188 170366 451208
rect 170310 451152 170366 451188
rect 169574 401920 169630 401976
rect 169482 397024 169538 397080
rect 169482 394168 169538 394224
rect 169390 375944 169446 376000
rect 169298 375264 169354 375320
rect 169114 282104 169170 282160
rect 168930 175752 168986 175808
rect 168838 174800 168894 174856
rect 168746 173032 168802 173088
rect 168930 171944 168986 172000
rect 168378 153040 168434 153096
rect 168378 151952 168434 152008
rect 169666 398792 169722 398848
rect 169574 289856 169630 289912
rect 170126 423580 170128 423600
rect 170128 423580 170180 423600
rect 170180 423580 170182 423600
rect 170126 423544 170182 423580
rect 169666 286728 169722 286784
rect 169666 285640 169722 285696
rect 169206 264016 169262 264072
rect 169850 251368 169906 251424
rect 170586 454008 170642 454064
rect 171138 584568 171194 584624
rect 170770 361664 170826 361720
rect 169298 177928 169354 177984
rect 168562 150356 168564 150376
rect 168564 150356 168616 150376
rect 168616 150356 168618 150376
rect 168562 150320 168618 150356
rect 168470 150048 168526 150104
rect 168378 39888 168434 39944
rect 168746 150048 168802 150104
rect 169114 170176 169170 170232
rect 169114 153040 169170 153096
rect 168838 66952 168894 67008
rect 168838 66000 168894 66056
rect 168838 63824 168894 63880
rect 168930 61104 168986 61160
rect 168838 60016 168894 60072
rect 168838 58248 168894 58304
rect 168562 38392 168618 38448
rect 168470 38120 168526 38176
rect 169390 62872 169446 62928
rect 170586 28736 170642 28792
rect 170494 27240 170550 27296
rect 172150 587152 172206 587208
rect 170678 26832 170734 26888
rect 170402 26152 170458 26208
rect 172426 475224 172482 475280
rect 172794 427624 172850 427680
rect 173070 455640 173126 455696
rect 173990 584296 174046 584352
rect 173714 427624 173770 427680
rect 175278 474988 175280 475008
rect 175280 474988 175332 475008
rect 175332 474988 175334 475008
rect 175278 474952 175334 474988
rect 176658 475088 176714 475144
rect 174634 26968 174690 27024
rect 178866 453192 178922 453248
rect 177302 27376 177358 27432
rect 177486 26696 177542 26752
rect 178682 28328 178738 28384
rect 181442 444896 181498 444952
rect 180154 352552 180210 352608
rect 178774 27104 178830 27160
rect 181534 28192 181590 28248
rect 187698 474816 187754 474872
rect 246302 659676 246304 659696
rect 246304 659676 246356 659696
rect 246356 659676 246358 659696
rect 246302 659640 246358 659676
rect 237286 654472 237342 654528
rect 237194 591640 237250 591696
rect 188342 28872 188398 28928
rect 192482 342896 192538 342952
rect 192942 445032 192998 445088
rect 193126 445304 193182 445360
rect 194322 445168 194378 445224
rect 196162 453192 196218 453248
rect 193954 24792 194010 24848
rect 196714 421368 196770 421424
rect 198370 574640 198426 574696
rect 196898 417152 196954 417208
rect 196806 402328 196862 402384
rect 197358 533160 197414 533216
rect 198278 473320 198334 473376
rect 198186 471688 198242 471744
rect 198094 470328 198150 470384
rect 198002 468832 198058 468888
rect 197818 467608 197874 467664
rect 197818 421640 197874 421696
rect 197358 419056 197414 419112
rect 197358 416608 197414 416664
rect 197358 414976 197414 415032
rect 197358 413480 197414 413536
rect 197358 412256 197414 412312
rect 197358 411032 197414 411088
rect 197358 409828 197414 409864
rect 197358 409808 197360 409828
rect 197360 409808 197412 409828
rect 197412 409808 197414 409828
rect 197450 408584 197506 408640
rect 197358 407904 197414 407960
rect 197726 406000 197782 406056
rect 197358 404776 197414 404832
rect 197358 403552 197414 403608
rect 197358 401104 197414 401160
rect 197358 399880 197414 399936
rect 197358 398656 197414 398712
rect 197450 397432 197506 397488
rect 197358 396072 197414 396128
rect 197358 394848 197414 394904
rect 197358 393624 197414 393680
rect 197358 392400 197414 392456
rect 197358 391176 197414 391232
rect 197358 389952 197414 390008
rect 197358 388728 197414 388784
rect 197358 387504 197414 387560
rect 197358 386300 197414 386336
rect 197358 386280 197360 386300
rect 197360 386280 197412 386300
rect 197412 386280 197414 386300
rect 197726 385056 197782 385112
rect 197358 384376 197414 384432
rect 197358 383152 197414 383208
rect 197358 381248 197414 381304
rect 197358 380024 197414 380080
rect 197358 378800 197414 378856
rect 197358 377576 197414 377632
rect 197358 376352 197414 376408
rect 197358 375128 197414 375184
rect 197358 373940 197360 373960
rect 197360 373940 197412 373960
rect 197412 373940 197414 373960
rect 197358 373904 197414 373940
rect 197358 372564 197414 372600
rect 197358 372544 197360 372564
rect 197360 372544 197412 372564
rect 197412 372544 197414 372564
rect 197450 371320 197506 371376
rect 197358 370096 197414 370152
rect 197358 368872 197414 368928
rect 197358 368328 197414 368384
rect 197358 367004 197360 367024
rect 197360 367004 197412 367024
rect 197412 367004 197414 367024
rect 197358 366968 197414 367004
rect 197358 365200 197414 365256
rect 197358 363976 197414 364032
rect 197358 362752 197414 362808
rect 197358 361392 197414 361448
rect 197450 360168 197506 360224
rect 197358 359624 197414 359680
rect 197358 357720 197414 357776
rect 197358 356496 197414 356552
rect 197358 355272 197414 355328
rect 197358 354048 197414 354104
rect 197358 352824 197414 352880
rect 197358 351600 197414 351656
rect 197358 350376 197414 350432
rect 197450 349036 197506 349072
rect 197450 349016 197452 349036
rect 197452 349016 197504 349036
rect 197504 349016 197506 349036
rect 197358 347792 197414 347848
rect 197358 346568 197414 346624
rect 197358 345344 197414 345400
rect 197358 344800 197414 344856
rect 197358 343440 197414 343496
rect 197358 341672 197414 341728
rect 197358 340448 197414 340504
rect 197358 339224 197414 339280
rect 197358 337864 197414 337920
rect 197450 336660 197506 336696
rect 197450 336640 197452 336660
rect 197452 336640 197504 336660
rect 197504 336640 197506 336660
rect 197358 336096 197414 336152
rect 197358 334192 197414 334248
rect 197358 332968 197414 333024
rect 197358 331744 197414 331800
rect 197358 330520 197414 330576
rect 197358 329296 197414 329352
rect 197358 328380 197360 328400
rect 197360 328380 197412 328400
rect 197412 328380 197414 328400
rect 197358 328344 197414 328380
rect 197358 327020 197360 327040
rect 197360 327020 197412 327040
rect 197412 327020 197414 327040
rect 197358 326984 197414 327020
rect 197358 325488 197414 325544
rect 197358 324264 197414 324320
rect 197450 323040 197506 323096
rect 197358 321816 197414 321872
rect 197358 320592 197414 320648
rect 197358 319368 197414 319424
rect 197358 318144 197414 318200
rect 197358 316920 197414 316976
rect 197358 315696 197414 315752
rect 197358 314336 197414 314392
rect 197358 313148 197360 313168
rect 197360 313148 197412 313168
rect 197412 313148 197414 313168
rect 197358 313112 197414 313148
rect 197450 312568 197506 312624
rect 197358 311344 197414 311400
rect 197358 309440 197414 309496
rect 197358 308216 197414 308272
rect 197726 306992 197782 307048
rect 197358 305768 197414 305824
rect 197358 304544 197414 304600
rect 197358 303456 197414 303512
rect 197358 301960 197414 302016
rect 197358 300772 197360 300792
rect 197360 300772 197412 300792
rect 197412 300772 197414 300792
rect 197358 300736 197414 300772
rect 197358 299532 197414 299568
rect 197358 299512 197360 299532
rect 197360 299512 197412 299532
rect 197412 299512 197414 299532
rect 197358 298288 197414 298344
rect 197358 297064 197414 297120
rect 197358 295432 197414 295488
rect 197358 294344 197414 294400
rect 197358 293392 197414 293448
rect 197358 292032 197414 292088
rect 197358 290808 197414 290864
rect 197358 289584 197414 289640
rect 197450 288360 197506 288416
rect 197358 287136 197414 287192
rect 197358 285912 197414 285968
rect 197358 284688 197414 284744
rect 197358 283464 197414 283520
rect 197358 282240 197414 282296
rect 197358 281016 197414 281072
rect 197358 279112 197414 279168
rect 197358 278432 197414 278488
rect 197450 277208 197506 277264
rect 197358 275984 197414 276040
rect 197358 274760 197414 274816
rect 197358 273536 197414 273592
rect 197358 272312 197414 272368
rect 197358 270564 197414 270600
rect 197358 270544 197360 270564
rect 197360 270544 197412 270564
rect 197412 270544 197414 270564
rect 197818 269864 197874 269920
rect 197358 268504 197414 268560
rect 197358 267280 197414 267336
rect 197358 266056 197414 266112
rect 197450 264832 197506 264888
rect 197358 263628 197414 263664
rect 197358 263608 197360 263628
rect 197360 263608 197412 263628
rect 197412 263608 197414 263628
rect 197358 262384 197414 262440
rect 197358 261160 197414 261216
rect 197358 258712 197414 258768
rect 197542 254768 197598 254824
rect 197450 252476 197506 252512
rect 197450 252456 197452 252476
rect 197452 252456 197504 252476
rect 197504 252456 197506 252476
rect 198002 448432 198058 448488
rect 197910 257352 197966 257408
rect 198094 448296 198150 448352
rect 198002 256128 198058 256184
rect 198186 448160 198242 448216
rect 198094 254768 198150 254824
rect 198278 448024 198334 448080
rect 198186 253816 198242 253872
rect 336738 603744 336794 603800
rect 238666 594632 238722 594688
rect 238574 593000 238630 593056
rect 253110 576136 253166 576192
rect 292486 576136 292542 576192
rect 284206 575320 284262 575376
rect 285310 575320 285366 575376
rect 286598 575320 286654 575376
rect 287886 575320 287942 575376
rect 280158 575048 280214 575104
rect 280250 574932 280306 574968
rect 280250 574912 280252 574932
rect 280252 574912 280304 574932
rect 280304 574912 280306 574932
rect 281538 574912 281594 574968
rect 253754 574368 253810 574424
rect 273258 574368 273314 574424
rect 276018 574368 276074 574424
rect 254582 574232 254638 574288
rect 269210 574232 269266 574288
rect 253846 574096 253902 574152
rect 269118 574096 269174 574152
rect 270498 574096 270554 574152
rect 271878 574096 271934 574152
rect 274638 574232 274694 574288
rect 284390 575184 284446 575240
rect 284298 574796 284354 574832
rect 284298 574776 284300 574796
rect 284300 574776 284352 574796
rect 284352 574776 284354 574796
rect 278778 574232 278834 574288
rect 285678 574232 285734 574288
rect 277674 574096 277730 574152
rect 278686 574096 278742 574152
rect 237286 542952 237342 543008
rect 287518 574912 287574 574968
rect 289818 575184 289874 575240
rect 291198 575048 291254 575104
rect 291106 574912 291162 574968
rect 288438 574776 288494 574832
rect 291014 574776 291070 574832
rect 289726 574504 289782 574560
rect 280066 574096 280122 574152
rect 281446 574096 281502 574152
rect 282826 574096 282882 574152
rect 284206 574096 284262 574152
rect 217598 539688 217654 539744
rect 218058 539552 218114 539608
rect 205730 539144 205786 539200
rect 297914 575320 297970 575376
rect 300674 575320 300730 575376
rect 301870 575320 301926 575376
rect 302882 575320 302938 575376
rect 304630 575320 304686 575376
rect 305550 575320 305606 575376
rect 306286 575320 306342 575376
rect 307574 575320 307630 575376
rect 320454 575320 320510 575376
rect 330206 575320 330262 575376
rect 330482 575320 330538 575376
rect 293958 575204 294014 575240
rect 293958 575184 293960 575204
rect 293960 575184 294012 575204
rect 294012 575184 294014 575204
rect 293958 575068 294014 575104
rect 293958 575048 293960 575068
rect 293960 575048 294012 575068
rect 294012 575048 294014 575068
rect 292578 574776 292634 574832
rect 296534 574504 296590 574560
rect 293774 574368 293830 574424
rect 294694 574368 294750 574424
rect 295338 574096 295394 574152
rect 298926 574504 298982 574560
rect 299202 574504 299258 574560
rect 299478 574504 299534 574560
rect 298190 574232 298246 574288
rect 298098 574096 298154 574152
rect 303618 574232 303674 574288
rect 300858 574096 300914 574152
rect 302238 574096 302294 574152
rect 304998 574096 305054 574152
rect 306470 574116 306526 574152
rect 306470 574096 306472 574116
rect 306472 574096 306524 574116
rect 306524 574096 306526 574116
rect 318706 574096 318762 574152
rect 288898 453736 288954 453792
rect 213182 453600 213238 453656
rect 284298 453600 284354 453656
rect 286782 453600 286838 453656
rect 198278 252456 198334 252512
rect 197542 251504 197598 251560
rect 197358 251232 197414 251288
rect 197266 248784 197322 248840
rect 197358 246336 197414 246392
rect 197358 244976 197414 245032
rect 197358 243752 197414 243808
rect 197358 242528 197414 242584
rect 197542 241304 197598 241360
rect 197450 239536 197506 239592
rect 197358 238892 197360 238912
rect 197360 238892 197412 238912
rect 197412 238892 197414 238912
rect 197358 238856 197414 238892
rect 197358 236408 197414 236464
rect 197726 235184 197782 235240
rect 197358 233824 197414 233880
rect 197358 232600 197414 232656
rect 197818 232600 197874 232656
rect 197358 231648 197414 231704
rect 197542 230152 197598 230208
rect 197358 224032 197414 224088
rect 197358 220224 197414 220280
rect 197358 217776 197414 217832
rect 197358 216552 197414 216608
rect 197358 214104 197414 214160
rect 197358 212880 197414 212936
rect 197358 210296 197414 210352
rect 197358 208292 197360 208312
rect 197360 208292 197412 208312
rect 197412 208292 197414 208312
rect 197358 208256 197414 208292
rect 197358 206624 197414 206680
rect 197358 205400 197414 205456
rect 197358 204196 197414 204232
rect 197358 204176 197360 204196
rect 197360 204176 197412 204196
rect 197412 204176 197414 204196
rect 197358 201728 197414 201784
rect 197358 200504 197414 200560
rect 197358 199144 197414 199200
rect 197358 197956 197360 197976
rect 197360 197956 197412 197976
rect 197412 197956 197414 197976
rect 197358 197920 197414 197956
rect 197358 196696 197414 196752
rect 197358 195472 197414 195528
rect 197358 194248 197414 194304
rect 197358 193024 197414 193080
rect 197358 190576 197414 190632
rect 197358 189352 197414 189408
rect 197358 188128 197414 188184
rect 197358 186768 197414 186824
rect 197358 185580 197360 185600
rect 197360 185580 197412 185600
rect 197412 185580 197414 185600
rect 197358 185544 197414 185580
rect 197358 184204 197414 184240
rect 197358 184184 197360 184204
rect 197360 184184 197412 184204
rect 197412 184184 197414 184204
rect 197358 182844 197414 182880
rect 197358 182824 197360 182844
rect 197360 182824 197412 182844
rect 197412 182824 197414 182844
rect 197358 181872 197414 181928
rect 197358 180648 197414 180704
rect 197358 179460 197360 179480
rect 197360 179460 197412 179480
rect 197412 179460 197414 179480
rect 197358 179424 197414 179460
rect 197358 176976 197414 177032
rect 197358 175652 197360 175672
rect 197360 175652 197412 175672
rect 197412 175652 197414 175672
rect 197358 175616 197414 175652
rect 197358 174392 197414 174448
rect 197358 173204 197360 173224
rect 197360 173204 197412 173224
rect 197412 173204 197414 173224
rect 197358 173168 197414 173204
rect 197358 171944 197414 172000
rect 197358 170720 197414 170776
rect 197358 169496 197414 169552
rect 197358 167728 197414 167784
rect 197358 165824 197414 165880
rect 197358 164464 197414 164520
rect 197358 163240 197414 163296
rect 197358 162016 197414 162072
rect 197358 160792 197414 160848
rect 197358 159432 197414 159488
rect 197358 158364 197414 158400
rect 197358 158344 197360 158364
rect 197360 158344 197412 158364
rect 197412 158344 197414 158364
rect 197358 157120 197414 157176
rect 197358 155896 197414 155952
rect 197358 153448 197414 153504
rect 197358 152768 197414 152824
rect 197358 150476 197414 150512
rect 197358 150456 197360 150476
rect 197360 150456 197412 150476
rect 197412 150456 197414 150476
rect 197358 149640 197414 149696
rect 197358 147192 197414 147248
rect 197358 145968 197414 146024
rect 197358 144764 197414 144800
rect 197358 144744 197360 144764
rect 197360 144744 197412 144764
rect 197412 144744 197414 144764
rect 197358 143556 197360 143576
rect 197360 143556 197412 143576
rect 197412 143556 197414 143576
rect 197358 143520 197414 143556
rect 197358 142296 197414 142352
rect 197542 226480 197598 226536
rect 197634 211656 197690 211712
rect 198370 228928 198426 228984
rect 198554 226480 198610 226536
rect 198462 225256 198518 225312
rect 198646 224032 198702 224088
rect 199290 425720 199346 425776
rect 199382 259528 199438 259584
rect 200118 421504 200174 421560
rect 231766 452512 231822 452568
rect 234526 452512 234582 452568
rect 235906 452512 235962 452568
rect 238666 452512 238722 452568
rect 241426 452512 241482 452568
rect 243174 452512 243230 452568
rect 245566 452512 245622 452568
rect 253846 452512 253902 452568
rect 255686 452512 255742 452568
rect 260746 452512 260802 452568
rect 263506 452512 263562 452568
rect 265622 452512 265678 452568
rect 269026 452512 269082 452568
rect 271786 452512 271842 452568
rect 273166 452512 273222 452568
rect 275834 452512 275890 452568
rect 213366 452376 213422 452432
rect 213182 451424 213238 451480
rect 204534 447888 204590 447944
rect 206834 445304 206890 445360
rect 208030 445168 208086 445224
rect 209318 445032 209374 445088
rect 240782 447752 240838 447808
rect 248234 451288 248290 451344
rect 251086 451288 251142 451344
rect 249522 447888 249578 447944
rect 248326 439456 248382 439512
rect 250810 447616 250866 447672
rect 259366 451288 259422 451344
rect 278686 452512 278742 452568
rect 280158 452512 280214 452568
rect 294786 453736 294842 453792
rect 282090 452512 282146 452568
rect 284206 452512 284262 452568
rect 285586 452512 285642 452568
rect 288346 452512 288402 452568
rect 283194 452240 283250 452296
rect 281446 452104 281502 452160
rect 290186 453600 290242 453656
rect 291198 453600 291254 453656
rect 293682 453600 293738 453656
rect 297086 453600 297142 453656
rect 298466 453600 298522 453656
rect 299570 453600 299626 453656
rect 311070 453600 311126 453656
rect 312358 453600 312414 453656
rect 297086 452648 297142 452704
rect 291106 452512 291162 452568
rect 292578 452512 292634 452568
rect 293038 452512 293094 452568
rect 296626 452512 296682 452568
rect 294786 451968 294842 452024
rect 293590 451832 293646 451888
rect 297362 452104 297418 452160
rect 299386 452512 299442 452568
rect 300766 452512 300822 452568
rect 300122 452240 300178 452296
rect 301962 452512 302018 452568
rect 303066 452512 303122 452568
rect 304170 452512 304226 452568
rect 305274 452548 305276 452568
rect 305276 452548 305328 452568
rect 305328 452548 305330 452568
rect 305274 452512 305330 452548
rect 306378 452512 306434 452568
rect 307850 452512 307906 452568
rect 308954 452512 309010 452568
rect 309874 452512 309930 452568
rect 303526 452240 303582 452296
rect 306286 452240 306342 452296
rect 307390 445032 307446 445088
rect 309046 451288 309102 451344
rect 313370 452532 313426 452568
rect 313370 452512 313372 452532
rect 313372 452512 313424 452532
rect 313424 452512 313426 452532
rect 314658 452512 314714 452568
rect 320178 452512 320234 452568
rect 319442 452240 319498 452296
rect 336922 585248 336978 585304
rect 340142 659640 340198 659696
rect 339406 612176 339462 612232
rect 339406 610952 339462 611008
rect 338302 609184 338358 609240
rect 338118 608096 338174 608152
rect 337382 583616 337438 583672
rect 337014 574232 337070 574288
rect 337106 574096 337162 574152
rect 338026 575320 338082 575376
rect 337566 575184 337622 575240
rect 338394 606464 338450 606520
rect 339406 605512 339462 605568
rect 339222 603764 339278 603800
rect 339222 603744 339224 603764
rect 339224 603744 339276 603764
rect 339276 603744 339278 603764
rect 339222 585248 339278 585304
rect 339406 583616 339462 583672
rect 338486 575048 338542 575104
rect 339406 490864 339462 490920
rect 339314 489912 339370 489968
rect 338854 486784 338910 486840
rect 339406 485016 339462 485072
rect 338854 482160 338910 482216
rect 339406 463936 339462 463992
rect 339130 462304 339186 462360
rect 339038 461488 339094 461544
rect 340050 487736 340106 487792
rect 340050 483928 340106 483984
rect 341246 574912 341302 574968
rect 341062 574776 341118 574832
rect 341154 574640 341210 574696
rect 341614 543088 341670 543144
rect 341522 450880 341578 450936
rect 337382 421776 337438 421832
rect 338854 421776 338910 421832
rect 340050 421776 340106 421832
rect 341614 428032 341670 428088
rect 390098 421640 390154 421696
rect 391386 419600 391442 419656
rect 407118 612176 407174 612232
rect 407118 610952 407174 611008
rect 407118 609184 407174 609240
rect 407118 608096 407174 608152
rect 407118 606464 407174 606520
rect 407118 605512 407174 605568
rect 407118 603764 407174 603800
rect 407118 603744 407120 603764
rect 407120 603744 407172 603764
rect 407172 603744 407174 603764
rect 407118 585248 407174 585304
rect 407118 583616 407174 583672
rect 405186 572192 405242 572248
rect 405554 572328 405610 572384
rect 405370 572056 405426 572112
rect 405370 452104 405426 452160
rect 405554 451968 405610 452024
rect 407118 490864 407174 490920
rect 407210 489912 407266 489968
rect 407118 487736 407174 487792
rect 407118 486784 407174 486840
rect 407118 485016 407174 485072
rect 407118 483928 407174 483984
rect 407118 482160 407174 482216
rect 407118 463936 407174 463992
rect 407118 462304 407174 462360
rect 407118 462032 407174 462088
rect 406474 445032 406530 445088
rect 408222 574776 408278 574832
rect 407946 571920 408002 571976
rect 408222 451832 408278 451888
rect 396354 421504 396410 421560
rect 395066 421368 395122 421424
rect 409142 575048 409198 575104
rect 409326 574912 409382 574968
rect 488906 659640 488962 659696
rect 499854 659676 499856 659696
rect 499856 659676 499908 659696
rect 499908 659676 499910 659696
rect 499854 659640 499910 659676
rect 507858 654472 507914 654528
rect 506570 594632 506626 594688
rect 506478 593000 506534 593056
rect 492678 577768 492734 577824
rect 441802 576952 441858 577008
rect 462870 576952 462926 577008
rect 415398 575320 415454 575376
rect 425058 575320 425114 575376
rect 426438 575184 426494 575240
rect 437478 575184 437534 575240
rect 438858 574796 438914 574832
rect 438858 574776 438860 574796
rect 438860 574776 438912 574796
rect 438912 574776 438914 574796
rect 433338 574368 433394 574424
rect 436098 574232 436154 574288
rect 440330 574232 440386 574288
rect 434718 574096 434774 574152
rect 433338 572328 433394 572384
rect 434718 572192 434774 572248
rect 436190 574096 436246 574152
rect 437570 574096 437626 574152
rect 438950 574096 439006 574152
rect 440238 574096 440294 574152
rect 436098 572056 436154 572112
rect 441618 574096 441674 574152
rect 455510 576136 455566 576192
rect 459282 576136 459338 576192
rect 448518 575048 448574 575104
rect 444378 574776 444434 574832
rect 451278 574660 451334 574696
rect 451278 574640 451280 574660
rect 451280 574640 451332 574660
rect 451332 574640 451334 574660
rect 451278 574524 451334 574560
rect 451278 574504 451280 574524
rect 451280 574504 451332 574524
rect 451332 574504 451334 574524
rect 455418 574504 455474 574560
rect 443090 574232 443146 574288
rect 444562 574232 444618 574288
rect 445850 574232 445906 574288
rect 447230 574232 447286 574288
rect 449990 574232 450046 574288
rect 452750 574232 452806 574288
rect 454130 574232 454186 574288
rect 442998 574096 443054 574152
rect 444470 574096 444526 574152
rect 445758 574096 445814 574152
rect 447138 574096 447194 574152
rect 448610 574096 448666 574152
rect 449898 574096 449954 574152
rect 451278 574096 451334 574152
rect 452658 574096 452714 574152
rect 454038 574096 454094 574152
rect 458178 574388 458234 574424
rect 458178 574368 458180 574388
rect 458180 574368 458232 574388
rect 458232 574368 458234 574388
rect 456890 574232 456946 574288
rect 455602 574096 455658 574152
rect 456798 574096 456854 574152
rect 458362 574096 458418 574152
rect 459558 574368 459614 574424
rect 468482 576136 468538 576192
rect 466458 575184 466514 575240
rect 463790 574504 463846 574560
rect 461122 574232 461178 574288
rect 459650 574096 459706 574152
rect 461306 574096 461362 574152
rect 462410 574096 462466 574152
rect 463698 574096 463754 574152
rect 465078 574368 465134 574424
rect 464342 574232 464398 574288
rect 466458 574096 466514 574152
rect 466642 574096 466698 574152
rect 467838 574096 467894 574152
rect 492954 576816 493010 576872
rect 470690 574232 470746 574288
rect 470598 574096 470654 574152
rect 471978 574096 472034 574152
rect 473358 574096 473414 574152
rect 474738 574096 474794 574152
rect 476118 574096 476174 574152
rect 492678 574368 492734 574424
rect 492770 574252 492826 574288
rect 492770 574232 492772 574252
rect 492772 574232 492824 574252
rect 492824 574232 492826 574252
rect 506570 576000 506626 576056
rect 507950 591640 508006 591696
rect 507858 542952 507914 543008
rect 527178 540268 527180 540288
rect 527180 540268 527232 540288
rect 527232 540268 527234 540288
rect 527178 540232 527234 540268
rect 528834 539688 528890 539744
rect 540794 538736 540850 538792
rect 443642 453600 443698 453656
rect 425426 452512 425482 452568
rect 426898 452512 426954 452568
rect 428462 452512 428518 452568
rect 432050 452512 432106 452568
rect 433706 452512 433762 452568
rect 434718 452512 434774 452568
rect 436282 452512 436338 452568
rect 401598 421232 401654 421288
rect 405186 421096 405242 421152
rect 411442 420960 411498 421016
rect 431866 444896 431922 444952
rect 433154 450744 433210 450800
rect 438674 452240 438730 452296
rect 437662 451560 437718 451616
rect 437570 451288 437626 451344
rect 438122 450608 438178 450664
rect 441618 452104 441674 452160
rect 442998 452104 443054 452160
rect 440238 451560 440294 451616
rect 438950 451288 439006 451344
rect 441526 451288 441582 451344
rect 450266 452512 450322 452568
rect 452842 452512 452898 452568
rect 466182 452532 466238 452568
rect 466182 452512 466184 452532
rect 466184 452512 466236 452532
rect 466236 452512 466238 452532
rect 445758 452104 445814 452160
rect 447046 452104 447102 452160
rect 448610 452104 448666 452160
rect 444470 451288 444526 451344
rect 445666 450472 445722 450528
rect 443182 438096 443238 438152
rect 441618 425584 441674 425640
rect 445850 451288 445906 451344
rect 447230 451288 447286 451344
rect 448518 451288 448574 451344
rect 451370 452104 451426 452160
rect 451186 451288 451242 451344
rect 452750 451288 452806 451344
rect 466550 452512 466606 452568
rect 454130 452240 454186 452296
rect 462318 452240 462374 452296
rect 453670 452104 453726 452160
rect 456706 452104 456762 452160
rect 459742 452104 459798 452160
rect 455510 451288 455566 451344
rect 453210 432520 453266 432576
rect 459466 451560 459522 451616
rect 456890 451288 456946 451344
rect 458270 451288 458326 451344
rect 461030 449248 461086 449304
rect 462226 449112 462282 449168
rect 462410 452104 462466 452160
rect 463606 452104 463662 452160
rect 465078 452104 465134 452160
rect 463790 451288 463846 451344
rect 467930 452512 467986 452568
rect 468022 452240 468078 452296
rect 468666 452512 468722 452568
rect 471886 452512 471942 452568
rect 473542 452532 473598 452568
rect 473542 452512 473544 452532
rect 473544 452512 473596 452532
rect 473596 452512 473598 452532
rect 476026 452512 476082 452568
rect 478418 452512 478474 452568
rect 481086 452532 481142 452568
rect 481086 452512 481088 452532
rect 481088 452512 481140 452532
rect 481140 452512 481142 452532
rect 483478 452512 483534 452568
rect 487066 452512 487122 452568
rect 488446 452512 488502 452568
rect 491022 452512 491078 452568
rect 493598 452532 493654 452568
rect 493598 452512 493600 452532
rect 493600 452512 493652 452532
rect 493652 452512 493654 452532
rect 495990 452512 496046 452568
rect 499486 452512 499542 452568
rect 501234 452512 501290 452568
rect 503534 452532 503590 452568
rect 503534 452512 503536 452532
rect 503536 452512 503588 452532
rect 503588 452512 503590 452532
rect 505926 452532 505982 452568
rect 505926 452512 505928 452532
rect 505928 452512 505980 452532
rect 505980 452512 505982 452532
rect 509146 452512 509202 452568
rect 511906 452512 511962 452568
rect 514666 452512 514722 452568
rect 516046 452512 516102 452568
rect 580446 697176 580502 697232
rect 549258 533160 549314 533216
rect 549350 473320 549406 473376
rect 549442 471688 549498 471744
rect 549534 470328 549590 470384
rect 549626 468832 549682 468888
rect 549718 467608 549774 467664
rect 549626 448432 549682 448488
rect 549534 448296 549590 448352
rect 549442 448160 549498 448216
rect 549350 448024 549406 448080
rect 549258 422864 549314 422920
rect 560206 415112 560262 415168
rect 560114 407088 560170 407144
rect 560022 399064 560078 399120
rect 560206 391176 560262 391232
rect 559194 383152 559250 383208
rect 560206 375128 560262 375184
rect 559194 367240 559250 367296
rect 559378 319368 559434 319424
rect 559286 303320 559342 303376
rect 559010 295296 559066 295352
rect 560206 359216 560262 359272
rect 559654 351192 559710 351248
rect 560206 343304 560262 343360
rect 560206 335300 560262 335336
rect 560206 335280 560208 335300
rect 560208 335280 560260 335300
rect 560260 335280 560262 335300
rect 559930 327256 559986 327312
rect 560206 311344 560262 311400
rect 560206 287408 560262 287464
rect 559930 279384 559986 279440
rect 559562 271360 559618 271416
rect 560206 263508 560208 263528
rect 560208 263508 560260 263528
rect 560260 263508 560262 263528
rect 560206 263472 560262 263508
rect 199474 258712 199530 258768
rect 560022 255448 560078 255504
rect 560206 247424 560262 247480
rect 560206 239572 560208 239592
rect 560208 239572 560260 239592
rect 560260 239572 560262 239592
rect 560206 239536 560262 239572
rect 199290 237632 199346 237688
rect 559194 231512 559250 231568
rect 199198 230152 199254 230208
rect 199106 227704 199162 227760
rect 560206 223524 560208 223544
rect 560208 223524 560260 223544
rect 560260 223524 560262 223544
rect 560206 223488 560262 223524
rect 199566 222876 199622 222932
rect 198922 221448 198978 221504
rect 198738 220224 198794 220280
rect 197910 219000 197966 219056
rect 559194 215600 559250 215656
rect 198094 215364 198096 215384
rect 198096 215364 198148 215384
rect 198148 215364 198150 215384
rect 198094 215328 198150 215364
rect 197726 209072 197782 209128
rect 197726 202952 197782 203008
rect 197726 192344 197782 192400
rect 197542 167592 197598 167648
rect 197542 154672 197598 154728
rect 197542 148416 197598 148472
rect 560206 207576 560262 207632
rect 559562 199552 559618 199608
rect 560206 191700 560208 191720
rect 560208 191700 560260 191720
rect 560260 191700 560262 191720
rect 560206 191664 560262 191700
rect 560022 183640 560078 183696
rect 197910 178236 197912 178256
rect 197912 178236 197964 178256
rect 197964 178236 197966 178256
rect 197910 178200 197966 178236
rect 560206 175616 560262 175672
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 578882 630808 578938 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 578974 537784 579030 537840
rect 578882 351872 578938 351928
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 579894 431568 579950 431624
rect 580630 484608 580686 484664
rect 580354 418240 580410 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579618 365064 579674 365120
rect 580078 325216 580134 325272
rect 580170 298696 580226 298752
rect 580446 312024 580502 312080
rect 579802 272176 579858 272232
rect 580170 258848 580226 258904
rect 580262 245520 580318 245576
rect 579802 232328 579858 232384
rect 579894 219000 579950 219056
rect 580262 205672 580318 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 559010 167592 559066 167648
rect 580170 165824 580226 165880
rect 559562 159704 559618 159760
rect 580262 152632 580318 152688
rect 559562 151680 559618 151736
rect 197266 140936 197322 140992
rect 197358 139712 197414 139768
rect 560022 143656 560078 143712
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 197450 138488 197506 138544
rect 197358 137264 197414 137320
rect 197358 136312 197414 136368
rect 559286 135768 559342 135824
rect 197358 134816 197414 134872
rect 197358 133592 197414 133648
rect 197358 132404 197360 132424
rect 197360 132404 197412 132424
rect 197412 132404 197414 132424
rect 197358 132368 197414 132404
rect 197450 131144 197506 131200
rect 197358 129784 197414 129840
rect 197358 129240 197414 129296
rect 197358 128016 197414 128072
rect 559562 127744 559618 127800
rect 197358 126112 197414 126168
rect 197358 124888 197414 124944
rect 197358 123664 197414 123720
rect 197358 122440 197414 122496
rect 197358 121216 197414 121272
rect 197358 120028 197360 120048
rect 197360 120028 197412 120048
rect 197412 120028 197414 120048
rect 197358 119992 197414 120028
rect 558918 119720 558974 119776
rect 197450 118768 197506 118824
rect 197358 117408 197414 117464
rect 197358 116184 197414 116240
rect 197358 114960 197414 115016
rect 197358 113736 197414 113792
rect 197358 113092 197360 113112
rect 197360 113092 197412 113112
rect 197412 113092 197414 113112
rect 197358 113056 197414 113092
rect 559194 111852 559250 111888
rect 559194 111832 559196 111852
rect 559196 111832 559248 111852
rect 559248 111832 559250 111852
rect 197358 111732 197360 111752
rect 197360 111732 197412 111752
rect 197412 111732 197414 111752
rect 197358 111696 197414 111732
rect 197358 110064 197414 110120
rect 197358 108876 197360 108896
rect 197360 108876 197412 108896
rect 197412 108876 197414 108896
rect 197358 108840 197414 108876
rect 197542 107616 197598 107672
rect 197450 106256 197506 106312
rect 197358 105032 197414 105088
rect 197358 103808 197414 103864
rect 197358 102584 197414 102640
rect 197358 101360 197414 101416
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 560206 103828 560262 103864
rect 560206 103808 560208 103828
rect 560208 103808 560260 103828
rect 560260 103808 560262 103828
rect 197358 100136 197414 100192
rect 197358 98912 197414 98968
rect 198002 97688 198058 97744
rect 197358 94560 197414 94616
rect 197358 92656 197414 92712
rect 197358 91432 197414 91488
rect 197358 90208 197414 90264
rect 197358 88984 197414 89040
rect 197358 87216 197414 87272
rect 197358 86536 197414 86592
rect 197358 85312 197414 85368
rect 197358 84088 197414 84144
rect 197450 82728 197506 82784
rect 197358 81504 197414 81560
rect 197358 80144 197414 80200
rect 197358 78784 197414 78840
rect 197358 77832 197414 77888
rect 197358 76608 197414 76664
rect 197358 75384 197414 75440
rect 197358 74160 197414 74216
rect 197358 72936 197414 72992
rect 197358 70388 197360 70408
rect 197360 70388 197412 70408
rect 197412 70388 197414 70408
rect 197358 70352 197414 70388
rect 197358 63824 197414 63880
rect 197910 63008 197966 63064
rect 197358 61784 197414 61840
rect 197542 60560 197598 60616
rect 198094 95920 198150 95976
rect 559746 95784 559802 95840
rect 198186 93880 198242 93936
rect 560206 87896 560262 87952
rect 560022 79872 560078 79928
rect 559194 71868 559250 71904
rect 559194 71848 559196 71868
rect 559196 71848 559248 71868
rect 559248 71848 559250 71868
rect 198278 71032 198334 71088
rect 198370 69128 198426 69184
rect 198462 67904 198518 67960
rect 198554 66680 198610 66736
rect 198646 65456 198702 65512
rect 560206 63960 560262 64016
rect 196806 26288 196862 26344
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 579618 19760 579674 19816
rect 580170 6568 580226 6624
rect 580354 33088 580410 33144
<< metal3 >>
rect 154113 700634 154179 700637
rect 196566 700634 196572 700636
rect 154113 700632 196572 700634
rect 154113 700576 154118 700632
rect 154174 700576 196572 700632
rect 154113 700574 196572 700576
rect 154113 700571 154179 700574
rect 196566 700572 196572 700574
rect 196636 700572 196642 700636
rect 89161 700498 89227 700501
rect 174670 700498 174676 700500
rect 89161 700496 174676 700498
rect 89161 700440 89166 700496
rect 89222 700440 174676 700496
rect 89161 700438 174676 700440
rect 89161 700435 89227 700438
rect 174670 700436 174676 700438
rect 174740 700436 174746 700500
rect 40493 700362 40559 700365
rect 174486 700362 174492 700364
rect 40493 700360 174492 700362
rect 40493 700304 40498 700360
rect 40554 700304 174492 700360
rect 40493 700302 174492 700304
rect 40493 700299 40559 700302
rect 174486 700300 174492 700302
rect 174556 700300 174562 700364
rect -960 697220 480 697460
rect 580441 697234 580507 697237
rect 583520 697234 584960 697324
rect 580441 697232 584960 697234
rect 580441 697176 580446 697232
rect 580502 697176 584960 697232
rect 580441 697174 584960 697176
rect 580441 697171 580507 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect 34513 674930 34579 674933
rect 35750 674930 35756 674932
rect 34513 674928 35756 674930
rect 34513 674872 34518 674928
rect 34574 674872 35756 674928
rect 34513 674870 35756 674872
rect 34513 674867 34579 674870
rect 35750 674868 35756 674870
rect 35820 674868 35826 674932
rect 46197 674930 46263 674933
rect 46790 674930 46796 674932
rect 46197 674928 46796 674930
rect 46197 674872 46202 674928
rect 46258 674872 46796 674928
rect 46197 674870 46796 674872
rect 46197 674867 46263 674870
rect 46790 674868 46796 674870
rect 46860 674868 46866 674932
rect 46933 674930 46999 674933
rect 48078 674930 48084 674932
rect 46933 674928 48084 674930
rect 46933 674872 46938 674928
rect 46994 674872 48084 674928
rect 46933 674870 48084 674872
rect 46933 674867 46999 674870
rect 48078 674868 48084 674870
rect 48148 674868 48154 674932
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 28165 669218 28231 669221
rect 28165 669216 30062 669218
rect 28165 669160 28170 669216
rect 28226 669160 30062 669216
rect 28165 669158 30062 669160
rect 28165 669155 28231 669158
rect 246297 659700 246363 659701
rect 340137 659700 340203 659701
rect 246246 659698 246252 659700
rect 246206 659638 246252 659698
rect 246316 659696 246363 659700
rect 246358 659640 246363 659696
rect 246246 659636 246252 659638
rect 246316 659636 246363 659640
rect 256550 659636 256556 659700
rect 256620 659698 256626 659700
rect 340086 659698 340092 659700
rect 256620 659638 340092 659698
rect 340156 659696 340203 659700
rect 340198 659640 340203 659696
rect 256620 659636 256626 659638
rect 340086 659636 340092 659638
rect 340156 659636 340203 659640
rect 246297 659635 246363 659636
rect 340137 659635 340203 659636
rect 488901 659700 488967 659701
rect 488901 659696 488948 659700
rect 489012 659698 489018 659700
rect 499849 659698 499915 659701
rect 499982 659698 499988 659700
rect 488901 659640 488906 659696
rect 488901 659636 488948 659640
rect 489012 659638 489058 659698
rect 499849 659696 499988 659698
rect 499849 659640 499854 659696
rect 499910 659640 499988 659696
rect 499849 659638 499988 659640
rect 489012 659636 489018 659638
rect 488901 659635 488967 659636
rect 499849 659635 499915 659638
rect 499982 659636 499988 659638
rect 500052 659636 500058 659700
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect 237281 654530 237347 654533
rect 507853 654530 507919 654533
rect 237281 654528 239506 654530
rect 237281 654472 237286 654528
rect 237342 654500 239506 654528
rect 506430 654528 507919 654530
rect 506430 654500 507858 654528
rect 237342 654472 240028 654500
rect 237281 654470 240028 654472
rect 237281 654467 237347 654470
rect 239446 654440 240028 654470
rect 505908 654472 507858 654500
rect 507914 654472 507919 654528
rect 505908 654470 507919 654472
rect 505908 654440 506490 654470
rect 507853 654467 507919 654470
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 578877 630866 578943 630869
rect 583520 630866 584960 630956
rect 578877 630864 584960 630866
rect 578877 630808 578882 630864
rect 578938 630808 584960 630864
rect 578877 630806 584960 630808
rect 578877 630803 578943 630806
rect 583520 630716 584960 630806
rect 166612 626922 167194 626924
rect 169017 626922 169083 626925
rect 166612 626920 169083 626922
rect 166612 626864 169022 626920
rect 169078 626864 169083 626920
rect 167134 626862 169083 626864
rect 169017 626859 169083 626862
rect 166612 625970 167194 625972
rect 169109 625970 169175 625973
rect 166612 625968 169175 625970
rect 166612 625912 169114 625968
rect 169170 625912 169175 625968
rect 167134 625910 169175 625912
rect 169109 625907 169175 625910
rect 166612 623794 167194 623796
rect 169201 623794 169267 623797
rect 166612 623792 169267 623794
rect 166612 623736 169206 623792
rect 169262 623736 169267 623792
rect 167134 623734 169267 623736
rect 169201 623731 169267 623734
rect 166612 622842 167194 622844
rect 169293 622842 169359 622845
rect 166612 622840 169359 622842
rect 166612 622784 169298 622840
rect 169354 622784 169359 622840
rect 167134 622782 169359 622784
rect 169293 622779 169359 622782
rect 166612 621074 167194 621076
rect 169477 621074 169543 621077
rect 166612 621072 169543 621074
rect 166612 621016 169482 621072
rect 169538 621016 169543 621072
rect 167134 621014 169543 621016
rect 169477 621011 169543 621014
rect 166612 619986 167194 619988
rect 169385 619986 169451 619989
rect 166612 619984 169451 619986
rect 166612 619928 169390 619984
rect 169446 619928 169451 619984
rect 167134 619926 169451 619928
rect 169385 619923 169451 619926
rect -960 619170 480 619260
rect 2957 619170 3023 619173
rect -960 619168 3023 619170
rect -960 619112 2962 619168
rect 3018 619112 3023 619168
rect -960 619110 3023 619112
rect -960 619020 480 619110
rect 2957 619107 3023 619110
rect 166612 618218 167194 618220
rect 168557 618218 168623 618221
rect 166612 618216 168623 618218
rect 166612 618160 168562 618216
rect 168618 618160 168623 618216
rect 167134 618158 168623 618160
rect 168557 618155 168623 618158
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 338246 612234 338252 612236
rect 336414 612204 338252 612234
rect 335892 612174 338252 612204
rect 335892 612144 336474 612174
rect 338246 612172 338252 612174
rect 338316 612234 338322 612236
rect 339401 612234 339467 612237
rect 338316 612232 339467 612234
rect 338316 612176 339406 612232
rect 339462 612176 339467 612232
rect 338316 612174 339467 612176
rect 338316 612172 338322 612174
rect 339401 612171 339467 612174
rect 407113 612234 407179 612237
rect 407113 612232 409522 612234
rect 407113 612176 407118 612232
rect 407174 612204 409522 612232
rect 407174 612176 410032 612204
rect 407113 612174 410032 612176
rect 407113 612171 407179 612174
rect 409462 612144 410032 612174
rect 338062 611010 338068 611012
rect 336414 610980 338068 611010
rect 335892 610950 338068 610980
rect 335892 610920 336474 610950
rect 338062 610948 338068 610950
rect 338132 611010 338138 611012
rect 339401 611010 339467 611013
rect 338132 611008 339467 611010
rect 338132 610952 339406 611008
rect 339462 610952 339467 611008
rect 338132 610950 339467 610952
rect 338132 610948 338138 610950
rect 339401 610947 339467 610950
rect 407113 611010 407179 611013
rect 407113 611008 409522 611010
rect 407113 610952 407118 611008
rect 407174 610980 409522 611008
rect 407174 610952 410032 610980
rect 407113 610950 410032 610952
rect 407113 610947 407179 610950
rect 409462 610920 410032 610950
rect 27429 609378 27495 609381
rect 27429 609376 30062 609378
rect 27429 609320 27434 609376
rect 27490 609320 30062 609376
rect 27429 609318 30062 609320
rect 27429 609315 27495 609318
rect 338297 609242 338363 609245
rect 336414 609240 338363 609242
rect 336414 609212 338302 609240
rect 335892 609184 338302 609212
rect 338358 609184 338363 609240
rect 335892 609182 338363 609184
rect 335892 609152 336474 609182
rect 338297 609179 338363 609182
rect 407113 609242 407179 609245
rect 407113 609240 409522 609242
rect 407113 609184 407118 609240
rect 407174 609212 409522 609240
rect 407174 609184 410032 609212
rect 407113 609182 410032 609184
rect 407113 609179 407179 609182
rect 409462 609152 410032 609182
rect 338113 608154 338179 608157
rect 336414 608152 338179 608154
rect 336414 608124 338118 608152
rect 335892 608096 338118 608124
rect 338174 608096 338179 608152
rect 335892 608094 338179 608096
rect 335892 608064 336474 608094
rect 338113 608091 338179 608094
rect 407113 608154 407179 608157
rect 407113 608152 409522 608154
rect 407113 608096 407118 608152
rect 407174 608124 409522 608152
rect 407174 608096 410032 608124
rect 407113 608094 410032 608096
rect 407113 608091 407179 608094
rect 409462 608064 410032 608094
rect 27337 607746 27403 607749
rect 27337 607744 30062 607746
rect 27337 607688 27342 607744
rect 27398 607688 30062 607744
rect 27337 607686 30062 607688
rect 27337 607683 27403 607686
rect 338389 606522 338455 606525
rect 336414 606520 338455 606522
rect 336414 606492 338394 606520
rect 335892 606464 338394 606492
rect 338450 606464 338455 606520
rect 335892 606462 338455 606464
rect 335892 606432 336474 606462
rect 338389 606459 338455 606462
rect 407113 606522 407179 606525
rect 407113 606520 409522 606522
rect 407113 606464 407118 606520
rect 407174 606492 409522 606520
rect 407174 606464 410032 606492
rect 407113 606462 410032 606464
rect 407113 606459 407179 606462
rect 409462 606432 410032 606462
rect 27521 606386 27587 606389
rect 27521 606384 30062 606386
rect 27521 606328 27526 606384
rect 27582 606328 30062 606384
rect 27521 606326 30062 606328
rect 27521 606323 27587 606326
rect -960 606114 480 606204
rect 3693 606114 3759 606117
rect -960 606112 3759 606114
rect -960 606056 3698 606112
rect 3754 606056 3759 606112
rect -960 606054 3759 606056
rect -960 605964 480 606054
rect 3693 606051 3759 606054
rect 339401 605570 339467 605573
rect 336414 605568 339467 605570
rect 336414 605540 339406 605568
rect 335892 605512 339406 605540
rect 339462 605512 339467 605568
rect 335892 605510 339467 605512
rect 335892 605480 336474 605510
rect 339401 605507 339467 605510
rect 407113 605570 407179 605573
rect 407113 605568 409522 605570
rect 407113 605512 407118 605568
rect 407174 605540 409522 605568
rect 407174 605512 410032 605540
rect 407113 605510 410032 605512
rect 407113 605507 407179 605510
rect 409462 605480 410032 605510
rect 27153 604890 27219 604893
rect 27153 604888 30062 604890
rect 27153 604832 27158 604888
rect 27214 604832 30062 604888
rect 27153 604830 30062 604832
rect 27153 604827 27219 604830
rect 583520 604060 584960 604300
rect 336733 603802 336799 603805
rect 339217 603802 339283 603805
rect 336414 603800 339283 603802
rect 336414 603772 336738 603800
rect 335892 603744 336738 603772
rect 336794 603744 339222 603800
rect 339278 603744 339283 603800
rect 335892 603742 339283 603744
rect 335892 603712 336474 603742
rect 336733 603739 336799 603742
rect 339217 603739 339283 603742
rect 407113 603802 407179 603805
rect 407113 603800 409522 603802
rect 407113 603744 407118 603800
rect 407174 603772 409522 603800
rect 407174 603744 410032 603772
rect 407113 603742 410032 603744
rect 407113 603739 407179 603742
rect 409462 603712 410032 603742
rect 27245 603666 27311 603669
rect 27245 603664 30062 603666
rect 27245 603608 27250 603664
rect 27306 603608 30062 603664
rect 27245 603606 30062 603608
rect 27245 603603 27311 603606
rect 166612 599994 167194 599996
rect 168925 599994 168991 599997
rect 166612 599992 168991 599994
rect 166612 599936 168930 599992
rect 168986 599936 168991 599992
rect 167134 599934 168991 599936
rect 168925 599931 168991 599934
rect 166612 598362 167194 598364
rect 169661 598362 169727 598365
rect 166612 598360 169727 598362
rect 166612 598304 169666 598360
rect 169722 598304 169727 598360
rect 167134 598302 169727 598304
rect 169661 598299 169727 598302
rect 166612 598090 167194 598092
rect 168741 598090 168807 598093
rect 166612 598088 168807 598090
rect 166612 598032 168746 598088
rect 168802 598032 168807 598088
rect 167134 598030 168807 598032
rect 168741 598027 168807 598030
rect 238661 594690 238727 594693
rect 506565 594690 506631 594693
rect 238661 594688 239506 594690
rect 238661 594632 238666 594688
rect 238722 594660 239506 594688
rect 506430 594688 506631 594690
rect 506430 594660 506570 594688
rect 238722 594632 240028 594660
rect 238661 594630 240028 594632
rect 238661 594627 238727 594630
rect 239446 594600 240028 594630
rect 505908 594632 506570 594660
rect 506626 594632 506631 594688
rect 505908 594630 506631 594632
rect 505908 594600 506490 594630
rect 506565 594627 506631 594630
rect -960 592908 480 593148
rect 238569 593058 238635 593061
rect 506473 593058 506539 593061
rect 238569 593056 239506 593058
rect 238569 593000 238574 593056
rect 238630 593028 239506 593056
rect 506430 593056 506539 593058
rect 506430 593028 506478 593056
rect 238630 593000 240028 593028
rect 238569 592998 240028 593000
rect 238569 592995 238635 592998
rect 239446 592968 240028 592998
rect 505908 593000 506478 593028
rect 506534 593000 506539 593056
rect 505908 592995 506539 593000
rect 505908 592968 506490 592995
rect 237189 591698 237255 591701
rect 507945 591698 508011 591701
rect 237189 591696 239506 591698
rect 237189 591640 237194 591696
rect 237250 591668 239506 591696
rect 506430 591696 508011 591698
rect 506430 591668 507950 591696
rect 237250 591640 240028 591668
rect 237189 591638 240028 591640
rect 237189 591635 237255 591638
rect 239446 591608 240028 591638
rect 505908 591640 507950 591668
rect 508006 591640 508011 591696
rect 505908 591638 508011 591640
rect 505908 591608 506490 591638
rect 507945 591635 508011 591638
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect 144784 589732 144790 589796
rect 144854 589794 144860 589796
rect 146008 589794 146014 589796
rect 144854 589734 146014 589794
rect 144854 589732 144860 589734
rect 146008 589732 146014 589734
rect 146078 589732 146084 589796
rect 43110 588100 43116 588164
rect 43180 588100 43186 588164
rect 63166 588100 63172 588164
rect 63236 588100 63242 588164
rect 73102 588100 73108 588164
rect 73172 588100 73178 588164
rect 83038 588100 83044 588164
rect 83108 588100 83114 588164
rect 85614 588100 85620 588164
rect 85684 588100 85690 588164
rect 95550 588100 95556 588164
rect 95620 588100 95626 588164
rect 103094 588100 103100 588164
rect 103164 588100 103170 588164
rect 109534 588100 109540 588164
rect 109604 588100 109610 588164
rect 112110 588100 112116 588164
rect 112180 588100 112186 588164
rect 113030 588100 113036 588164
rect 113100 588100 113106 588164
rect 115606 588100 115612 588164
rect 115676 588100 115682 588164
rect 122966 588100 122972 588164
rect 123036 588100 123042 588164
rect 129590 588100 129596 588164
rect 129660 588100 129666 588164
rect 133086 588100 133092 588164
rect 133156 588100 133162 588164
rect 143390 588100 143396 588164
rect 143460 588100 143466 588164
rect 149462 588100 149468 588164
rect 149532 588100 149538 588164
rect 43118 587893 43178 588100
rect 43069 587888 43178 587893
rect 43069 587832 43074 587888
rect 43130 587832 43178 587888
rect 43069 587830 43178 587832
rect 43529 587890 43595 587893
rect 60641 587892 60707 587893
rect 43662 587890 43668 587892
rect 43529 587888 43668 587890
rect 43529 587832 43534 587888
rect 43590 587832 43668 587888
rect 43529 587830 43668 587832
rect 43069 587827 43135 587830
rect 43529 587827 43595 587830
rect 43662 587828 43668 587830
rect 43732 587828 43738 587892
rect 60590 587890 60596 587892
rect 60550 587830 60596 587890
rect 60660 587888 60707 587892
rect 60702 587832 60707 587888
rect 60590 587828 60596 587830
rect 60660 587828 60707 587832
rect 60641 587827 60707 587828
rect 62941 587890 63007 587893
rect 63174 587890 63234 588100
rect 62941 587888 63234 587890
rect 62941 587832 62946 587888
rect 63002 587832 63234 587888
rect 62941 587830 63234 587832
rect 62941 587827 63007 587830
rect 68134 587828 68140 587892
rect 68204 587890 68210 587892
rect 68921 587890 68987 587893
rect 68204 587888 68987 587890
rect 68204 587832 68926 587888
rect 68982 587832 68987 587888
rect 68204 587830 68987 587832
rect 73110 587890 73170 588100
rect 74441 587890 74507 587893
rect 73110 587888 74507 587890
rect 73110 587832 74446 587888
rect 74502 587832 74507 587888
rect 73110 587830 74507 587832
rect 83046 587890 83106 588100
rect 83825 587890 83891 587893
rect 83046 587888 83891 587890
rect 83046 587832 83830 587888
rect 83886 587832 83891 587888
rect 83046 587830 83891 587832
rect 85622 587890 85682 588100
rect 86401 587890 86467 587893
rect 88241 587892 88307 587893
rect 88190 587890 88196 587892
rect 85622 587888 86467 587890
rect 85622 587832 86406 587888
rect 86462 587832 86467 587888
rect 85622 587830 86467 587832
rect 88150 587830 88196 587890
rect 88260 587888 88307 587892
rect 88302 587832 88307 587888
rect 68204 587828 68210 587830
rect 68921 587827 68987 587830
rect 74441 587827 74507 587830
rect 83825 587827 83891 587830
rect 86401 587827 86467 587830
rect 88190 587828 88196 587830
rect 88260 587828 88307 587832
rect 88241 587827 88307 587828
rect 95233 587890 95299 587893
rect 95558 587890 95618 588100
rect 103102 587893 103162 588100
rect 109542 587893 109602 588100
rect 95233 587888 95618 587890
rect 95233 587832 95238 587888
rect 95294 587832 95618 587888
rect 95233 587830 95618 587832
rect 95233 587827 95299 587830
rect 98310 587828 98316 587892
rect 98380 587890 98386 587892
rect 99189 587890 99255 587893
rect 100569 587892 100635 587893
rect 100518 587890 100524 587892
rect 98380 587888 99255 587890
rect 98380 587832 99194 587888
rect 99250 587832 99255 587888
rect 98380 587830 99255 587832
rect 100478 587830 100524 587890
rect 100588 587888 100635 587892
rect 100630 587832 100635 587888
rect 98380 587828 98386 587830
rect 99189 587827 99255 587830
rect 100518 587828 100524 587830
rect 100588 587828 100635 587832
rect 103102 587888 103211 587893
rect 103102 587832 103150 587888
rect 103206 587832 103211 587888
rect 103102 587830 103211 587832
rect 100569 587827 100635 587828
rect 103145 587827 103211 587830
rect 105077 587890 105143 587893
rect 105302 587890 105308 587892
rect 105077 587888 105308 587890
rect 105077 587832 105082 587888
rect 105138 587832 105308 587888
rect 105077 587830 105308 587832
rect 105077 587827 105143 587830
rect 105302 587828 105308 587830
rect 105372 587828 105378 587892
rect 106273 587890 106339 587893
rect 107326 587890 107332 587892
rect 106273 587888 107332 587890
rect 106273 587832 106278 587888
rect 106334 587832 107332 587888
rect 106273 587830 107332 587832
rect 106273 587827 106339 587830
rect 107326 587828 107332 587830
rect 107396 587828 107402 587892
rect 107745 587890 107811 587893
rect 108430 587890 108436 587892
rect 107745 587888 108436 587890
rect 107745 587832 107750 587888
rect 107806 587832 108436 587888
rect 107745 587830 108436 587832
rect 107745 587827 107811 587830
rect 108430 587828 108436 587830
rect 108500 587828 108506 587892
rect 109493 587888 109602 587893
rect 110505 587892 110571 587893
rect 110454 587890 110460 587892
rect 109493 587832 109498 587888
rect 109554 587832 109602 587888
rect 109493 587830 109602 587832
rect 110414 587830 110460 587890
rect 110524 587888 110571 587892
rect 110566 587832 110571 587888
rect 109493 587827 109559 587830
rect 110454 587828 110460 587830
rect 110524 587828 110571 587832
rect 110822 587828 110828 587892
rect 110892 587890 110898 587892
rect 111609 587890 111675 587893
rect 110892 587888 111675 587890
rect 110892 587832 111614 587888
rect 111670 587832 111675 587888
rect 110892 587830 111675 587832
rect 112118 587890 112178 588100
rect 113038 587893 113098 588100
rect 112529 587890 112595 587893
rect 112118 587888 112595 587890
rect 112118 587832 112534 587888
rect 112590 587832 112595 587888
rect 112118 587830 112595 587832
rect 113038 587888 113147 587893
rect 113038 587832 113086 587888
rect 113142 587832 113147 587888
rect 113038 587830 113147 587832
rect 110892 587828 110898 587830
rect 110505 587827 110571 587828
rect 111609 587827 111675 587830
rect 112529 587827 112595 587830
rect 113081 587827 113147 587830
rect 113817 587890 113883 587893
rect 114318 587890 114324 587892
rect 113817 587888 114324 587890
rect 113817 587832 113822 587888
rect 113878 587832 114324 587888
rect 113817 587830 114324 587832
rect 113817 587827 113883 587830
rect 114318 587828 114324 587830
rect 114388 587828 114394 587892
rect 114829 587890 114895 587893
rect 115238 587890 115244 587892
rect 114829 587888 115244 587890
rect 114829 587832 114834 587888
rect 114890 587832 115244 587888
rect 114829 587830 115244 587832
rect 114829 587827 114895 587830
rect 115238 587828 115244 587830
rect 115308 587828 115314 587892
rect 113766 587692 113772 587756
rect 113836 587754 113842 587756
rect 114369 587754 114435 587757
rect 113836 587752 114435 587754
rect 113836 587696 114374 587752
rect 114430 587696 114435 587752
rect 113836 587694 114435 587696
rect 113836 587692 113842 587694
rect 114369 587691 114435 587694
rect 114553 587754 114619 587757
rect 115614 587754 115674 588100
rect 116710 587828 116716 587892
rect 116780 587890 116786 587892
rect 117129 587890 117195 587893
rect 116780 587888 117195 587890
rect 116780 587832 117134 587888
rect 117190 587832 117195 587888
rect 116780 587830 117195 587832
rect 116780 587828 116786 587830
rect 117129 587827 117195 587830
rect 118918 587828 118924 587892
rect 118988 587890 118994 587892
rect 119797 587890 119863 587893
rect 120257 587892 120323 587893
rect 120206 587890 120212 587892
rect 118988 587888 119863 587890
rect 118988 587832 119802 587888
rect 119858 587832 119863 587888
rect 118988 587830 119863 587832
rect 120166 587830 120212 587890
rect 120276 587888 120323 587892
rect 120318 587832 120323 587888
rect 118988 587828 118994 587830
rect 119797 587827 119863 587830
rect 120206 587828 120212 587830
rect 120276 587828 120323 587832
rect 120257 587827 120323 587828
rect 120533 587890 120599 587893
rect 122649 587892 122715 587893
rect 121310 587890 121316 587892
rect 120533 587888 121316 587890
rect 120533 587832 120538 587888
rect 120594 587832 121316 587888
rect 120533 587830 121316 587832
rect 120533 587827 120599 587830
rect 121310 587828 121316 587830
rect 121380 587828 121386 587892
rect 122598 587890 122604 587892
rect 122558 587830 122604 587890
rect 122668 587888 122715 587892
rect 122710 587832 122715 587888
rect 122598 587828 122604 587830
rect 122668 587828 122715 587832
rect 122649 587827 122715 587828
rect 122833 587890 122899 587893
rect 122974 587890 123034 588100
rect 129598 587893 129658 588100
rect 133094 587893 133154 588100
rect 143398 587893 143458 588100
rect 149470 587893 149530 588100
rect 122833 587888 123034 587890
rect 122833 587832 122838 587888
rect 122894 587832 123034 587888
rect 122833 587830 123034 587832
rect 122833 587827 122899 587830
rect 124806 587828 124812 587892
rect 124876 587890 124882 587892
rect 125041 587890 125107 587893
rect 124876 587888 125107 587890
rect 124876 587832 125046 587888
rect 125102 587832 125107 587888
rect 124876 587830 125107 587832
rect 124876 587828 124882 587830
rect 125041 587827 125107 587830
rect 126278 587828 126284 587892
rect 126348 587890 126354 587892
rect 126881 587890 126947 587893
rect 126348 587888 126947 587890
rect 126348 587832 126886 587888
rect 126942 587832 126947 587888
rect 126348 587830 126947 587832
rect 126348 587828 126354 587830
rect 126881 587827 126947 587830
rect 128486 587828 128492 587892
rect 128556 587890 128562 587892
rect 129365 587890 129431 587893
rect 128556 587888 129431 587890
rect 128556 587832 129370 587888
rect 129426 587832 129431 587888
rect 128556 587830 129431 587832
rect 129598 587888 129707 587893
rect 129598 587832 129646 587888
rect 129702 587832 129707 587888
rect 129598 587830 129707 587832
rect 128556 587828 128562 587830
rect 129365 587827 129431 587830
rect 129641 587827 129707 587830
rect 130561 587890 130627 587893
rect 130694 587890 130700 587892
rect 130561 587888 130700 587890
rect 130561 587832 130566 587888
rect 130622 587832 130700 587888
rect 130561 587830 130700 587832
rect 130561 587827 130627 587830
rect 130694 587828 130700 587830
rect 130764 587828 130770 587892
rect 131113 587890 131179 587893
rect 131614 587890 131620 587892
rect 131113 587888 131620 587890
rect 131113 587832 131118 587888
rect 131174 587832 131620 587888
rect 131113 587830 131620 587832
rect 131113 587827 131179 587830
rect 131614 587828 131620 587830
rect 131684 587828 131690 587892
rect 132585 587890 132651 587893
rect 132718 587890 132724 587892
rect 132585 587888 132724 587890
rect 132585 587832 132590 587888
rect 132646 587832 132724 587888
rect 132585 587830 132724 587832
rect 132585 587827 132651 587830
rect 132718 587828 132724 587830
rect 132788 587828 132794 587892
rect 133094 587888 133203 587893
rect 133094 587832 133142 587888
rect 133198 587832 133203 587888
rect 133094 587830 133203 587832
rect 133137 587827 133203 587830
rect 136214 587828 136220 587892
rect 136284 587890 136290 587892
rect 136449 587890 136515 587893
rect 137921 587892 137987 587893
rect 137870 587890 137876 587892
rect 136284 587888 136515 587890
rect 136284 587832 136454 587888
rect 136510 587832 136515 587888
rect 136284 587830 136515 587832
rect 137830 587830 137876 587890
rect 137940 587888 137987 587892
rect 137982 587832 137987 587888
rect 136284 587828 136290 587830
rect 136449 587827 136515 587830
rect 137870 587828 137876 587830
rect 137940 587828 137987 587832
rect 138238 587828 138244 587892
rect 138308 587890 138314 587892
rect 139301 587890 139367 587893
rect 140129 587892 140195 587893
rect 142705 587892 142771 587893
rect 140078 587890 140084 587892
rect 138308 587888 139367 587890
rect 138308 587832 139306 587888
rect 139362 587832 139367 587888
rect 138308 587830 139367 587832
rect 140038 587830 140084 587890
rect 140148 587888 140195 587892
rect 142654 587890 142660 587892
rect 140190 587832 140195 587888
rect 138308 587828 138314 587830
rect 137921 587827 137987 587828
rect 139301 587827 139367 587830
rect 140078 587828 140084 587830
rect 140148 587828 140195 587832
rect 142614 587830 142660 587890
rect 142724 587888 142771 587892
rect 142766 587832 142771 587888
rect 142654 587828 142660 587830
rect 142724 587828 142771 587832
rect 143398 587888 143507 587893
rect 143398 587832 143446 587888
rect 143502 587832 143507 587888
rect 143398 587830 143507 587832
rect 140129 587827 140195 587828
rect 142705 587827 142771 587828
rect 143441 587827 143507 587830
rect 147070 587828 147076 587892
rect 147140 587890 147146 587892
rect 147673 587890 147739 587893
rect 148358 587890 148364 587892
rect 147140 587888 148364 587890
rect 147140 587832 147678 587888
rect 147734 587832 148364 587888
rect 147140 587830 148364 587832
rect 147140 587828 147146 587830
rect 147673 587827 147739 587830
rect 148358 587828 148364 587830
rect 148428 587828 148434 587892
rect 149470 587888 149579 587893
rect 149470 587832 149518 587888
rect 149574 587832 149579 587888
rect 149470 587830 149579 587832
rect 149513 587827 149579 587830
rect 150566 587828 150572 587892
rect 150636 587890 150642 587892
rect 150709 587890 150775 587893
rect 150636 587888 150775 587890
rect 150636 587832 150714 587888
rect 150770 587832 150775 587888
rect 150636 587830 150775 587832
rect 150636 587828 150642 587830
rect 150709 587827 150775 587830
rect 114553 587752 115674 587754
rect 114553 587696 114558 587752
rect 114614 587696 115674 587752
rect 114553 587694 115674 587696
rect 120165 587754 120231 587757
rect 120574 587754 120580 587756
rect 120165 587752 120580 587754
rect 120165 587696 120170 587752
rect 120226 587696 120580 587752
rect 120165 587694 120580 587696
rect 114553 587691 114619 587694
rect 120165 587691 120231 587694
rect 120574 587692 120580 587694
rect 120644 587692 120650 587756
rect 130510 587692 130516 587756
rect 130580 587754 130586 587756
rect 131021 587754 131087 587757
rect 130580 587752 131087 587754
rect 130580 587696 131026 587752
rect 131082 587696 131087 587752
rect 130580 587694 131087 587696
rect 130580 587692 130586 587694
rect 131021 587691 131087 587694
rect 134190 587692 134196 587756
rect 134260 587754 134266 587756
rect 166942 587754 166948 587756
rect 134260 587694 166948 587754
rect 134260 587692 134266 587694
rect 166942 587692 166948 587694
rect 167012 587692 167018 587756
rect 135294 587556 135300 587620
rect 135364 587618 135370 587620
rect 170070 587618 170076 587620
rect 135364 587558 170076 587618
rect 135364 587556 135370 587558
rect 170070 587556 170076 587558
rect 170140 587556 170146 587620
rect 127198 587420 127204 587484
rect 127268 587482 127274 587484
rect 173157 587482 173223 587485
rect 127268 587480 173223 587482
rect 127268 587424 173162 587480
rect 173218 587424 173223 587480
rect 127268 587422 173223 587424
rect 127268 587420 127274 587422
rect 173157 587419 173223 587422
rect 123702 587284 123708 587348
rect 123772 587346 123778 587348
rect 170254 587346 170260 587348
rect 123772 587286 170260 587346
rect 123772 587284 123778 587286
rect 170254 587284 170260 587286
rect 170324 587284 170330 587348
rect 172145 587210 172211 587213
rect 122790 587208 172211 587210
rect 122790 587152 172150 587208
rect 172206 587152 172211 587208
rect 122790 587150 172211 587152
rect 117814 587012 117820 587076
rect 117884 587074 117890 587076
rect 122790 587074 122850 587150
rect 172145 587147 172211 587150
rect 117884 587014 122850 587074
rect 136541 587076 136607 587077
rect 139025 587076 139091 587077
rect 136541 587072 136588 587076
rect 136652 587074 136658 587076
rect 138974 587074 138980 587076
rect 136541 587016 136546 587072
rect 117884 587012 117890 587014
rect 136541 587012 136588 587016
rect 136652 587014 136698 587074
rect 138934 587014 138980 587074
rect 139044 587072 139091 587076
rect 139086 587016 139091 587072
rect 136652 587012 136658 587014
rect 138974 587012 138980 587014
rect 139044 587012 139091 587016
rect 136541 587011 136607 587012
rect 139025 587011 139091 587012
rect 70710 586666 70716 586668
rect 70350 586606 70716 586666
rect 64873 586532 64939 586533
rect 64822 586468 64828 586532
rect 64892 586530 64939 586532
rect 64892 586528 64984 586530
rect 64934 586472 64984 586528
rect 64892 586470 64984 586472
rect 64892 586468 64939 586470
rect 64873 586467 64939 586468
rect 70350 586394 70410 586606
rect 70710 586604 70716 586606
rect 70780 586604 70786 586668
rect 75310 586666 75316 586668
rect 74582 586606 75316 586666
rect 71681 586394 71747 586397
rect 70350 586392 71747 586394
rect 70350 586336 71686 586392
rect 71742 586336 71747 586392
rect 70350 586334 71747 586336
rect 74582 586394 74642 586606
rect 75310 586604 75316 586606
rect 75380 586604 75386 586668
rect 78070 586666 78076 586668
rect 77342 586606 78076 586666
rect 75821 586394 75887 586397
rect 74582 586392 75887 586394
rect 74582 586336 75826 586392
rect 75882 586336 75887 586392
rect 74582 586334 75887 586336
rect 77342 586394 77402 586606
rect 78070 586604 78076 586606
rect 78140 586604 78146 586668
rect 80646 586666 80652 586668
rect 80102 586606 80652 586666
rect 78581 586394 78647 586397
rect 77342 586392 78647 586394
rect 77342 586336 78586 586392
rect 78642 586336 78647 586392
rect 77342 586334 78647 586336
rect 80102 586394 80162 586606
rect 80646 586604 80652 586606
rect 80716 586604 80722 586668
rect 90582 586666 90588 586668
rect 90038 586606 90588 586666
rect 81341 586394 81407 586397
rect 80102 586392 81407 586394
rect 80102 586336 81346 586392
rect 81402 586336 81407 586392
rect 80102 586334 81407 586336
rect 90038 586394 90098 586606
rect 90582 586604 90588 586606
rect 90652 586604 90658 586668
rect 92790 586666 92796 586668
rect 92614 586606 92796 586666
rect 91001 586394 91067 586397
rect 90038 586392 91067 586394
rect 90038 586336 91006 586392
rect 91062 586336 91067 586392
rect 90038 586334 91067 586336
rect 92614 586394 92674 586606
rect 92790 586604 92796 586606
rect 92860 586604 92866 586668
rect 108062 586666 108068 586668
rect 107886 586606 108068 586666
rect 93761 586394 93827 586397
rect 92614 586392 93827 586394
rect 92614 586336 93766 586392
rect 93822 586336 93827 586392
rect 92614 586334 93827 586336
rect 107886 586394 107946 586606
rect 108062 586604 108068 586606
rect 108132 586604 108138 586668
rect 118182 586666 118188 586668
rect 117270 586606 118188 586666
rect 108941 586394 109007 586397
rect 107886 586392 109007 586394
rect 107886 586336 108946 586392
rect 109002 586336 109007 586392
rect 107886 586334 109007 586336
rect 117270 586394 117330 586606
rect 118182 586604 118188 586606
rect 118252 586604 118258 586668
rect 125358 586666 125364 586668
rect 124262 586606 125364 586666
rect 118601 586394 118667 586397
rect 117270 586392 118667 586394
rect 117270 586336 118606 586392
rect 118662 586336 118667 586392
rect 117270 586334 118667 586336
rect 124262 586394 124322 586606
rect 125358 586604 125364 586606
rect 125428 586604 125434 586668
rect 128118 586666 128124 586668
rect 127022 586606 128124 586666
rect 125501 586394 125567 586397
rect 124262 586392 125567 586394
rect 124262 586336 125506 586392
rect 125562 586336 125567 586392
rect 124262 586334 125567 586336
rect 127022 586394 127082 586606
rect 128118 586604 128124 586606
rect 128188 586604 128194 586668
rect 140998 586666 141004 586668
rect 140822 586606 141004 586666
rect 128261 586394 128327 586397
rect 127022 586392 128327 586394
rect 127022 586336 128266 586392
rect 128322 586336 128327 586392
rect 127022 586334 128327 586336
rect 140822 586394 140882 586606
rect 140998 586604 141004 586606
rect 141068 586604 141074 586668
rect 142061 586394 142127 586397
rect 140822 586392 142127 586394
rect 140822 586336 142066 586392
rect 142122 586336 142127 586392
rect 140822 586334 142127 586336
rect 71681 586331 71747 586334
rect 75821 586331 75887 586334
rect 78581 586331 78647 586334
rect 81341 586331 81407 586334
rect 91001 586331 91067 586334
rect 93761 586331 93827 586334
rect 108941 586331 109007 586334
rect 118601 586331 118667 586334
rect 125501 586331 125567 586334
rect 128261 586331 128327 586334
rect 142061 586331 142127 586334
rect 336917 585306 336983 585309
rect 339217 585306 339283 585309
rect 336414 585304 339283 585306
rect 336414 585276 336922 585304
rect 335892 585248 336922 585276
rect 336978 585248 339222 585304
rect 339278 585248 339283 585304
rect 335892 585246 339283 585248
rect 335892 585216 336474 585246
rect 336917 585243 336983 585246
rect 339217 585243 339283 585246
rect 407113 585306 407179 585309
rect 407113 585304 409522 585306
rect 407113 585248 407118 585304
rect 407174 585276 409522 585304
rect 407174 585248 410032 585276
rect 407113 585246 410032 585248
rect 407113 585243 407179 585246
rect 409462 585216 410032 585246
rect 120257 584898 120323 584901
rect 168414 584898 168420 584900
rect 120257 584896 168420 584898
rect 120257 584840 120262 584896
rect 120318 584840 168420 584896
rect 120257 584838 168420 584840
rect 120257 584835 120323 584838
rect 168414 584836 168420 584838
rect 168484 584836 168490 584900
rect 119797 584762 119863 584765
rect 167126 584762 167132 584764
rect 119797 584760 167132 584762
rect 119797 584704 119802 584760
rect 119858 584704 167132 584760
rect 119797 584702 167132 584704
rect 119797 584699 119863 584702
rect 167126 584700 167132 584702
rect 167196 584700 167202 584764
rect 114369 584626 114435 584629
rect 171133 584626 171199 584629
rect 114369 584624 171199 584626
rect 114369 584568 114374 584624
rect 114430 584568 171138 584624
rect 171194 584568 171199 584624
rect 114369 584566 171199 584568
rect 114369 584563 114435 584566
rect 171133 584563 171199 584566
rect 111609 584490 111675 584493
rect 172646 584490 172652 584492
rect 111609 584488 172652 584490
rect 111609 584432 111614 584488
rect 111670 584432 172652 584488
rect 111609 584430 172652 584432
rect 111609 584427 111675 584430
rect 172646 584428 172652 584430
rect 172716 584428 172722 584492
rect 112529 584354 112595 584357
rect 173985 584354 174051 584357
rect 112529 584352 174051 584354
rect 112529 584296 112534 584352
rect 112590 584296 173990 584352
rect 174046 584296 174051 584352
rect 112529 584294 174051 584296
rect 112529 584291 112595 584294
rect 173985 584291 174051 584294
rect 337377 583674 337443 583677
rect 339401 583674 339467 583677
rect 336414 583672 339467 583674
rect 336414 583644 337382 583672
rect 335892 583616 337382 583644
rect 337438 583616 339406 583672
rect 339462 583616 339467 583672
rect 335892 583614 339467 583616
rect 335892 583584 336474 583614
rect 337377 583611 337443 583614
rect 339401 583611 339467 583614
rect 407113 583674 407179 583677
rect 407113 583672 409522 583674
rect 407113 583616 407118 583672
rect 407174 583644 409522 583672
rect 407174 583616 410032 583644
rect 407113 583614 410032 583616
rect 407113 583611 407179 583614
rect 409462 583584 410032 583614
rect 107745 581770 107811 581773
rect 168598 581770 168604 581772
rect 107745 581768 168604 581770
rect 107745 581712 107750 581768
rect 107806 581712 168604 581768
rect 107745 581710 168604 581712
rect 107745 581707 107811 581710
rect 168598 581708 168604 581710
rect 168668 581708 168674 581772
rect 106273 581634 106339 581637
rect 167678 581634 167684 581636
rect 106273 581632 167684 581634
rect 106273 581576 106278 581632
rect 106334 581576 167684 581632
rect 106273 581574 167684 581576
rect 106273 581571 106339 581574
rect 167678 581572 167684 581574
rect 167748 581572 167754 581636
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 492673 577828 492739 577829
rect 252502 577764 252508 577828
rect 252572 577826 252578 577828
rect 252920 577826 252926 577828
rect 252572 577766 252926 577826
rect 252572 577764 252578 577766
rect 252920 577764 252926 577766
rect 252990 577764 252996 577828
rect 284886 577764 284892 577828
rect 284956 577826 284962 577828
rect 285288 577826 285294 577828
rect 284956 577766 285294 577826
rect 284956 577764 284962 577766
rect 285288 577764 285294 577766
rect 285358 577764 285364 577828
rect 445150 577764 445156 577828
rect 445220 577826 445226 577828
rect 445496 577826 445502 577828
rect 445220 577766 445502 577826
rect 445220 577764 445226 577766
rect 445496 577764 445502 577766
rect 445566 577764 445572 577828
rect 492673 577826 492694 577828
rect 492602 577824 492694 577826
rect 492602 577768 492678 577824
rect 492602 577766 492694 577768
rect 492673 577764 492694 577766
rect 492758 577764 492764 577828
rect 493096 577764 493102 577828
rect 493166 577764 493172 577828
rect 492673 577763 492739 577764
rect 492622 577628 492628 577692
rect 492692 577690 492698 577692
rect 493104 577690 493164 577764
rect 492692 577630 493164 577690
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 492692 577628 492698 577630
rect 580165 577627 580231 577630
rect 280102 577492 280108 577556
rect 280172 577554 280178 577556
rect 281480 577554 281486 577556
rect 280172 577494 281486 577554
rect 280172 577492 280178 577494
rect 281480 577492 281486 577494
rect 281550 577492 281556 577556
rect 583520 577540 584960 577630
rect 441797 577012 441863 577013
rect 462865 577012 462931 577013
rect 441797 577010 441844 577012
rect 441752 577008 441844 577010
rect 441752 576952 441802 577008
rect 441752 576950 441844 576952
rect 441797 576948 441844 576950
rect 441908 576948 441914 577012
rect 462814 576948 462820 577012
rect 462884 577010 462931 577012
rect 462884 577008 462976 577010
rect 462926 576952 462976 577008
rect 462884 576950 462976 576952
rect 462884 576948 462931 576950
rect 441797 576947 441863 576948
rect 462865 576947 462931 576948
rect 492949 576876 493015 576877
rect 492949 576874 492996 576876
rect 492904 576872 492996 576874
rect 492904 576816 492954 576872
rect 492904 576814 492996 576816
rect 492949 576812 492996 576814
rect 493060 576812 493066 576876
rect 492949 576811 493015 576812
rect 253105 576196 253171 576197
rect 292481 576196 292547 576197
rect 455505 576196 455571 576197
rect 253054 576194 253060 576196
rect 253014 576134 253060 576194
rect 253124 576192 253171 576196
rect 292430 576194 292436 576196
rect 253166 576136 253171 576192
rect 253054 576132 253060 576134
rect 253124 576132 253171 576136
rect 292390 576134 292436 576194
rect 292500 576192 292547 576196
rect 292542 576136 292547 576192
rect 292430 576132 292436 576134
rect 292500 576132 292547 576136
rect 455454 576132 455460 576196
rect 455524 576194 455571 576196
rect 459277 576196 459343 576197
rect 459277 576194 459324 576196
rect 455524 576192 455616 576194
rect 455566 576136 455616 576192
rect 455524 576134 455616 576136
rect 459232 576192 459324 576194
rect 459232 576136 459282 576192
rect 459232 576134 459324 576136
rect 455524 576132 455571 576134
rect 253105 576131 253171 576132
rect 292481 576131 292547 576132
rect 455505 576131 455571 576132
rect 459277 576132 459324 576134
rect 459388 576132 459394 576196
rect 468477 576194 468543 576197
rect 469254 576194 469260 576196
rect 468477 576192 469260 576194
rect 468477 576136 468482 576192
rect 468538 576136 469260 576192
rect 468477 576134 469260 576136
rect 459277 576131 459343 576132
rect 468477 576131 468543 576134
rect 469254 576132 469260 576134
rect 469324 576132 469330 576196
rect 341558 575996 341564 576060
rect 341628 576058 341634 576060
rect 506565 576058 506631 576061
rect 341628 576056 506631 576058
rect 341628 576000 506570 576056
rect 506626 576000 506631 576056
rect 341628 575998 506631 576000
rect 341628 575996 341634 575998
rect 506565 575995 506631 575998
rect 284201 575380 284267 575381
rect 285305 575380 285371 575381
rect 286593 575380 286659 575381
rect 284150 575378 284156 575380
rect 284110 575318 284156 575378
rect 284220 575376 284267 575380
rect 285254 575378 285260 575380
rect 284262 575320 284267 575376
rect 284150 575316 284156 575318
rect 284220 575316 284267 575320
rect 285214 575318 285260 575378
rect 285324 575376 285371 575380
rect 286542 575378 286548 575380
rect 285366 575320 285371 575376
rect 285254 575316 285260 575318
rect 285324 575316 285371 575320
rect 286502 575318 286548 575378
rect 286612 575376 286659 575380
rect 286654 575320 286659 575376
rect 286542 575316 286548 575318
rect 286612 575316 286659 575320
rect 287646 575316 287652 575380
rect 287716 575378 287722 575380
rect 287881 575378 287947 575381
rect 287716 575376 287947 575378
rect 287716 575320 287886 575376
rect 287942 575320 287947 575376
rect 287716 575318 287947 575320
rect 287716 575316 287722 575318
rect 284201 575315 284267 575316
rect 285305 575315 285371 575316
rect 286593 575315 286659 575316
rect 287881 575315 287947 575318
rect 297030 575316 297036 575380
rect 297100 575378 297106 575380
rect 297909 575378 297975 575381
rect 297100 575376 297975 575378
rect 297100 575320 297914 575376
rect 297970 575320 297975 575376
rect 297100 575318 297975 575320
rect 297100 575316 297106 575318
rect 297909 575315 297975 575318
rect 300526 575316 300532 575380
rect 300596 575378 300602 575380
rect 300669 575378 300735 575381
rect 300596 575376 300735 575378
rect 300596 575320 300674 575376
rect 300730 575320 300735 575376
rect 300596 575318 300735 575320
rect 300596 575316 300602 575318
rect 300669 575315 300735 575318
rect 301630 575316 301636 575380
rect 301700 575378 301706 575380
rect 301865 575378 301931 575381
rect 301700 575376 301931 575378
rect 301700 575320 301870 575376
rect 301926 575320 301931 575376
rect 301700 575318 301931 575320
rect 301700 575316 301706 575318
rect 301865 575315 301931 575318
rect 302734 575316 302740 575380
rect 302804 575378 302810 575380
rect 302877 575378 302943 575381
rect 302804 575376 302943 575378
rect 302804 575320 302882 575376
rect 302938 575320 302943 575376
rect 302804 575318 302943 575320
rect 302804 575316 302810 575318
rect 302877 575315 302943 575318
rect 304206 575316 304212 575380
rect 304276 575378 304282 575380
rect 304625 575378 304691 575381
rect 304276 575376 304691 575378
rect 304276 575320 304630 575376
rect 304686 575320 304691 575376
rect 304276 575318 304691 575320
rect 304276 575316 304282 575318
rect 304625 575315 304691 575318
rect 305126 575316 305132 575380
rect 305196 575378 305202 575380
rect 305545 575378 305611 575381
rect 306281 575380 306347 575381
rect 307569 575380 307635 575381
rect 320449 575380 320515 575381
rect 330201 575380 330267 575381
rect 306230 575378 306236 575380
rect 305196 575376 305611 575378
rect 305196 575320 305550 575376
rect 305606 575320 305611 575376
rect 305196 575318 305611 575320
rect 306190 575318 306236 575378
rect 306300 575376 306347 575380
rect 307518 575378 307524 575380
rect 306342 575320 306347 575376
rect 305196 575316 305202 575318
rect 305545 575315 305611 575318
rect 306230 575316 306236 575318
rect 306300 575316 306347 575320
rect 307478 575318 307524 575378
rect 307588 575376 307635 575380
rect 320398 575378 320404 575380
rect 307630 575320 307635 575376
rect 307518 575316 307524 575318
rect 307588 575316 307635 575320
rect 320358 575318 320404 575378
rect 320468 575376 320515 575380
rect 330150 575378 330156 575380
rect 320510 575320 320515 575376
rect 320398 575316 320404 575318
rect 320468 575316 320515 575320
rect 330110 575318 330156 575378
rect 330220 575376 330267 575380
rect 330262 575320 330267 575376
rect 330150 575316 330156 575318
rect 330220 575316 330267 575320
rect 306281 575315 306347 575316
rect 307569 575315 307635 575316
rect 320449 575315 320515 575316
rect 330201 575315 330267 575316
rect 330477 575378 330543 575381
rect 336958 575378 336964 575380
rect 330477 575376 336964 575378
rect 330477 575320 330482 575376
rect 330538 575320 336964 575376
rect 330477 575318 336964 575320
rect 330477 575315 330543 575318
rect 336958 575316 336964 575318
rect 337028 575378 337034 575380
rect 338021 575378 338087 575381
rect 415393 575380 415459 575381
rect 337028 575376 338087 575378
rect 337028 575320 338026 575376
rect 338082 575320 338087 575376
rect 337028 575318 338087 575320
rect 337028 575316 337034 575318
rect 338021 575315 338087 575318
rect 415342 575316 415348 575380
rect 415412 575378 415459 575380
rect 425053 575378 425119 575381
rect 425278 575378 425284 575380
rect 415412 575376 415504 575378
rect 415454 575320 415504 575376
rect 415412 575318 415504 575320
rect 425053 575376 425284 575378
rect 425053 575320 425058 575376
rect 425114 575320 425284 575376
rect 425053 575318 425284 575320
rect 415412 575316 415459 575318
rect 415393 575315 415459 575316
rect 425053 575315 425119 575318
rect 425278 575316 425284 575318
rect 425348 575316 425354 575380
rect 284385 575242 284451 575245
rect 284886 575242 284892 575244
rect 284385 575240 284892 575242
rect 284385 575184 284390 575240
rect 284446 575184 284892 575240
rect 284385 575182 284892 575184
rect 284385 575179 284451 575182
rect 284886 575180 284892 575182
rect 284956 575180 284962 575244
rect 289813 575242 289879 575245
rect 293953 575244 294019 575245
rect 290222 575242 290228 575244
rect 289813 575240 290228 575242
rect 289813 575184 289818 575240
rect 289874 575184 290228 575240
rect 289813 575182 290228 575184
rect 289813 575179 289879 575182
rect 290222 575180 290228 575182
rect 290292 575180 290298 575244
rect 293902 575180 293908 575244
rect 293972 575242 294019 575244
rect 293972 575240 294064 575242
rect 294014 575184 294064 575240
rect 293972 575182 294064 575184
rect 293972 575180 294019 575182
rect 314510 575180 314516 575244
rect 314580 575242 314586 575244
rect 337561 575242 337627 575245
rect 314580 575240 337627 575242
rect 314580 575184 337566 575240
rect 337622 575184 337627 575240
rect 314580 575182 337627 575184
rect 314580 575180 314586 575182
rect 293953 575179 294019 575180
rect 337561 575179 337627 575182
rect 426433 575242 426499 575245
rect 426750 575242 426756 575244
rect 426433 575240 426756 575242
rect 426433 575184 426438 575240
rect 426494 575184 426756 575240
rect 426433 575182 426756 575184
rect 426433 575179 426499 575182
rect 426750 575180 426756 575182
rect 426820 575180 426826 575244
rect 437473 575242 437539 575245
rect 438342 575242 438348 575244
rect 437473 575240 438348 575242
rect 437473 575184 437478 575240
rect 437534 575184 438348 575240
rect 437473 575182 438348 575184
rect 437473 575179 437539 575182
rect 438342 575180 438348 575182
rect 438412 575180 438418 575244
rect 466453 575242 466519 575245
rect 467598 575242 467604 575244
rect 466453 575240 467604 575242
rect 466453 575184 466458 575240
rect 466514 575184 467604 575240
rect 466453 575182 467604 575184
rect 466453 575179 466519 575182
rect 467598 575180 467604 575182
rect 467668 575180 467674 575244
rect 280153 575108 280219 575109
rect 280102 575044 280108 575108
rect 280172 575106 280219 575108
rect 291193 575106 291259 575109
rect 291510 575106 291516 575108
rect 280172 575104 280264 575106
rect 280214 575048 280264 575104
rect 280172 575046 280264 575048
rect 291193 575104 291516 575106
rect 291193 575048 291198 575104
rect 291254 575048 291516 575104
rect 291193 575046 291516 575048
rect 280172 575044 280219 575046
rect 280153 575043 280219 575044
rect 291193 575043 291259 575046
rect 291510 575044 291516 575046
rect 291580 575044 291586 575108
rect 293953 575106 294019 575109
rect 295190 575106 295196 575108
rect 293953 575104 295196 575106
rect 293953 575048 293958 575104
rect 294014 575048 295196 575104
rect 293953 575046 295196 575048
rect 293953 575043 294019 575046
rect 295190 575044 295196 575046
rect 295260 575044 295266 575108
rect 312670 575044 312676 575108
rect 312740 575106 312746 575108
rect 338481 575106 338547 575109
rect 312740 575104 338547 575106
rect 312740 575048 338486 575104
rect 338542 575048 338547 575104
rect 312740 575046 338547 575048
rect 312740 575044 312746 575046
rect 338481 575043 338547 575046
rect 409137 575106 409203 575109
rect 442758 575106 442764 575108
rect 409137 575104 442764 575106
rect 409137 575048 409142 575104
rect 409198 575048 442764 575104
rect 409137 575046 442764 575048
rect 409137 575043 409203 575046
rect 442758 575044 442764 575046
rect 442828 575044 442834 575108
rect 448513 575106 448579 575109
rect 448830 575106 448836 575108
rect 448513 575104 448836 575106
rect 448513 575048 448518 575104
rect 448574 575048 448836 575104
rect 448513 575046 448836 575048
rect 448513 575043 448579 575046
rect 448830 575044 448836 575046
rect 448900 575044 448906 575108
rect 280245 574972 280311 574973
rect 280245 574970 280292 574972
rect 280200 574968 280292 574970
rect 280200 574912 280250 574968
rect 280200 574910 280292 574912
rect 280245 574908 280292 574910
rect 280356 574908 280362 574972
rect 281533 574970 281599 574973
rect 282678 574970 282684 574972
rect 281533 574968 282684 574970
rect 281533 574912 281538 574968
rect 281594 574912 282684 574968
rect 281533 574910 282684 574912
rect 280245 574907 280311 574908
rect 281533 574907 281599 574910
rect 282678 574908 282684 574910
rect 282748 574908 282754 574972
rect 287513 574970 287579 574973
rect 288014 574970 288020 574972
rect 287513 574968 288020 574970
rect 287513 574912 287518 574968
rect 287574 574912 288020 574968
rect 287513 574910 288020 574912
rect 287513 574907 287579 574910
rect 288014 574908 288020 574910
rect 288084 574908 288090 574972
rect 290038 574908 290044 574972
rect 290108 574970 290114 574972
rect 291101 574970 291167 574973
rect 290108 574968 291167 574970
rect 290108 574912 291106 574968
rect 291162 574912 291167 574968
rect 290108 574910 291167 574912
rect 290108 574908 290114 574910
rect 291101 574907 291167 574910
rect 310830 574908 310836 574972
rect 310900 574970 310906 574972
rect 341241 574970 341307 574973
rect 310900 574968 341307 574970
rect 310900 574912 341246 574968
rect 341302 574912 341307 574968
rect 310900 574910 341307 574912
rect 310900 574908 310906 574910
rect 341241 574907 341307 574910
rect 409321 574970 409387 574973
rect 431350 574970 431356 574972
rect 409321 574968 431356 574970
rect 409321 574912 409326 574968
rect 409382 574912 431356 574968
rect 409321 574910 431356 574912
rect 409321 574907 409387 574910
rect 431350 574908 431356 574910
rect 431420 574908 431426 574972
rect 284293 574834 284359 574837
rect 284518 574834 284524 574836
rect 284293 574832 284524 574834
rect 284293 574776 284298 574832
rect 284354 574776 284524 574832
rect 284293 574774 284524 574776
rect 284293 574771 284359 574774
rect 284518 574772 284524 574774
rect 284588 574772 284594 574836
rect 288433 574834 288499 574837
rect 291009 574836 291075 574837
rect 288934 574834 288940 574836
rect 288433 574832 288940 574834
rect 288433 574776 288438 574832
rect 288494 574776 288940 574832
rect 288433 574774 288940 574776
rect 288433 574771 288499 574774
rect 288934 574772 288940 574774
rect 289004 574772 289010 574836
rect 290958 574834 290964 574836
rect 290918 574774 290964 574834
rect 291028 574832 291075 574836
rect 291070 574776 291075 574832
rect 290958 574772 290964 574774
rect 291028 574772 291075 574776
rect 291009 574771 291075 574772
rect 292573 574834 292639 574837
rect 292798 574834 292804 574836
rect 292573 574832 292804 574834
rect 292573 574776 292578 574832
rect 292634 574776 292804 574832
rect 292573 574774 292804 574776
rect 292573 574771 292639 574774
rect 292798 574772 292804 574774
rect 292868 574772 292874 574836
rect 310094 574772 310100 574836
rect 310164 574834 310170 574836
rect 341057 574834 341123 574837
rect 310164 574832 341123 574834
rect 310164 574776 341062 574832
rect 341118 574776 341123 574832
rect 310164 574774 341123 574776
rect 310164 574772 310170 574774
rect 341057 574771 341123 574774
rect 408217 574834 408283 574837
rect 432638 574834 432644 574836
rect 408217 574832 432644 574834
rect 408217 574776 408222 574832
rect 408278 574776 432644 574832
rect 408217 574774 432644 574776
rect 408217 574771 408283 574774
rect 432638 574772 432644 574774
rect 432708 574772 432714 574836
rect 438853 574834 438919 574837
rect 439998 574834 440004 574836
rect 438853 574832 440004 574834
rect 438853 574776 438858 574832
rect 438914 574776 440004 574832
rect 438853 574774 440004 574776
rect 438853 574771 438919 574774
rect 439998 574772 440004 574774
rect 440068 574772 440074 574836
rect 444373 574834 444439 574837
rect 445150 574834 445156 574836
rect 444373 574832 445156 574834
rect 444373 574776 444378 574832
rect 444434 574776 445156 574832
rect 444373 574774 445156 574776
rect 444373 574771 444439 574774
rect 445150 574772 445156 574774
rect 445220 574772 445226 574836
rect 198365 574698 198431 574701
rect 307886 574698 307892 574700
rect 198365 574696 307892 574698
rect 198365 574640 198370 574696
rect 198426 574640 307892 574696
rect 198365 574638 307892 574640
rect 198365 574635 198431 574638
rect 307886 574636 307892 574638
rect 307956 574636 307962 574700
rect 308622 574636 308628 574700
rect 308692 574698 308698 574700
rect 341149 574698 341215 574701
rect 308692 574696 341215 574698
rect 308692 574640 341154 574696
rect 341210 574640 341215 574696
rect 308692 574638 341215 574640
rect 308692 574636 308698 574638
rect 341149 574635 341215 574638
rect 451273 574698 451339 574701
rect 452510 574698 452516 574700
rect 451273 574696 452516 574698
rect 451273 574640 451278 574696
rect 451334 574640 452516 574696
rect 451273 574638 452516 574640
rect 451273 574635 451339 574638
rect 452510 574636 452516 574638
rect 452580 574636 452586 574700
rect 288750 574500 288756 574564
rect 288820 574562 288826 574564
rect 289721 574562 289787 574565
rect 288820 574560 289787 574562
rect 288820 574504 289726 574560
rect 289782 574504 289787 574560
rect 288820 574502 289787 574504
rect 288820 574500 288826 574502
rect 289721 574499 289787 574502
rect 296294 574500 296300 574564
rect 296364 574562 296370 574564
rect 296529 574562 296595 574565
rect 296364 574560 296595 574562
rect 296364 574504 296534 574560
rect 296590 574504 296595 574560
rect 296364 574502 296595 574504
rect 296364 574500 296370 574502
rect 296529 574499 296595 574502
rect 298318 574500 298324 574564
rect 298388 574562 298394 574564
rect 298921 574562 298987 574565
rect 298388 574560 298987 574562
rect 298388 574504 298926 574560
rect 298982 574504 298987 574560
rect 298388 574502 298987 574504
rect 298388 574500 298394 574502
rect 298921 574499 298987 574502
rect 299054 574500 299060 574564
rect 299124 574562 299130 574564
rect 299197 574562 299263 574565
rect 299124 574560 299263 574562
rect 299124 574504 299202 574560
rect 299258 574504 299263 574560
rect 299124 574502 299263 574504
rect 299124 574500 299130 574502
rect 299197 574499 299263 574502
rect 299473 574562 299539 574565
rect 300158 574562 300164 574564
rect 299473 574560 300164 574562
rect 299473 574504 299478 574560
rect 299534 574504 300164 574560
rect 299473 574502 300164 574504
rect 299473 574499 299539 574502
rect 300158 574500 300164 574502
rect 300228 574500 300234 574564
rect 451273 574562 451339 574565
rect 451406 574562 451412 574564
rect 451273 574560 451412 574562
rect 451273 574504 451278 574560
rect 451334 574504 451412 574560
rect 451273 574502 451412 574504
rect 451273 574499 451339 574502
rect 451406 574500 451412 574502
rect 451476 574500 451482 574564
rect 455413 574562 455479 574565
rect 456374 574562 456380 574564
rect 455413 574560 456380 574562
rect 455413 574504 455418 574560
rect 455474 574504 456380 574560
rect 455413 574502 456380 574504
rect 455413 574499 455479 574502
rect 456374 574500 456380 574502
rect 456444 574500 456450 574564
rect 463785 574562 463851 574565
rect 463918 574562 463924 574564
rect 463785 574560 463924 574562
rect 463785 574504 463790 574560
rect 463846 574504 463924 574560
rect 463785 574502 463924 574504
rect 463785 574499 463851 574502
rect 463918 574500 463924 574502
rect 463988 574500 463994 574564
rect 253749 574428 253815 574429
rect 253749 574424 253796 574428
rect 253860 574426 253866 574428
rect 273253 574426 273319 574429
rect 274030 574426 274036 574428
rect 253749 574368 253754 574424
rect 253749 574364 253796 574368
rect 253860 574366 253906 574426
rect 273253 574424 274036 574426
rect 273253 574368 273258 574424
rect 273314 574368 274036 574424
rect 273253 574366 274036 574368
rect 253860 574364 253866 574366
rect 253749 574363 253815 574364
rect 273253 574363 273319 574366
rect 274030 574364 274036 574366
rect 274100 574364 274106 574428
rect 276013 574426 276079 574429
rect 293769 574428 293835 574429
rect 294689 574428 294755 574429
rect 276606 574426 276612 574428
rect 276013 574424 276612 574426
rect 276013 574368 276018 574424
rect 276074 574368 276612 574424
rect 276013 574366 276612 574368
rect 276013 574363 276079 574366
rect 276606 574364 276612 574366
rect 276676 574364 276682 574428
rect 293718 574426 293724 574428
rect 293678 574366 293724 574426
rect 293788 574424 293835 574428
rect 294638 574426 294644 574428
rect 293830 574368 293835 574424
rect 293718 574364 293724 574366
rect 293788 574364 293835 574368
rect 294598 574366 294644 574426
rect 294708 574424 294755 574428
rect 294750 574368 294755 574424
rect 294638 574364 294644 574366
rect 294708 574364 294755 574368
rect 293769 574363 293835 574364
rect 294689 574363 294755 574364
rect 433333 574426 433399 574429
rect 458173 574428 458239 574429
rect 433742 574426 433748 574428
rect 433333 574424 433748 574426
rect 433333 574368 433338 574424
rect 433394 574368 433748 574424
rect 433333 574366 433748 574368
rect 433333 574363 433399 574366
rect 433742 574364 433748 574366
rect 433812 574364 433818 574428
rect 458173 574426 458220 574428
rect 458128 574424 458220 574426
rect 458128 574368 458178 574424
rect 458128 574366 458220 574368
rect 458173 574364 458220 574366
rect 458284 574364 458290 574428
rect 459553 574426 459619 574429
rect 465073 574428 465139 574429
rect 492673 574428 492739 574429
rect 460790 574426 460796 574428
rect 459553 574424 460796 574426
rect 459553 574368 459558 574424
rect 459614 574368 460796 574424
rect 459553 574366 460796 574368
rect 458173 574363 458239 574364
rect 459553 574363 459619 574366
rect 460790 574364 460796 574366
rect 460860 574364 460866 574428
rect 465022 574364 465028 574428
rect 465092 574426 465139 574428
rect 465092 574424 465184 574426
rect 465134 574368 465184 574424
rect 465092 574366 465184 574368
rect 465092 574364 465139 574366
rect 492622 574364 492628 574428
rect 492692 574426 492739 574428
rect 492692 574424 492784 574426
rect 492734 574368 492784 574424
rect 492692 574366 492784 574368
rect 492692 574364 492739 574366
rect 465073 574363 465139 574364
rect 492673 574363 492739 574364
rect 252686 574228 252692 574292
rect 252756 574290 252762 574292
rect 254577 574290 254643 574293
rect 252756 574288 254643 574290
rect 252756 574232 254582 574288
rect 254638 574232 254643 574288
rect 252756 574230 254643 574232
rect 252756 574228 252762 574230
rect 254577 574227 254643 574230
rect 269205 574290 269271 574293
rect 270350 574290 270356 574292
rect 269205 574288 270356 574290
rect 269205 574232 269210 574288
rect 269266 574232 270356 574288
rect 269205 574230 270356 574232
rect 269205 574227 269271 574230
rect 270350 574228 270356 574230
rect 270420 574228 270426 574292
rect 274633 574290 274699 574293
rect 278773 574292 278839 574293
rect 275318 574290 275324 574292
rect 274633 574288 275324 574290
rect 274633 574232 274638 574288
rect 274694 574232 275324 574288
rect 274633 574230 275324 574232
rect 274633 574227 274699 574230
rect 275318 574228 275324 574230
rect 275388 574228 275394 574292
rect 278773 574290 278820 574292
rect 278728 574288 278820 574290
rect 278728 574232 278778 574288
rect 278728 574230 278820 574232
rect 278773 574228 278820 574230
rect 278884 574228 278890 574292
rect 285673 574290 285739 574293
rect 286726 574290 286732 574292
rect 285673 574288 286732 574290
rect 285673 574232 285678 574288
rect 285734 574232 286732 574288
rect 285673 574230 286732 574232
rect 278773 574227 278839 574228
rect 285673 574227 285739 574230
rect 286726 574228 286732 574230
rect 286796 574228 286802 574292
rect 298185 574290 298251 574293
rect 298870 574290 298876 574292
rect 298185 574288 298876 574290
rect 298185 574232 298190 574288
rect 298246 574232 298876 574288
rect 298185 574230 298876 574232
rect 298185 574227 298251 574230
rect 298870 574228 298876 574230
rect 298940 574228 298946 574292
rect 303613 574290 303679 574293
rect 303838 574290 303844 574292
rect 303613 574288 303844 574290
rect 303613 574232 303618 574288
rect 303674 574232 303844 574288
rect 303613 574230 303844 574232
rect 303613 574227 303679 574230
rect 303838 574228 303844 574230
rect 303908 574228 303914 574292
rect 313774 574228 313780 574292
rect 313844 574290 313850 574292
rect 337009 574290 337075 574293
rect 313844 574288 337075 574290
rect 313844 574232 337014 574288
rect 337070 574232 337075 574288
rect 313844 574230 337075 574232
rect 313844 574228 313850 574230
rect 337009 574227 337075 574230
rect 436093 574290 436159 574293
rect 436318 574290 436324 574292
rect 436093 574288 436324 574290
rect 436093 574232 436098 574288
rect 436154 574232 436324 574288
rect 436093 574230 436324 574232
rect 436093 574227 436159 574230
rect 436318 574228 436324 574230
rect 436388 574228 436394 574292
rect 440325 574290 440391 574293
rect 440734 574290 440740 574292
rect 440325 574288 440740 574290
rect 440325 574232 440330 574288
rect 440386 574232 440740 574288
rect 440325 574230 440740 574232
rect 440325 574227 440391 574230
rect 440734 574228 440740 574230
rect 440804 574228 440810 574292
rect 443085 574290 443151 574293
rect 444046 574290 444052 574292
rect 443085 574288 444052 574290
rect 443085 574232 443090 574288
rect 443146 574232 444052 574288
rect 443085 574230 444052 574232
rect 443085 574227 443151 574230
rect 444046 574228 444052 574230
rect 444116 574228 444122 574292
rect 444557 574290 444623 574293
rect 445334 574290 445340 574292
rect 444557 574288 445340 574290
rect 444557 574232 444562 574288
rect 444618 574232 445340 574288
rect 444557 574230 445340 574232
rect 444557 574227 444623 574230
rect 445334 574228 445340 574230
rect 445404 574228 445410 574292
rect 445845 574290 445911 574293
rect 446622 574290 446628 574292
rect 445845 574288 446628 574290
rect 445845 574232 445850 574288
rect 445906 574232 446628 574288
rect 445845 574230 446628 574232
rect 445845 574227 445911 574230
rect 446622 574228 446628 574230
rect 446692 574228 446698 574292
rect 447225 574290 447291 574293
rect 447542 574290 447548 574292
rect 447225 574288 447548 574290
rect 447225 574232 447230 574288
rect 447286 574232 447548 574288
rect 447225 574230 447548 574232
rect 447225 574227 447291 574230
rect 447542 574228 447548 574230
rect 447612 574228 447618 574292
rect 449985 574290 450051 574293
rect 452745 574292 452811 574293
rect 450302 574290 450308 574292
rect 449985 574288 450308 574290
rect 449985 574232 449990 574288
rect 450046 574232 450308 574288
rect 449985 574230 450308 574232
rect 449985 574227 450051 574230
rect 450302 574228 450308 574230
rect 450372 574228 450378 574292
rect 452694 574228 452700 574292
rect 452764 574290 452811 574292
rect 454125 574290 454191 574293
rect 454902 574290 454908 574292
rect 452764 574288 452856 574290
rect 452806 574232 452856 574288
rect 452764 574230 452856 574232
rect 454125 574288 454908 574290
rect 454125 574232 454130 574288
rect 454186 574232 454908 574288
rect 454125 574230 454908 574232
rect 452764 574228 452811 574230
rect 452745 574227 452811 574228
rect 454125 574227 454191 574230
rect 454902 574228 454908 574230
rect 454972 574228 454978 574292
rect 456885 574290 456951 574293
rect 457110 574290 457116 574292
rect 456885 574288 457116 574290
rect 456885 574232 456890 574288
rect 456946 574232 457116 574288
rect 456885 574230 457116 574232
rect 456885 574227 456951 574230
rect 457110 574228 457116 574230
rect 457180 574228 457186 574292
rect 461117 574290 461183 574293
rect 461342 574290 461348 574292
rect 461117 574288 461348 574290
rect 461117 574232 461122 574288
rect 461178 574232 461348 574288
rect 461117 574230 461348 574232
rect 461117 574227 461183 574230
rect 461342 574228 461348 574230
rect 461412 574228 461418 574292
rect 464337 574290 464403 574293
rect 465206 574290 465212 574292
rect 464337 574288 465212 574290
rect 464337 574232 464342 574288
rect 464398 574232 465212 574288
rect 464337 574230 465212 574232
rect 464337 574227 464403 574230
rect 465206 574228 465212 574230
rect 465276 574228 465282 574292
rect 470685 574290 470751 574293
rect 471462 574290 471468 574292
rect 470685 574288 471468 574290
rect 470685 574232 470690 574288
rect 470746 574232 471468 574288
rect 470685 574230 471468 574232
rect 470685 574227 470751 574230
rect 471462 574228 471468 574230
rect 471532 574228 471538 574292
rect 492622 574228 492628 574292
rect 492692 574290 492698 574292
rect 492765 574290 492831 574293
rect 492692 574288 492831 574290
rect 492692 574232 492770 574288
rect 492826 574232 492831 574288
rect 492692 574230 492831 574232
rect 492692 574228 492698 574230
rect 492765 574227 492831 574230
rect 252502 574092 252508 574156
rect 252572 574154 252578 574156
rect 253841 574154 253907 574157
rect 269113 574156 269179 574157
rect 252572 574152 253907 574154
rect 252572 574096 253846 574152
rect 253902 574096 253907 574152
rect 252572 574094 253907 574096
rect 252572 574092 252578 574094
rect 253841 574091 253907 574094
rect 269062 574092 269068 574156
rect 269132 574154 269179 574156
rect 270493 574154 270559 574157
rect 271454 574154 271460 574156
rect 269132 574152 269224 574154
rect 269174 574096 269224 574152
rect 269132 574094 269224 574096
rect 270493 574152 271460 574154
rect 270493 574096 270498 574152
rect 270554 574096 271460 574152
rect 270493 574094 271460 574096
rect 269132 574092 269179 574094
rect 269113 574091 269179 574092
rect 270493 574091 270559 574094
rect 271454 574092 271460 574094
rect 271524 574092 271530 574156
rect 271873 574154 271939 574157
rect 272742 574154 272748 574156
rect 271873 574152 272748 574154
rect 271873 574096 271878 574152
rect 271934 574096 272748 574152
rect 271873 574094 272748 574096
rect 271873 574091 271939 574094
rect 272742 574092 272748 574094
rect 272812 574092 272818 574156
rect 277669 574154 277735 574157
rect 278078 574154 278084 574156
rect 277669 574152 278084 574154
rect 277669 574096 277674 574152
rect 277730 574096 278084 574152
rect 277669 574094 278084 574096
rect 277669 574091 277735 574094
rect 278078 574092 278084 574094
rect 278148 574092 278154 574156
rect 278262 574092 278268 574156
rect 278332 574154 278338 574156
rect 278681 574154 278747 574157
rect 278332 574152 278747 574154
rect 278332 574096 278686 574152
rect 278742 574096 278747 574152
rect 278332 574094 278747 574096
rect 278332 574092 278338 574094
rect 278681 574091 278747 574094
rect 278998 574092 279004 574156
rect 279068 574154 279074 574156
rect 280061 574154 280127 574157
rect 279068 574152 280127 574154
rect 279068 574096 280066 574152
rect 280122 574096 280127 574152
rect 279068 574094 280127 574096
rect 279068 574092 279074 574094
rect 280061 574091 280127 574094
rect 280654 574092 280660 574156
rect 280724 574154 280730 574156
rect 281441 574154 281507 574157
rect 280724 574152 281507 574154
rect 280724 574096 281446 574152
rect 281502 574096 281507 574152
rect 280724 574094 281507 574096
rect 280724 574092 280730 574094
rect 281441 574091 281507 574094
rect 282494 574092 282500 574156
rect 282564 574154 282570 574156
rect 282821 574154 282887 574157
rect 282564 574152 282887 574154
rect 282564 574096 282826 574152
rect 282882 574096 282887 574152
rect 282564 574094 282887 574096
rect 282564 574092 282570 574094
rect 282821 574091 282887 574094
rect 283782 574092 283788 574156
rect 283852 574154 283858 574156
rect 284201 574154 284267 574157
rect 283852 574152 284267 574154
rect 283852 574096 284206 574152
rect 284262 574096 284267 574152
rect 283852 574094 284267 574096
rect 283852 574092 283858 574094
rect 284201 574091 284267 574094
rect 295333 574154 295399 574157
rect 298093 574156 298159 574157
rect 296478 574154 296484 574156
rect 295333 574152 296484 574154
rect 295333 574096 295338 574152
rect 295394 574096 296484 574152
rect 295333 574094 296484 574096
rect 295333 574091 295399 574094
rect 296478 574092 296484 574094
rect 296548 574092 296554 574156
rect 298093 574154 298140 574156
rect 298048 574152 298140 574154
rect 298048 574096 298098 574152
rect 298048 574094 298140 574096
rect 298093 574092 298140 574094
rect 298204 574092 298210 574156
rect 300853 574154 300919 574157
rect 301446 574154 301452 574156
rect 300853 574152 301452 574154
rect 300853 574096 300858 574152
rect 300914 574096 301452 574152
rect 300853 574094 301452 574096
rect 298093 574091 298159 574092
rect 300853 574091 300919 574094
rect 301446 574092 301452 574094
rect 301516 574092 301522 574156
rect 302233 574154 302299 574157
rect 302550 574154 302556 574156
rect 302233 574152 302556 574154
rect 302233 574096 302238 574152
rect 302294 574096 302556 574152
rect 302233 574094 302556 574096
rect 302233 574091 302299 574094
rect 302550 574092 302556 574094
rect 302620 574092 302626 574156
rect 304993 574154 305059 574157
rect 305310 574154 305316 574156
rect 304993 574152 305316 574154
rect 304993 574096 304998 574152
rect 305054 574096 305316 574152
rect 304993 574094 305316 574096
rect 304993 574091 305059 574094
rect 305310 574092 305316 574094
rect 305380 574092 305386 574156
rect 306465 574154 306531 574157
rect 306598 574154 306604 574156
rect 306465 574152 306604 574154
rect 306465 574096 306470 574152
rect 306526 574096 306604 574152
rect 306465 574094 306604 574096
rect 306465 574091 306531 574094
rect 306598 574092 306604 574094
rect 306668 574092 306674 574156
rect 318701 574154 318767 574157
rect 318926 574154 318932 574156
rect 318701 574152 318932 574154
rect 318701 574096 318706 574152
rect 318762 574096 318932 574152
rect 318701 574094 318932 574096
rect 318701 574091 318767 574094
rect 318926 574092 318932 574094
rect 318996 574092 319002 574156
rect 336774 574092 336780 574156
rect 336844 574154 336850 574156
rect 337101 574154 337167 574157
rect 336844 574152 337167 574154
rect 336844 574096 337106 574152
rect 337162 574096 337167 574152
rect 336844 574094 337167 574096
rect 336844 574092 336850 574094
rect 337101 574091 337167 574094
rect 434713 574154 434779 574157
rect 434846 574154 434852 574156
rect 434713 574152 434852 574154
rect 434713 574096 434718 574152
rect 434774 574096 434852 574152
rect 434713 574094 434852 574096
rect 434713 574091 434779 574094
rect 434846 574092 434852 574094
rect 434916 574092 434922 574156
rect 436185 574154 436251 574157
rect 437238 574154 437244 574156
rect 436185 574152 437244 574154
rect 436185 574096 436190 574152
rect 436246 574096 437244 574152
rect 436185 574094 437244 574096
rect 436185 574091 436251 574094
rect 437238 574092 437244 574094
rect 437308 574092 437314 574156
rect 437565 574154 437631 574157
rect 437790 574154 437796 574156
rect 437565 574152 437796 574154
rect 437565 574096 437570 574152
rect 437626 574096 437796 574152
rect 437565 574094 437796 574096
rect 437565 574091 437631 574094
rect 437790 574092 437796 574094
rect 437860 574092 437866 574156
rect 438945 574154 439011 574157
rect 439078 574154 439084 574156
rect 438945 574152 439084 574154
rect 438945 574096 438950 574152
rect 439006 574096 439084 574152
rect 438945 574094 439084 574096
rect 438945 574091 439011 574094
rect 439078 574092 439084 574094
rect 439148 574092 439154 574156
rect 440233 574154 440299 574157
rect 440366 574154 440372 574156
rect 440233 574152 440372 574154
rect 440233 574096 440238 574152
rect 440294 574096 440372 574152
rect 440233 574094 440372 574096
rect 440233 574091 440299 574094
rect 440366 574092 440372 574094
rect 440436 574092 440442 574156
rect 441613 574154 441679 574157
rect 442574 574154 442580 574156
rect 441613 574152 442580 574154
rect 441613 574096 441618 574152
rect 441674 574096 442580 574152
rect 441613 574094 442580 574096
rect 441613 574091 441679 574094
rect 442574 574092 442580 574094
rect 442644 574092 442650 574156
rect 442993 574154 443059 574157
rect 444465 574156 444531 574157
rect 443678 574154 443684 574156
rect 442993 574152 443684 574154
rect 442993 574096 442998 574152
rect 443054 574096 443684 574152
rect 442993 574094 443684 574096
rect 442993 574091 443059 574094
rect 443678 574092 443684 574094
rect 443748 574092 443754 574156
rect 444414 574154 444420 574156
rect 444374 574094 444420 574154
rect 444484 574152 444531 574156
rect 444526 574096 444531 574152
rect 444414 574092 444420 574094
rect 444484 574092 444531 574096
rect 444465 574091 444531 574092
rect 445753 574154 445819 574157
rect 446806 574154 446812 574156
rect 445753 574152 446812 574154
rect 445753 574096 445758 574152
rect 445814 574096 446812 574152
rect 445753 574094 446812 574096
rect 445753 574091 445819 574094
rect 446806 574092 446812 574094
rect 446876 574092 446882 574156
rect 447133 574154 447199 574157
rect 447910 574154 447916 574156
rect 447133 574152 447916 574154
rect 447133 574096 447138 574152
rect 447194 574096 447916 574152
rect 447133 574094 447916 574096
rect 447133 574091 447199 574094
rect 447910 574092 447916 574094
rect 447980 574092 447986 574156
rect 448605 574154 448671 574157
rect 449014 574154 449020 574156
rect 448605 574152 449020 574154
rect 448605 574096 448610 574152
rect 448666 574096 449020 574152
rect 448605 574094 449020 574096
rect 448605 574091 448671 574094
rect 449014 574092 449020 574094
rect 449084 574092 449090 574156
rect 449893 574154 449959 574157
rect 450670 574154 450676 574156
rect 449893 574152 450676 574154
rect 449893 574096 449898 574152
rect 449954 574096 450676 574152
rect 449893 574094 450676 574096
rect 449893 574091 449959 574094
rect 450670 574092 450676 574094
rect 450740 574092 450746 574156
rect 451273 574154 451339 574157
rect 451590 574154 451596 574156
rect 451273 574152 451596 574154
rect 451273 574096 451278 574152
rect 451334 574096 451596 574152
rect 451273 574094 451596 574096
rect 451273 574091 451339 574094
rect 451590 574092 451596 574094
rect 451660 574092 451666 574156
rect 452653 574154 452719 574157
rect 453798 574154 453804 574156
rect 452653 574152 453804 574154
rect 452653 574096 452658 574152
rect 452714 574096 453804 574152
rect 452653 574094 453804 574096
rect 452653 574091 452719 574094
rect 453798 574092 453804 574094
rect 453868 574092 453874 574156
rect 454033 574154 454099 574157
rect 454350 574154 454356 574156
rect 454033 574152 454356 574154
rect 454033 574096 454038 574152
rect 454094 574096 454356 574152
rect 454033 574094 454356 574096
rect 454033 574091 454099 574094
rect 454350 574092 454356 574094
rect 454420 574092 454426 574156
rect 455597 574154 455663 574157
rect 456558 574154 456564 574156
rect 455597 574152 456564 574154
rect 455597 574096 455602 574152
rect 455658 574096 456564 574152
rect 455597 574094 456564 574096
rect 455597 574091 455663 574094
rect 456558 574092 456564 574094
rect 456628 574092 456634 574156
rect 456793 574154 456859 574157
rect 457846 574154 457852 574156
rect 456793 574152 457852 574154
rect 456793 574096 456798 574152
rect 456854 574096 457852 574152
rect 456793 574094 457852 574096
rect 456793 574091 456859 574094
rect 457846 574092 457852 574094
rect 457916 574092 457922 574156
rect 458357 574154 458423 574157
rect 458950 574154 458956 574156
rect 458357 574152 458956 574154
rect 458357 574096 458362 574152
rect 458418 574096 458956 574152
rect 458357 574094 458956 574096
rect 458357 574091 458423 574094
rect 458950 574092 458956 574094
rect 459020 574092 459026 574156
rect 459645 574154 459711 574157
rect 460606 574154 460612 574156
rect 459645 574152 460612 574154
rect 459645 574096 459650 574152
rect 459706 574096 460612 574152
rect 459645 574094 460612 574096
rect 459645 574091 459711 574094
rect 460606 574092 460612 574094
rect 460676 574092 460682 574156
rect 461301 574154 461367 574157
rect 461526 574154 461532 574156
rect 461301 574152 461532 574154
rect 461301 574096 461306 574152
rect 461362 574096 461532 574152
rect 461301 574094 461532 574096
rect 461301 574091 461367 574094
rect 461526 574092 461532 574094
rect 461596 574092 461602 574156
rect 462405 574154 462471 574157
rect 462630 574154 462636 574156
rect 462405 574152 462636 574154
rect 462405 574096 462410 574152
rect 462466 574096 462636 574152
rect 462405 574094 462636 574096
rect 462405 574091 462471 574094
rect 462630 574092 462636 574094
rect 462700 574092 462706 574156
rect 463693 574154 463759 574157
rect 466453 574156 466519 574157
rect 464286 574154 464292 574156
rect 463693 574152 464292 574154
rect 463693 574096 463698 574152
rect 463754 574096 464292 574152
rect 463693 574094 464292 574096
rect 463693 574091 463759 574094
rect 464286 574092 464292 574094
rect 464356 574092 464362 574156
rect 466453 574154 466500 574156
rect 466408 574152 466500 574154
rect 466408 574096 466458 574152
rect 466408 574094 466500 574096
rect 466453 574092 466500 574094
rect 466564 574092 466570 574156
rect 466637 574154 466703 574157
rect 467833 574156 467899 574157
rect 470593 574156 470659 574157
rect 466862 574154 466868 574156
rect 466637 574152 466868 574154
rect 466637 574096 466642 574152
rect 466698 574096 466868 574152
rect 466637 574094 466868 574096
rect 466453 574091 466519 574092
rect 466637 574091 466703 574094
rect 466862 574092 466868 574094
rect 466932 574092 466938 574156
rect 467782 574154 467788 574156
rect 467742 574094 467788 574154
rect 467852 574152 467899 574156
rect 467894 574096 467899 574152
rect 467782 574092 467788 574094
rect 467852 574092 467899 574096
rect 470542 574092 470548 574156
rect 470612 574154 470659 574156
rect 471973 574154 472039 574157
rect 472750 574154 472756 574156
rect 470612 574152 470704 574154
rect 470654 574096 470704 574152
rect 470612 574094 470704 574096
rect 471973 574152 472756 574154
rect 471973 574096 471978 574152
rect 472034 574096 472756 574152
rect 471973 574094 472756 574096
rect 470612 574092 470659 574094
rect 467833 574091 467899 574092
rect 470593 574091 470659 574092
rect 471973 574091 472039 574094
rect 472750 574092 472756 574094
rect 472820 574092 472826 574156
rect 473353 574154 473419 574157
rect 474222 574154 474228 574156
rect 473353 574152 474228 574154
rect 473353 574096 473358 574152
rect 473414 574096 474228 574152
rect 473353 574094 474228 574096
rect 473353 574091 473419 574094
rect 474222 574092 474228 574094
rect 474292 574092 474298 574156
rect 474733 574154 474799 574157
rect 475326 574154 475332 574156
rect 474733 574152 475332 574154
rect 474733 574096 474738 574152
rect 474794 574096 475332 574152
rect 474733 574094 475332 574096
rect 474733 574091 474799 574094
rect 475326 574092 475332 574094
rect 475396 574092 475402 574156
rect 476113 574154 476179 574157
rect 476798 574154 476804 574156
rect 476113 574152 476804 574154
rect 476113 574096 476118 574152
rect 476174 574096 476804 574152
rect 476113 574094 476804 574096
rect 476113 574091 476179 574094
rect 476798 574092 476804 574094
rect 476868 574092 476874 574156
rect 405549 572386 405615 572389
rect 433333 572386 433399 572389
rect 405549 572384 433399 572386
rect 405549 572328 405554 572384
rect 405610 572328 433338 572384
rect 433394 572328 433399 572384
rect 405549 572326 433399 572328
rect 405549 572323 405615 572326
rect 433333 572323 433399 572326
rect 405181 572250 405247 572253
rect 434713 572250 434779 572253
rect 405181 572248 434779 572250
rect 405181 572192 405186 572248
rect 405242 572192 434718 572248
rect 434774 572192 434779 572248
rect 405181 572190 434779 572192
rect 405181 572187 405247 572190
rect 434713 572187 434779 572190
rect 405365 572114 405431 572117
rect 436093 572114 436159 572117
rect 405365 572112 436159 572114
rect 405365 572056 405370 572112
rect 405426 572056 436098 572112
rect 436154 572056 436159 572112
rect 405365 572054 436159 572056
rect 405365 572051 405431 572054
rect 436093 572051 436159 572054
rect 3509 571978 3575 571981
rect 407941 571978 408007 571981
rect 3509 571976 408007 571978
rect 3509 571920 3514 571976
rect 3570 571920 407946 571976
rect 408002 571920 408007 571976
rect 3509 571918 408007 571920
rect 3509 571915 3575 571918
rect 407941 571915 408007 571918
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 35709 563140 35775 563141
rect 46749 563140 46815 563141
rect 35709 563136 35756 563140
rect 35820 563138 35826 563140
rect 35709 563080 35714 563136
rect 35709 563076 35756 563080
rect 35820 563078 35866 563138
rect 46749 563136 46796 563140
rect 46860 563138 46866 563140
rect 46749 563080 46754 563136
rect 35820 563076 35826 563078
rect 46749 563076 46796 563080
rect 46860 563078 46906 563138
rect 46860 563076 46866 563078
rect 35709 563075 35775 563076
rect 46749 563075 46815 563076
rect 48037 561780 48103 561781
rect 48037 561776 48094 561780
rect 48158 561778 48164 561780
rect 48037 561720 48042 561776
rect 48037 561716 48094 561720
rect 48158 561718 48194 561778
rect 48158 561716 48164 561718
rect 48037 561715 48103 561716
rect 29318 557160 30032 557220
rect 28809 557154 28875 557157
rect 29318 557154 29378 557160
rect 28809 557152 29378 557154
rect 28809 557096 28814 557152
rect 28870 557096 29378 557152
rect 28809 557094 29378 557096
rect 28809 557091 28875 557094
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect 341609 543148 341675 543149
rect 341558 543084 341564 543148
rect 341628 543146 341675 543148
rect 341628 543144 341720 543146
rect 341670 543088 341720 543144
rect 341628 543086 341720 543088
rect 341628 543084 341675 543086
rect 341609 543083 341675 543084
rect 237281 543010 237347 543013
rect 337142 543010 337148 543012
rect 237281 543008 337148 543010
rect 237281 542952 237286 543008
rect 237342 542952 337148 543008
rect 237281 542950 337148 542952
rect 237281 542947 237347 542950
rect 337142 542948 337148 542950
rect 337212 542948 337218 543012
rect 338982 542948 338988 543012
rect 339052 543010 339058 543012
rect 507853 543010 507919 543013
rect 339052 543008 507919 543010
rect 339052 542952 507858 543008
rect 507914 542952 507919 543008
rect 339052 542950 507919 542952
rect 339052 542948 339058 542950
rect 507853 542947 507919 542950
rect -960 540684 480 540924
rect 527173 540290 527239 540293
rect 528318 540290 528324 540292
rect 527173 540288 528324 540290
rect 527173 540232 527178 540288
rect 527234 540232 528324 540288
rect 527173 540230 528324 540232
rect 527173 540227 527239 540230
rect 528318 540228 528324 540230
rect 528388 540228 528394 540292
rect 198590 539684 198596 539748
rect 198660 539746 198666 539748
rect 216806 539746 216812 539748
rect 198660 539686 216812 539746
rect 198660 539684 198666 539686
rect 216806 539684 216812 539686
rect 216876 539746 216882 539748
rect 217593 539746 217659 539749
rect 216876 539744 217659 539746
rect 216876 539688 217598 539744
rect 217654 539688 217659 539744
rect 216876 539686 217659 539688
rect 216876 539684 216882 539686
rect 217593 539683 217659 539686
rect 528829 539746 528895 539749
rect 529054 539746 529060 539748
rect 528829 539744 529060 539746
rect 528829 539688 528834 539744
rect 528890 539688 529060 539744
rect 528829 539686 529060 539688
rect 528829 539683 528895 539686
rect 529054 539684 529060 539686
rect 529124 539684 529130 539748
rect 218053 539612 218119 539613
rect 218053 539608 218100 539612
rect 218164 539610 218170 539612
rect 218053 539552 218058 539608
rect 218053 539548 218100 539552
rect 218164 539550 218210 539610
rect 218164 539548 218170 539550
rect 218053 539547 218119 539548
rect 205725 539204 205791 539205
rect 205725 539202 205772 539204
rect 205680 539200 205772 539202
rect 205680 539144 205730 539200
rect 205680 539142 205772 539144
rect 205725 539140 205772 539142
rect 205836 539140 205842 539204
rect 205725 539139 205791 539140
rect 540789 538796 540855 538797
rect 540789 538794 540836 538796
rect 540744 538792 540836 538794
rect 540744 538736 540794 538792
rect 540744 538734 540836 538736
rect 540789 538732 540836 538734
rect 540900 538732 540906 538796
rect 540789 538731 540855 538732
rect 578969 537842 579035 537845
rect 583520 537842 584960 537932
rect 578969 537840 584960 537842
rect 578969 537784 578974 537840
rect 579030 537784 584960 537840
rect 578969 537782 584960 537784
rect 578969 537779 579035 537782
rect 583520 537692 584960 537782
rect 197353 533218 197419 533221
rect 199334 533218 200008 533220
rect 197353 533216 200008 533218
rect 197353 533160 197358 533216
rect 197414 533160 200008 533216
rect 546572 533218 547154 533220
rect 549253 533218 549319 533221
rect 546572 533216 549319 533218
rect 546572 533160 549258 533216
rect 549314 533160 549319 533216
rect 197353 533158 199394 533160
rect 547094 533158 549319 533160
rect 197353 533155 197419 533158
rect 549253 533155 549319 533158
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 168373 514994 168439 514997
rect 169017 514994 169083 514997
rect 166766 514992 169083 514994
rect -960 514858 480 514948
rect 166766 514936 168378 514992
rect 168434 514936 169022 514992
rect 169078 514936 169083 514992
rect 166766 514934 169083 514936
rect 166766 514924 166826 514934
rect 168373 514931 168439 514934
rect 169017 514931 169083 514934
rect 166612 514864 166826 514924
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 166612 513912 166826 513972
rect 166766 513906 166826 513912
rect 169109 513906 169175 513909
rect 169569 513906 169635 513909
rect 166766 513904 169635 513906
rect 166766 513848 169114 513904
rect 169170 513848 169574 513904
rect 169630 513848 169635 513904
rect 166766 513846 169635 513848
rect 169109 513843 169175 513846
rect 169569 513843 169635 513846
rect 168649 512002 168715 512005
rect 169293 512002 169359 512005
rect 168649 512000 169359 512002
rect 168649 511944 168654 512000
rect 168710 511944 169298 512000
rect 169354 511944 169359 512000
rect 168649 511942 169359 511944
rect 168649 511939 168715 511942
rect 169293 511939 169359 511942
rect 168465 511866 168531 511869
rect 169201 511866 169267 511869
rect 166766 511864 169267 511866
rect 166766 511808 168470 511864
rect 168526 511808 169206 511864
rect 169262 511808 169267 511864
rect 166766 511806 169267 511808
rect 166766 511796 166826 511806
rect 168465 511803 168531 511806
rect 169201 511803 169267 511806
rect 166612 511736 166826 511796
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 166612 510784 166826 510844
rect 166766 510778 166826 510784
rect 168649 510778 168715 510781
rect 166766 510776 168715 510778
rect 166766 510720 168654 510776
rect 168710 510720 168715 510776
rect 166766 510718 168715 510720
rect 168649 510715 168715 510718
rect 166612 509016 166826 509076
rect 166766 509010 166826 509016
rect 169477 509010 169543 509013
rect 166766 509008 169543 509010
rect 166766 508952 169482 509008
rect 169538 508952 169543 509008
rect 166766 508950 169543 508952
rect 169477 508947 169543 508950
rect 166612 507928 166826 507988
rect 166766 507922 166826 507928
rect 169017 507922 169083 507925
rect 166766 507920 169083 507922
rect 166766 507864 169022 507920
rect 169078 507864 169083 507920
rect 166766 507862 169083 507864
rect 169017 507859 169083 507862
rect 166612 506160 166826 506220
rect 166766 506154 166826 506160
rect 168557 506154 168623 506157
rect 169109 506154 169175 506157
rect 166766 506152 169175 506154
rect 166766 506096 168562 506152
rect 168618 506096 169114 506152
rect 169170 506096 169175 506152
rect 166766 506094 169175 506096
rect 168557 506091 168623 506094
rect 169109 506091 169175 506094
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect 29686 497320 30032 497380
rect 27429 497314 27495 497317
rect 29686 497314 29746 497320
rect 27429 497312 29746 497314
rect 27429 497256 27434 497312
rect 27490 497256 29746 497312
rect 27429 497254 29746 497256
rect 27429 497251 27495 497254
rect 29686 495688 30032 495748
rect 27337 495682 27403 495685
rect 29686 495682 29746 495688
rect 27337 495680 29746 495682
rect 27337 495624 27342 495680
rect 27398 495624 29746 495680
rect 27337 495622 29746 495624
rect 27337 495619 27403 495622
rect 29686 494328 30032 494388
rect 27061 494322 27127 494325
rect 27521 494322 27587 494325
rect 29686 494322 29746 494328
rect 27061 494320 29746 494322
rect 27061 494264 27066 494320
rect 27122 494264 27526 494320
rect 27582 494264 29746 494320
rect 27061 494262 29746 494264
rect 27061 494259 27127 494262
rect 27521 494259 27587 494262
rect 27153 494050 27219 494053
rect 27521 494050 27587 494053
rect 27153 494048 27587 494050
rect 27153 493992 27158 494048
rect 27214 493992 27526 494048
rect 27582 493992 27587 494048
rect 27153 493990 27587 493992
rect 27153 493987 27219 493990
rect 27521 493987 27587 493990
rect 29686 492832 30032 492892
rect 27521 492826 27587 492829
rect 29686 492826 29746 492832
rect 27521 492824 29746 492826
rect 27521 492768 27526 492824
rect 27582 492768 29746 492824
rect 27521 492766 29746 492768
rect 27521 492763 27587 492766
rect 29686 491608 30032 491668
rect 27245 491602 27311 491605
rect 29686 491602 29746 491608
rect 27245 491600 29746 491602
rect 27245 491544 27250 491600
rect 27306 491544 29746 491600
rect 27245 491542 29746 491544
rect 27245 491539 27311 491542
rect 339401 490922 339467 490925
rect 336558 490920 339467 490922
rect 336558 490864 339406 490920
rect 339462 490864 339467 490920
rect 336558 490862 339467 490864
rect 339401 490859 339467 490862
rect 407113 490922 407179 490925
rect 407113 490920 410062 490922
rect 407113 490864 407118 490920
rect 407174 490864 410062 490920
rect 407113 490862 410062 490864
rect 407113 490859 407179 490862
rect 339309 489970 339375 489973
rect 336558 489968 339375 489970
rect 336558 489912 339314 489968
rect 339370 489912 339375 489968
rect 336558 489910 339375 489912
rect 339309 489907 339375 489910
rect 407205 489970 407271 489973
rect 407205 489968 410062 489970
rect 407205 489912 407210 489968
rect 407266 489912 410062 489968
rect 407205 489910 410062 489912
rect 407205 489907 407271 489910
rect -960 488596 480 488836
rect 166612 487936 166826 487996
rect 166766 487930 166826 487936
rect 168925 487930 168991 487933
rect 166766 487928 168991 487930
rect 166766 487872 168930 487928
rect 168986 487872 168991 487928
rect 166766 487870 168991 487872
rect 168925 487867 168991 487870
rect 340045 487794 340111 487797
rect 336558 487792 340111 487794
rect 336558 487736 340050 487792
rect 340106 487736 340111 487792
rect 336558 487734 340111 487736
rect 340045 487731 340111 487734
rect 407113 487794 407179 487797
rect 407113 487792 410062 487794
rect 407113 487736 407118 487792
rect 407174 487736 410062 487792
rect 407113 487734 410062 487736
rect 407113 487731 407179 487734
rect 168925 487250 168991 487253
rect 169385 487250 169451 487253
rect 168925 487248 169451 487250
rect 168925 487192 168930 487248
rect 168986 487192 169390 487248
rect 169446 487192 169451 487248
rect 168925 487190 169451 487192
rect 168925 487187 168991 487190
rect 169385 487187 169451 487190
rect 338849 486842 338915 486845
rect 336558 486840 338915 486842
rect 336558 486784 338854 486840
rect 338910 486784 338915 486840
rect 336558 486782 338915 486784
rect 338849 486779 338915 486782
rect 407113 486842 407179 486845
rect 407113 486840 410062 486842
rect 407113 486784 407118 486840
rect 407174 486784 410062 486840
rect 407113 486782 410062 486784
rect 407113 486779 407179 486782
rect 166612 486304 166826 486364
rect 166766 486298 166826 486304
rect 169661 486298 169727 486301
rect 166766 486296 169727 486298
rect 166766 486240 169666 486296
rect 169722 486240 169727 486296
rect 166766 486238 169727 486240
rect 169661 486235 169727 486238
rect 168833 486162 168899 486165
rect 167134 486160 168899 486162
rect 167134 486104 168838 486160
rect 168894 486104 168899 486160
rect 167134 486102 168899 486104
rect 167134 486092 167194 486102
rect 168833 486099 168899 486102
rect 166612 486032 167194 486092
rect 339401 485074 339467 485077
rect 336558 485072 339467 485074
rect 336558 485016 339406 485072
rect 339462 485016 339467 485072
rect 336558 485014 339467 485016
rect 339401 485011 339467 485014
rect 407113 485074 407179 485077
rect 407113 485072 410062 485074
rect 407113 485016 407118 485072
rect 407174 485016 410062 485072
rect 407113 485014 410062 485016
rect 407113 485011 407179 485014
rect 580625 484666 580691 484669
rect 583520 484666 584960 484756
rect 580625 484664 584960 484666
rect 580625 484608 580630 484664
rect 580686 484608 584960 484664
rect 580625 484606 584960 484608
rect 580625 484603 580691 484606
rect 583520 484516 584960 484606
rect 340045 483986 340111 483989
rect 336558 483984 340111 483986
rect 336558 483928 340050 483984
rect 340106 483928 340111 483984
rect 336558 483926 340111 483928
rect 340045 483923 340111 483926
rect 407113 483986 407179 483989
rect 407113 483984 410062 483986
rect 407113 483928 407118 483984
rect 407174 483928 410062 483984
rect 407113 483926 410062 483928
rect 407113 483923 407179 483926
rect 338849 482218 338915 482221
rect 336558 482216 338915 482218
rect 336558 482160 338854 482216
rect 338910 482160 338915 482216
rect 336558 482158 338915 482160
rect 338849 482155 338915 482158
rect 407113 482218 407179 482221
rect 407113 482216 410062 482218
rect 407113 482160 407118 482216
rect 407174 482160 410062 482216
rect 407113 482158 410062 482160
rect 407113 482155 407179 482158
rect 115473 477868 115539 477869
rect 122649 477868 122715 477869
rect 115408 477804 115414 477868
rect 115478 477866 115539 477868
rect 115478 477864 115570 477866
rect 115534 477808 115570 477864
rect 115478 477806 115570 477808
rect 115478 477804 115539 477806
rect 122616 477804 122622 477868
rect 122686 477866 122715 477868
rect 122686 477864 122778 477866
rect 122710 477808 122778 477864
rect 122686 477806 122778 477808
rect 122686 477804 122715 477806
rect 115473 477803 115539 477804
rect 122649 477803 122715 477804
rect 63166 476172 63172 476236
rect 63236 476172 63242 476236
rect 65742 476172 65748 476236
rect 65812 476172 65818 476236
rect 83038 476172 83044 476236
rect 83108 476172 83114 476236
rect 85614 476172 85620 476236
rect 85684 476172 85690 476236
rect 105670 476172 105676 476236
rect 105740 476172 105746 476236
rect 113030 476172 113036 476236
rect 113100 476172 113106 476236
rect 129590 476172 129596 476236
rect 129660 476172 129666 476236
rect 131982 476172 131988 476236
rect 132052 476172 132058 476236
rect 133086 476172 133092 476236
rect 133156 476172 133162 476236
rect 143390 476172 143396 476236
rect 143460 476172 143466 476236
rect 165429 476234 165495 476237
rect 167126 476234 167132 476236
rect 165429 476232 167132 476234
rect 165429 476176 165434 476232
rect 165490 476176 167132 476232
rect 165429 476174 167132 476176
rect 63174 476098 63234 476172
rect 63401 476098 63467 476101
rect 63174 476096 63467 476098
rect 63174 476040 63406 476096
rect 63462 476040 63467 476096
rect 63174 476038 63467 476040
rect 65750 476098 65810 476172
rect 66161 476098 66227 476101
rect 65750 476096 66227 476098
rect 65750 476040 66166 476096
rect 66222 476040 66227 476096
rect 65750 476038 66227 476040
rect 83046 476098 83106 476172
rect 84101 476098 84167 476101
rect 83046 476096 84167 476098
rect 83046 476040 84106 476096
rect 84162 476040 84167 476096
rect 83046 476038 84167 476040
rect 85622 476098 85682 476172
rect 86861 476098 86927 476101
rect 85622 476096 86927 476098
rect 85622 476040 86866 476096
rect 86922 476040 86927 476096
rect 85622 476038 86927 476040
rect 63401 476035 63467 476038
rect 66161 476035 66227 476038
rect 84101 476035 84167 476038
rect 86861 476035 86927 476038
rect 95366 476036 95372 476100
rect 95436 476098 95442 476100
rect 96521 476098 96587 476101
rect 95436 476096 96587 476098
rect 95436 476040 96526 476096
rect 96582 476040 96587 476096
rect 95436 476038 96587 476040
rect 105678 476098 105738 476172
rect 113038 476101 113098 476172
rect 129598 476101 129658 476172
rect 106181 476098 106247 476101
rect 105678 476096 106247 476098
rect 105678 476040 106186 476096
rect 106242 476040 106247 476096
rect 105678 476038 106247 476040
rect 95436 476036 95442 476038
rect 96521 476035 96587 476038
rect 106181 476035 106247 476038
rect 112989 476096 113098 476101
rect 112989 476040 112994 476096
rect 113050 476040 113098 476096
rect 112989 476038 113098 476040
rect 129549 476096 129658 476101
rect 129549 476040 129554 476096
rect 129610 476040 129658 476096
rect 129549 476038 129658 476040
rect 131990 476098 132050 476172
rect 132401 476098 132467 476101
rect 131990 476096 132467 476098
rect 131990 476040 132406 476096
rect 132462 476040 132467 476096
rect 131990 476038 132467 476040
rect 133094 476098 133154 476172
rect 143398 476101 143458 476172
rect 165429 476171 165495 476174
rect 167126 476172 167132 476174
rect 167196 476172 167202 476236
rect 133781 476098 133847 476101
rect 133094 476096 133847 476098
rect 133094 476040 133786 476096
rect 133842 476040 133847 476096
rect 133094 476038 133847 476040
rect 112989 476035 113055 476038
rect 129549 476035 129615 476038
rect 132401 476035 132467 476038
rect 133781 476035 133847 476038
rect 143349 476096 143458 476101
rect 148317 476100 148383 476101
rect 143349 476040 143354 476096
rect 143410 476040 143458 476096
rect 143349 476038 143458 476040
rect 143349 476035 143415 476038
rect 147070 476036 147076 476100
rect 147140 476098 147146 476100
rect 148317 476098 148364 476100
rect 147140 476096 148364 476098
rect 148428 476098 148434 476100
rect 147140 476040 148322 476096
rect 147140 476038 148364 476040
rect 147140 476036 147146 476038
rect 148317 476036 148364 476038
rect 148428 476038 148474 476098
rect 148428 476036 148434 476038
rect 148317 476035 148383 476036
rect -960 475690 480 475780
rect 122598 475764 122604 475828
rect 122668 475826 122674 475828
rect 124029 475826 124095 475829
rect 122668 475824 124095 475826
rect 122668 475768 124034 475824
rect 124090 475768 124095 475824
rect 122668 475766 124095 475768
rect 122668 475764 122674 475766
rect 124029 475763 124095 475766
rect 141182 475764 141188 475828
rect 141252 475826 141258 475828
rect 141785 475826 141851 475829
rect 141252 475824 141851 475826
rect 141252 475768 141790 475824
rect 141846 475768 141851 475824
rect 141252 475766 141851 475768
rect 141252 475764 141258 475766
rect 141785 475763 141851 475766
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 42793 475556 42859 475557
rect 42742 475492 42748 475556
rect 42812 475554 42859 475556
rect 42812 475552 42904 475554
rect 42854 475496 42904 475552
rect 42812 475494 42904 475496
rect 42812 475492 42859 475494
rect 120206 475492 120212 475556
rect 120276 475554 120282 475556
rect 121177 475554 121243 475557
rect 120276 475552 121243 475554
rect 120276 475496 121182 475552
rect 121238 475496 121243 475552
rect 120276 475494 121243 475496
rect 120276 475492 120282 475494
rect 42793 475491 42859 475492
rect 121177 475491 121243 475494
rect 124806 475492 124812 475556
rect 124876 475554 124882 475556
rect 124876 475494 132510 475554
rect 124876 475492 124882 475494
rect 42793 475418 42859 475421
rect 43662 475418 43668 475420
rect 42793 475416 43668 475418
rect 42793 475360 42798 475416
rect 42854 475360 43668 475416
rect 42793 475358 43668 475360
rect 42793 475355 42859 475358
rect 43662 475356 43668 475358
rect 43732 475356 43738 475420
rect 128486 475356 128492 475420
rect 128556 475418 128562 475420
rect 129641 475418 129707 475421
rect 128556 475416 129707 475418
rect 128556 475360 129646 475416
rect 129702 475360 129707 475416
rect 128556 475358 129707 475360
rect 132450 475418 132510 475494
rect 150566 475492 150572 475556
rect 150636 475554 150642 475556
rect 151353 475554 151419 475557
rect 150636 475552 151419 475554
rect 150636 475496 151358 475552
rect 151414 475496 151419 475552
rect 150636 475494 151419 475496
rect 150636 475492 150642 475494
rect 151353 475491 151419 475494
rect 196382 475418 196388 475420
rect 132450 475358 196388 475418
rect 128556 475356 128562 475358
rect 129641 475355 129707 475358
rect 196382 475356 196388 475358
rect 196452 475356 196458 475420
rect 126278 475220 126284 475284
rect 126348 475282 126354 475284
rect 126881 475282 126947 475285
rect 126348 475280 126947 475282
rect 126348 475224 126886 475280
rect 126942 475224 126947 475280
rect 126348 475222 126947 475224
rect 126348 475220 126354 475222
rect 126881 475219 126947 475222
rect 130694 475220 130700 475284
rect 130764 475282 130770 475284
rect 131021 475282 131087 475285
rect 130764 475280 131087 475282
rect 130764 475224 131026 475280
rect 131082 475224 131087 475280
rect 130764 475222 131087 475224
rect 130764 475220 130770 475222
rect 131021 475219 131087 475222
rect 138238 475220 138244 475284
rect 138308 475282 138314 475284
rect 139301 475282 139367 475285
rect 138308 475280 139367 475282
rect 138308 475224 139306 475280
rect 139362 475224 139367 475280
rect 138308 475222 139367 475224
rect 138308 475220 138314 475222
rect 139301 475219 139367 475222
rect 172421 475282 172487 475285
rect 199510 475282 199516 475284
rect 172421 475280 199516 475282
rect 172421 475224 172426 475280
rect 172482 475224 199516 475280
rect 172421 475222 199516 475224
rect 172421 475219 172487 475222
rect 199510 475220 199516 475222
rect 199580 475220 199586 475284
rect 127198 475084 127204 475148
rect 127268 475146 127274 475148
rect 128261 475146 128327 475149
rect 127268 475144 128327 475146
rect 127268 475088 128266 475144
rect 128322 475088 128327 475144
rect 127268 475086 128327 475088
rect 127268 475084 127274 475086
rect 128261 475083 128327 475086
rect 132718 475084 132724 475148
rect 132788 475146 132794 475148
rect 133689 475146 133755 475149
rect 132788 475144 133755 475146
rect 132788 475088 133694 475144
rect 133750 475088 133755 475144
rect 132788 475086 133755 475088
rect 132788 475084 132794 475086
rect 133689 475083 133755 475086
rect 176653 475146 176719 475149
rect 198038 475146 198044 475148
rect 176653 475144 198044 475146
rect 176653 475088 176658 475144
rect 176714 475088 198044 475144
rect 176653 475086 198044 475088
rect 176653 475083 176719 475086
rect 198038 475084 198044 475086
rect 198108 475084 198114 475148
rect 108062 474948 108068 475012
rect 108132 475010 108138 475012
rect 108849 475010 108915 475013
rect 108132 475008 108915 475010
rect 108132 474952 108854 475008
rect 108910 474952 108915 475008
rect 108132 474950 108915 474952
rect 108132 474948 108138 474950
rect 108849 474947 108915 474950
rect 110086 474948 110092 475012
rect 110156 475010 110162 475012
rect 110321 475010 110387 475013
rect 110156 475008 110387 475010
rect 110156 474952 110326 475008
rect 110382 474952 110387 475008
rect 110156 474950 110387 474952
rect 110156 474948 110162 474950
rect 110321 474947 110387 474950
rect 110454 474948 110460 475012
rect 110524 475010 110530 475012
rect 111609 475010 111675 475013
rect 110524 475008 111675 475010
rect 110524 474952 111614 475008
rect 111670 474952 111675 475008
rect 110524 474950 111675 474952
rect 110524 474948 110530 474950
rect 111609 474947 111675 474950
rect 113766 474948 113772 475012
rect 113836 475010 113842 475012
rect 114369 475010 114435 475013
rect 113836 475008 114435 475010
rect 113836 474952 114374 475008
rect 114430 474952 114435 475008
rect 113836 474950 114435 474952
rect 113836 474948 113842 474950
rect 114369 474947 114435 474950
rect 117814 474948 117820 475012
rect 117884 475010 117890 475012
rect 118601 475010 118667 475013
rect 121361 475012 121427 475013
rect 117884 475008 118667 475010
rect 117884 474952 118606 475008
rect 118662 474952 118667 475008
rect 117884 474950 118667 474952
rect 117884 474948 117890 474950
rect 118601 474947 118667 474950
rect 121310 474948 121316 475012
rect 121380 475010 121427 475012
rect 121380 475008 121472 475010
rect 121422 474952 121472 475008
rect 121380 474950 121472 474952
rect 121380 474948 121427 474950
rect 135294 474948 135300 475012
rect 135364 475010 135370 475012
rect 136449 475010 136515 475013
rect 135364 475008 136515 475010
rect 135364 474952 136454 475008
rect 136510 474952 136515 475008
rect 135364 474950 136515 474952
rect 135364 474948 135370 474950
rect 121361 474947 121427 474948
rect 136449 474947 136515 474950
rect 175273 475010 175339 475013
rect 199326 475010 199332 475012
rect 175273 475008 199332 475010
rect 175273 474952 175278 475008
rect 175334 474952 199332 475008
rect 175273 474950 199332 474952
rect 175273 474947 175339 474950
rect 199326 474948 199332 474950
rect 199396 474948 199402 475012
rect 60641 474876 60707 474877
rect 60590 474812 60596 474876
rect 60660 474874 60707 474876
rect 60660 474872 60752 474874
rect 60702 474816 60752 474872
rect 60660 474814 60752 474816
rect 60660 474812 60707 474814
rect 68134 474812 68140 474876
rect 68204 474874 68210 474876
rect 68921 474874 68987 474877
rect 68204 474872 68987 474874
rect 68204 474816 68926 474872
rect 68982 474816 68987 474872
rect 68204 474814 68987 474816
rect 68204 474812 68210 474814
rect 60641 474811 60707 474812
rect 68921 474811 68987 474814
rect 70710 474812 70716 474876
rect 70780 474874 70786 474876
rect 71681 474874 71747 474877
rect 70780 474872 71747 474874
rect 70780 474816 71686 474872
rect 71742 474816 71747 474872
rect 70780 474814 71747 474816
rect 70780 474812 70786 474814
rect 71681 474811 71747 474814
rect 73654 474812 73660 474876
rect 73724 474874 73730 474876
rect 74441 474874 74507 474877
rect 73724 474872 74507 474874
rect 73724 474816 74446 474872
rect 74502 474816 74507 474872
rect 73724 474814 74507 474816
rect 73724 474812 73730 474814
rect 74441 474811 74507 474814
rect 75310 474812 75316 474876
rect 75380 474874 75386 474876
rect 75821 474874 75887 474877
rect 75380 474872 75887 474874
rect 75380 474816 75826 474872
rect 75882 474816 75887 474872
rect 75380 474814 75887 474816
rect 75380 474812 75386 474814
rect 75821 474811 75887 474814
rect 78070 474812 78076 474876
rect 78140 474874 78146 474876
rect 78581 474874 78647 474877
rect 78140 474872 78647 474874
rect 78140 474816 78586 474872
rect 78642 474816 78647 474872
rect 78140 474814 78647 474816
rect 78140 474812 78146 474814
rect 78581 474811 78647 474814
rect 80646 474812 80652 474876
rect 80716 474874 80722 474876
rect 81341 474874 81407 474877
rect 88241 474876 88307 474877
rect 80716 474872 81407 474874
rect 80716 474816 81346 474872
rect 81402 474816 81407 474872
rect 80716 474814 81407 474816
rect 80716 474812 80722 474814
rect 81341 474811 81407 474814
rect 88190 474812 88196 474876
rect 88260 474874 88307 474876
rect 88260 474872 88352 474874
rect 88302 474816 88352 474872
rect 88260 474814 88352 474816
rect 88260 474812 88307 474814
rect 90766 474812 90772 474876
rect 90836 474874 90842 474876
rect 91001 474874 91067 474877
rect 93761 474876 93827 474877
rect 93710 474874 93716 474876
rect 90836 474872 91067 474874
rect 90836 474816 91006 474872
rect 91062 474816 91067 474872
rect 90836 474814 91067 474816
rect 93670 474814 93716 474874
rect 93780 474872 93827 474876
rect 93822 474816 93827 474872
rect 90836 474812 90842 474814
rect 88241 474811 88307 474812
rect 91001 474811 91067 474814
rect 93710 474812 93716 474814
rect 93780 474812 93827 474816
rect 98310 474812 98316 474876
rect 98380 474874 98386 474876
rect 99281 474874 99347 474877
rect 98380 474872 99347 474874
rect 98380 474816 99286 474872
rect 99342 474816 99347 474872
rect 98380 474814 99347 474816
rect 98380 474812 98386 474814
rect 93761 474811 93827 474812
rect 99281 474811 99347 474814
rect 100518 474812 100524 474876
rect 100588 474874 100594 474876
rect 100661 474874 100727 474877
rect 100588 474872 100727 474874
rect 100588 474816 100666 474872
rect 100722 474816 100727 474872
rect 100588 474814 100727 474816
rect 100588 474812 100594 474814
rect 100661 474811 100727 474814
rect 102726 474812 102732 474876
rect 102796 474874 102802 474876
rect 103421 474874 103487 474877
rect 102796 474872 103487 474874
rect 102796 474816 103426 474872
rect 103482 474816 103487 474872
rect 102796 474814 103487 474816
rect 102796 474812 102802 474814
rect 103421 474811 103487 474814
rect 107326 474812 107332 474876
rect 107396 474874 107402 474876
rect 107561 474874 107627 474877
rect 107396 474872 107627 474874
rect 107396 474816 107566 474872
rect 107622 474816 107627 474872
rect 107396 474814 107627 474816
rect 107396 474812 107402 474814
rect 107561 474811 107627 474814
rect 108430 474812 108436 474876
rect 108500 474874 108506 474876
rect 108941 474874 109007 474877
rect 108500 474872 109007 474874
rect 108500 474816 108946 474872
rect 109002 474816 109007 474872
rect 108500 474814 109007 474816
rect 108500 474812 108506 474814
rect 108941 474811 109007 474814
rect 110822 474812 110828 474876
rect 110892 474874 110898 474876
rect 111701 474874 111767 474877
rect 110892 474872 111767 474874
rect 110892 474816 111706 474872
rect 111762 474816 111767 474872
rect 110892 474814 111767 474816
rect 110892 474812 110898 474814
rect 111701 474811 111767 474814
rect 112662 474812 112668 474876
rect 112732 474874 112738 474876
rect 113081 474874 113147 474877
rect 112732 474872 113147 474874
rect 112732 474816 113086 474872
rect 113142 474816 113147 474872
rect 112732 474814 113147 474816
rect 112732 474812 112738 474814
rect 113081 474811 113147 474814
rect 114318 474812 114324 474876
rect 114388 474874 114394 474876
rect 114461 474874 114527 474877
rect 114388 474872 114527 474874
rect 114388 474816 114466 474872
rect 114522 474816 114527 474872
rect 114388 474814 114527 474816
rect 114388 474812 114394 474814
rect 114461 474811 114527 474814
rect 115238 474812 115244 474876
rect 115308 474874 115314 474876
rect 115749 474874 115815 474877
rect 115308 474872 115815 474874
rect 115308 474816 115754 474872
rect 115810 474816 115815 474872
rect 115308 474814 115815 474816
rect 115308 474812 115314 474814
rect 115749 474811 115815 474814
rect 116710 474812 116716 474876
rect 116780 474874 116786 474876
rect 117221 474874 117287 474877
rect 116780 474872 117287 474874
rect 116780 474816 117226 474872
rect 117282 474816 117287 474872
rect 116780 474814 117287 474816
rect 116780 474812 116786 474814
rect 117221 474811 117287 474814
rect 118366 474812 118372 474876
rect 118436 474874 118442 474876
rect 118509 474874 118575 474877
rect 118436 474872 118575 474874
rect 118436 474816 118514 474872
rect 118570 474816 118575 474872
rect 118436 474814 118575 474816
rect 118436 474812 118442 474814
rect 118509 474811 118575 474814
rect 118918 474812 118924 474876
rect 118988 474874 118994 474876
rect 119981 474874 120047 474877
rect 118988 474872 120047 474874
rect 118988 474816 119986 474872
rect 120042 474816 120047 474872
rect 118988 474814 120047 474816
rect 118988 474812 118994 474814
rect 119981 474811 120047 474814
rect 120574 474812 120580 474876
rect 120644 474874 120650 474876
rect 121269 474874 121335 474877
rect 120644 474872 121335 474874
rect 120644 474816 121274 474872
rect 121330 474816 121335 474872
rect 120644 474814 121335 474816
rect 120644 474812 120650 474814
rect 121269 474811 121335 474814
rect 123702 474812 123708 474876
rect 123772 474874 123778 474876
rect 124121 474874 124187 474877
rect 123772 474872 124187 474874
rect 123772 474816 124126 474872
rect 124182 474816 124187 474872
rect 123772 474814 124187 474816
rect 123772 474812 123778 474814
rect 124121 474811 124187 474814
rect 125358 474812 125364 474876
rect 125428 474874 125434 474876
rect 125501 474874 125567 474877
rect 125428 474872 125567 474874
rect 125428 474816 125506 474872
rect 125562 474816 125567 474872
rect 125428 474814 125567 474816
rect 125428 474812 125434 474814
rect 125501 474811 125567 474814
rect 128118 474812 128124 474876
rect 128188 474874 128194 474876
rect 128261 474874 128327 474877
rect 128188 474872 128327 474874
rect 128188 474816 128266 474872
rect 128322 474816 128327 474872
rect 128188 474814 128327 474816
rect 128188 474812 128194 474814
rect 128261 474811 128327 474814
rect 130510 474812 130516 474876
rect 130580 474874 130586 474876
rect 131021 474874 131087 474877
rect 130580 474872 131087 474874
rect 130580 474816 131026 474872
rect 131082 474816 131087 474872
rect 130580 474814 131087 474816
rect 130580 474812 130586 474814
rect 131021 474811 131087 474814
rect 134190 474812 134196 474876
rect 134260 474874 134266 474876
rect 135161 474874 135227 474877
rect 134260 474872 135227 474874
rect 134260 474816 135166 474872
rect 135222 474816 135227 474872
rect 134260 474814 135227 474816
rect 134260 474812 134266 474814
rect 135161 474811 135227 474814
rect 136214 474812 136220 474876
rect 136284 474874 136290 474876
rect 136357 474874 136423 474877
rect 136541 474876 136607 474877
rect 137921 474876 137987 474877
rect 136541 474874 136588 474876
rect 136284 474872 136423 474874
rect 136284 474816 136362 474872
rect 136418 474816 136423 474872
rect 136284 474814 136423 474816
rect 136496 474872 136588 474874
rect 136496 474816 136546 474872
rect 136496 474814 136588 474816
rect 136284 474812 136290 474814
rect 136357 474811 136423 474814
rect 136541 474812 136588 474814
rect 136652 474812 136658 474876
rect 137870 474812 137876 474876
rect 137940 474874 137987 474876
rect 137940 474872 138032 474874
rect 137982 474816 138032 474872
rect 137940 474814 138032 474816
rect 137940 474812 137987 474814
rect 138974 474812 138980 474876
rect 139044 474874 139050 474876
rect 139209 474874 139275 474877
rect 139044 474872 139275 474874
rect 139044 474816 139214 474872
rect 139270 474816 139275 474872
rect 139044 474814 139275 474816
rect 139044 474812 139050 474814
rect 136541 474811 136607 474812
rect 137921 474811 137987 474812
rect 139209 474811 139275 474814
rect 140078 474812 140084 474876
rect 140148 474874 140154 474876
rect 140681 474874 140747 474877
rect 140148 474872 140747 474874
rect 140148 474816 140686 474872
rect 140742 474816 140747 474872
rect 140148 474814 140747 474816
rect 140148 474812 140154 474814
rect 140681 474811 140747 474814
rect 142654 474812 142660 474876
rect 142724 474874 142730 474876
rect 143441 474874 143507 474877
rect 142724 474872 143507 474874
rect 142724 474816 143446 474872
rect 143502 474816 143507 474872
rect 142724 474814 143507 474816
rect 142724 474812 142730 474814
rect 143441 474811 143507 474814
rect 150014 474812 150020 474876
rect 150084 474874 150090 474876
rect 150341 474874 150407 474877
rect 150084 474872 150407 474874
rect 150084 474816 150346 474872
rect 150402 474816 150407 474872
rect 150084 474814 150407 474816
rect 150084 474812 150090 474814
rect 150341 474811 150407 474814
rect 187693 474874 187759 474877
rect 197854 474874 197860 474876
rect 187693 474872 197860 474874
rect 187693 474816 187698 474872
rect 187754 474816 197860 474872
rect 187693 474814 197860 474816
rect 187693 474811 187759 474814
rect 197854 474812 197860 474814
rect 197924 474812 197930 474876
rect 198273 473378 198339 473381
rect 199334 473378 200008 473380
rect 198273 473376 200008 473378
rect 198273 473320 198278 473376
rect 198334 473320 200008 473376
rect 546572 473378 547154 473380
rect 549345 473378 549411 473381
rect 546572 473376 549411 473378
rect 546572 473320 549350 473376
rect 549406 473320 549411 473376
rect 198273 473318 199394 473320
rect 547094 473318 549411 473320
rect 198273 473315 198339 473318
rect 549345 473315 549411 473318
rect 198181 471746 198247 471749
rect 199334 471746 200008 471748
rect 198181 471744 200008 471746
rect 198181 471688 198186 471744
rect 198242 471688 200008 471744
rect 546572 471746 547154 471748
rect 549437 471746 549503 471749
rect 546572 471744 549503 471746
rect 546572 471688 549442 471744
rect 549498 471688 549503 471744
rect 198181 471686 199394 471688
rect 547094 471686 549503 471688
rect 198181 471683 198247 471686
rect 549437 471683 549503 471686
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect 198089 470386 198155 470389
rect 199334 470386 200008 470388
rect 198089 470384 200008 470386
rect 198089 470328 198094 470384
rect 198150 470328 200008 470384
rect 546572 470386 547154 470388
rect 549529 470386 549595 470389
rect 546572 470384 549595 470386
rect 546572 470328 549534 470384
rect 549590 470328 549595 470384
rect 198089 470326 199394 470328
rect 547094 470326 549595 470328
rect 198089 470323 198155 470326
rect 549529 470323 549595 470326
rect 197997 468890 198063 468893
rect 199334 468890 200008 468892
rect 197997 468888 200008 468890
rect 197997 468832 198002 468888
rect 198058 468832 200008 468888
rect 546572 468890 547154 468892
rect 549621 468890 549687 468893
rect 546572 468888 549687 468890
rect 546572 468832 549626 468888
rect 549682 468832 549687 468888
rect 197997 468830 199394 468832
rect 547094 468830 549687 468832
rect 197997 468827 198063 468830
rect 549621 468827 549687 468830
rect 197813 467666 197879 467669
rect 199334 467666 200008 467668
rect 197813 467664 200008 467666
rect 197813 467608 197818 467664
rect 197874 467608 200008 467664
rect 546572 467666 547154 467668
rect 549713 467666 549779 467669
rect 546572 467664 549779 467666
rect 546572 467608 549718 467664
rect 549774 467608 549779 467664
rect 197813 467606 199394 467608
rect 547094 467606 549779 467608
rect 197813 467603 197879 467606
rect 549713 467603 549779 467606
rect 339401 463994 339467 463997
rect 336558 463992 339467 463994
rect 336558 463936 339406 463992
rect 339462 463936 339467 463992
rect 336558 463934 339467 463936
rect 339401 463931 339467 463934
rect 407113 463994 407179 463997
rect 407113 463992 410062 463994
rect 407113 463936 407118 463992
rect 407174 463936 410062 463992
rect 407113 463934 410062 463936
rect 407113 463931 407179 463934
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 336588 462362 337210 462364
rect 339125 462362 339191 462365
rect 336588 462360 339191 462362
rect 336588 462304 339130 462360
rect 339186 462304 339191 462360
rect 337150 462302 339191 462304
rect 339125 462299 339191 462302
rect 407113 462362 407179 462365
rect 409462 462362 410032 462364
rect 407113 462360 410032 462362
rect 407113 462304 407118 462360
rect 407174 462304 410032 462360
rect 407113 462302 409522 462304
rect 407113 462299 407179 462302
rect 338430 462090 338436 462092
rect 336558 462030 338436 462090
rect 338430 462028 338436 462030
rect 338500 462028 338506 462092
rect 407113 462090 407179 462093
rect 407113 462088 410062 462090
rect 407113 462032 407118 462088
rect 407174 462032 410062 462088
rect 407113 462030 410062 462032
rect 407113 462027 407179 462030
rect 338430 461484 338436 461548
rect 338500 461546 338506 461548
rect 339033 461546 339099 461549
rect 338500 461544 339099 461546
rect 338500 461488 339038 461544
rect 339094 461488 339099 461544
rect 338500 461486 339099 461488
rect 338500 461484 338506 461486
rect 339033 461483 339099 461486
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 107561 456242 107627 456245
rect 168557 456242 168623 456245
rect 107561 456240 168623 456242
rect 107561 456184 107566 456240
rect 107622 456184 168562 456240
rect 168618 456184 168623 456240
rect 107561 456182 168623 456184
rect 107561 456179 107627 456182
rect 168557 456179 168623 456182
rect 111701 456106 111767 456109
rect 111701 456104 161490 456106
rect 111701 456048 111706 456104
rect 111762 456048 161490 456104
rect 111701 456046 161490 456048
rect 111701 456043 111767 456046
rect 161430 455698 161490 456046
rect 168741 455834 168807 455837
rect 168966 455834 168972 455836
rect 168741 455832 168972 455834
rect 168741 455776 168746 455832
rect 168802 455776 168972 455832
rect 168741 455774 168972 455776
rect 168741 455771 168807 455774
rect 168966 455772 168972 455774
rect 169036 455772 169042 455836
rect 173065 455698 173131 455701
rect 198958 455698 198964 455700
rect 161430 455696 198964 455698
rect 161430 455640 173070 455696
rect 173126 455640 198964 455696
rect 161430 455638 198964 455640
rect 173065 455635 173131 455638
rect 198958 455636 198964 455638
rect 199028 455636 199034 455700
rect 168557 455562 168623 455565
rect 169201 455562 169267 455565
rect 197302 455562 197308 455564
rect 168557 455560 197308 455562
rect 168557 455504 168562 455560
rect 168618 455504 169206 455560
rect 169262 455504 197308 455560
rect 168557 455502 197308 455504
rect 168557 455499 168623 455502
rect 169201 455499 169267 455502
rect 197302 455500 197308 455502
rect 197372 455500 197378 455564
rect 108941 454746 109007 454749
rect 169845 454746 169911 454749
rect 108941 454744 169911 454746
rect 108941 454688 108946 454744
rect 109002 454688 169850 454744
rect 169906 454688 169911 454744
rect 108941 454686 169911 454688
rect 108941 454683 109007 454686
rect 169845 454683 169911 454686
rect 169845 454066 169911 454069
rect 170581 454066 170647 454069
rect 198774 454066 198780 454068
rect 169845 454064 198780 454066
rect 169845 454008 169850 454064
rect 169906 454008 170586 454064
rect 170642 454008 198780 454064
rect 169845 454006 198780 454008
rect 169845 454003 169911 454006
rect 170581 454003 170647 454006
rect 198774 454004 198780 454006
rect 198844 454004 198850 454068
rect 288893 453796 288959 453797
rect 294781 453796 294847 453797
rect 288893 453792 288950 453796
rect 289014 453794 289020 453796
rect 288893 453736 288898 453792
rect 288893 453732 288950 453736
rect 289014 453734 289050 453794
rect 294781 453792 294798 453796
rect 294862 453794 294868 453796
rect 294781 453736 294786 453792
rect 289014 453732 289020 453734
rect 294781 453732 294798 453736
rect 294862 453734 294938 453794
rect 294862 453732 294868 453734
rect 429584 453732 429590 453796
rect 429654 453794 429660 453796
rect 430536 453794 430542 453796
rect 429654 453734 430542 453794
rect 429654 453732 429660 453734
rect 430536 453732 430542 453734
rect 430606 453794 430612 453796
rect 431760 453794 431766 453796
rect 430606 453734 431766 453794
rect 430606 453732 430612 453734
rect 431760 453732 431766 453734
rect 431830 453732 431836 453796
rect 288893 453731 288959 453732
rect 294781 453731 294847 453732
rect 213177 453658 213243 453661
rect 284293 453660 284359 453661
rect 286777 453660 286843 453661
rect 290181 453660 290247 453661
rect 213328 453658 213334 453660
rect 213177 453656 213334 453658
rect 213177 453600 213182 453656
rect 213238 453600 213334 453656
rect 213177 453598 213334 453600
rect 213177 453595 213243 453598
rect 213328 453596 213334 453598
rect 213398 453596 213404 453660
rect 284293 453656 284326 453660
rect 284390 453658 284396 453660
rect 286768 453658 286774 453660
rect 284293 453600 284298 453656
rect 284293 453596 284326 453600
rect 284390 453598 284450 453658
rect 286686 453598 286774 453658
rect 284390 453596 284396 453598
rect 286768 453596 286774 453598
rect 286838 453596 286844 453660
rect 290168 453658 290174 453660
rect 290090 453598 290174 453658
rect 290238 453656 290247 453660
rect 290242 453600 290247 453656
rect 290168 453596 290174 453598
rect 290238 453596 290247 453600
rect 284293 453595 284359 453596
rect 286777 453595 286843 453596
rect 290181 453595 290247 453596
rect 291193 453660 291259 453661
rect 293677 453660 293743 453661
rect 297081 453660 297147 453661
rect 298461 453660 298527 453661
rect 299565 453660 299631 453661
rect 291193 453656 291262 453660
rect 291193 453600 291198 453656
rect 291254 453600 291262 453656
rect 291193 453596 291262 453600
rect 291326 453658 291332 453660
rect 291326 453598 291350 453658
rect 293677 453656 293710 453660
rect 293774 453658 293780 453660
rect 293677 453600 293682 453656
rect 291326 453596 291332 453598
rect 293677 453596 293710 453600
rect 293774 453598 293834 453658
rect 297081 453656 297110 453660
rect 297174 453658 297180 453660
rect 297081 453600 297086 453656
rect 293774 453596 293780 453598
rect 297081 453596 297110 453600
rect 297174 453598 297238 453658
rect 298461 453656 298470 453660
rect 298534 453658 298540 453660
rect 299552 453658 299558 453660
rect 298461 453600 298466 453656
rect 297174 453596 297180 453598
rect 298461 453596 298470 453600
rect 298534 453598 298618 453658
rect 299474 453598 299558 453658
rect 299622 453656 299631 453660
rect 299626 453600 299631 453656
rect 298534 453596 298540 453598
rect 299552 453596 299558 453598
rect 299622 453596 299631 453600
rect 291193 453595 291259 453596
rect 293677 453595 293743 453596
rect 297081 453595 297147 453596
rect 298461 453595 298527 453596
rect 299565 453595 299631 453596
rect 311065 453660 311131 453661
rect 312353 453660 312419 453661
rect 443637 453660 443703 453661
rect 311065 453656 311118 453660
rect 311182 453658 311188 453660
rect 312336 453658 312342 453660
rect 311065 453600 311070 453656
rect 311065 453596 311118 453600
rect 311182 453598 311222 453658
rect 312262 453598 312342 453658
rect 312406 453656 312419 453660
rect 443592 453658 443598 453660
rect 312414 453600 312419 453656
rect 311182 453596 311188 453598
rect 312336 453596 312342 453598
rect 312406 453596 312419 453600
rect 443546 453598 443598 453658
rect 443662 453656 443703 453660
rect 443698 453600 443703 453656
rect 443592 453596 443598 453598
rect 443662 453596 443703 453600
rect 532734 453596 532740 453660
rect 532804 453658 532810 453660
rect 533216 453658 533222 453660
rect 532804 453598 533222 453658
rect 532804 453596 532810 453598
rect 533216 453596 533222 453598
rect 533286 453596 533292 453660
rect 311065 453595 311131 453596
rect 312353 453595 312419 453596
rect 443637 453595 443703 453596
rect 178861 453250 178927 453253
rect 196157 453250 196223 453253
rect 196382 453250 196388 453252
rect 178861 453248 196388 453250
rect 178861 453192 178866 453248
rect 178922 453192 196162 453248
rect 196218 453192 196388 453248
rect 178861 453190 196388 453192
rect 178861 453187 178927 453190
rect 196157 453187 196223 453190
rect 196382 453188 196388 453190
rect 196452 453188 196458 453252
rect 199510 453052 199516 453116
rect 199580 453114 199586 453116
rect 279550 453114 279556 453116
rect 199580 453054 279556 453114
rect 199580 453052 199586 453054
rect 279550 453052 279556 453054
rect 279620 453052 279626 453116
rect 199326 452916 199332 452980
rect 199396 452978 199402 452980
rect 285254 452978 285260 452980
rect 199396 452918 285260 452978
rect 199396 452916 199402 452918
rect 285254 452916 285260 452918
rect 285324 452916 285330 452980
rect 198038 452780 198044 452844
rect 198108 452842 198114 452844
rect 295926 452842 295932 452844
rect 198108 452782 295932 452842
rect 198108 452780 198114 452782
rect 295926 452780 295932 452782
rect 295996 452780 296002 452844
rect 197854 452644 197860 452708
rect 197924 452706 197930 452708
rect 297081 452706 297147 452709
rect 197924 452704 297147 452706
rect 197924 452648 297086 452704
rect 297142 452648 297147 452704
rect 197924 452646 297147 452648
rect 197924 452644 197930 452646
rect 297081 452643 297147 452646
rect 34513 452570 34579 452573
rect 35198 452570 35204 452572
rect 34513 452568 35204 452570
rect 34513 452512 34518 452568
rect 34574 452512 35204 452568
rect 34513 452510 35204 452512
rect 34513 452507 34579 452510
rect 35198 452508 35204 452510
rect 35268 452508 35274 452572
rect 230606 452508 230612 452572
rect 230676 452570 230682 452572
rect 231761 452570 231827 452573
rect 230676 452568 231827 452570
rect 230676 452512 231766 452568
rect 231822 452512 231827 452568
rect 230676 452510 231827 452512
rect 230676 452508 230682 452510
rect 231761 452507 231827 452510
rect 233182 452508 233188 452572
rect 233252 452570 233258 452572
rect 234521 452570 234587 452573
rect 233252 452568 234587 452570
rect 233252 452512 234526 452568
rect 234582 452512 234587 452568
rect 233252 452510 234587 452512
rect 233252 452508 233258 452510
rect 234521 452507 234587 452510
rect 235574 452508 235580 452572
rect 235644 452570 235650 452572
rect 235901 452570 235967 452573
rect 235644 452568 235967 452570
rect 235644 452512 235906 452568
rect 235962 452512 235967 452568
rect 235644 452510 235967 452512
rect 235644 452508 235650 452510
rect 235901 452507 235967 452510
rect 238150 452508 238156 452572
rect 238220 452570 238226 452572
rect 238661 452570 238727 452573
rect 238220 452568 238727 452570
rect 238220 452512 238666 452568
rect 238722 452512 238727 452568
rect 238220 452510 238727 452512
rect 238220 452508 238226 452510
rect 238661 452507 238727 452510
rect 240726 452508 240732 452572
rect 240796 452570 240802 452572
rect 241421 452570 241487 452573
rect 243169 452572 243235 452573
rect 245561 452572 245627 452573
rect 243118 452570 243124 452572
rect 240796 452568 241487 452570
rect 240796 452512 241426 452568
rect 241482 452512 241487 452568
rect 240796 452510 241487 452512
rect 243078 452510 243124 452570
rect 243188 452568 243235 452572
rect 245510 452570 245516 452572
rect 243230 452512 243235 452568
rect 240796 452508 240802 452510
rect 241421 452507 241487 452510
rect 243118 452508 243124 452510
rect 243188 452508 243235 452512
rect 245470 452510 245516 452570
rect 245580 452568 245627 452572
rect 245622 452512 245627 452568
rect 245510 452508 245516 452510
rect 245580 452508 245627 452512
rect 253054 452508 253060 452572
rect 253124 452570 253130 452572
rect 253841 452570 253907 452573
rect 255681 452572 255747 452573
rect 255630 452570 255636 452572
rect 253124 452568 253907 452570
rect 253124 452512 253846 452568
rect 253902 452512 253907 452568
rect 253124 452510 253907 452512
rect 255590 452510 255636 452570
rect 255700 452568 255747 452572
rect 255742 452512 255747 452568
rect 253124 452508 253130 452510
rect 243169 452507 243235 452508
rect 245561 452507 245627 452508
rect 253841 452507 253907 452510
rect 255630 452508 255636 452510
rect 255700 452508 255747 452512
rect 260598 452508 260604 452572
rect 260668 452570 260674 452572
rect 260741 452570 260807 452573
rect 260668 452568 260807 452570
rect 260668 452512 260746 452568
rect 260802 452512 260807 452568
rect 260668 452510 260807 452512
rect 260668 452508 260674 452510
rect 255681 452507 255747 452508
rect 260741 452507 260807 452510
rect 263174 452508 263180 452572
rect 263244 452570 263250 452572
rect 263501 452570 263567 452573
rect 265617 452572 265683 452573
rect 265566 452570 265572 452572
rect 263244 452568 263567 452570
rect 263244 452512 263506 452568
rect 263562 452512 263567 452568
rect 263244 452510 263567 452512
rect 265526 452510 265572 452570
rect 265636 452568 265683 452572
rect 265678 452512 265683 452568
rect 263244 452508 263250 452510
rect 263501 452507 263567 452510
rect 265566 452508 265572 452510
rect 265636 452508 265683 452512
rect 268326 452508 268332 452572
rect 268396 452570 268402 452572
rect 269021 452570 269087 452573
rect 268396 452568 269087 452570
rect 268396 452512 269026 452568
rect 269082 452512 269087 452568
rect 268396 452510 269087 452512
rect 268396 452508 268402 452510
rect 265617 452507 265683 452508
rect 269021 452507 269087 452510
rect 270534 452508 270540 452572
rect 270604 452570 270610 452572
rect 271781 452570 271847 452573
rect 273161 452572 273227 452573
rect 273110 452570 273116 452572
rect 270604 452568 271847 452570
rect 270604 452512 271786 452568
rect 271842 452512 271847 452568
rect 270604 452510 271847 452512
rect 273070 452510 273116 452570
rect 273180 452568 273227 452572
rect 273222 452512 273227 452568
rect 270604 452508 270610 452510
rect 271781 452507 271847 452510
rect 273110 452508 273116 452510
rect 273180 452508 273227 452512
rect 275686 452508 275692 452572
rect 275756 452570 275762 452572
rect 275829 452570 275895 452573
rect 275756 452568 275895 452570
rect 275756 452512 275834 452568
rect 275890 452512 275895 452568
rect 275756 452510 275895 452512
rect 275756 452508 275762 452510
rect 273161 452507 273227 452508
rect 275829 452507 275895 452510
rect 278078 452508 278084 452572
rect 278148 452570 278154 452572
rect 278681 452570 278747 452573
rect 278148 452568 278747 452570
rect 278148 452512 278686 452568
rect 278742 452512 278747 452568
rect 278148 452510 278747 452512
rect 278148 452508 278154 452510
rect 278681 452507 278747 452510
rect 280153 452570 280219 452573
rect 282085 452572 282151 452573
rect 280470 452570 280476 452572
rect 280153 452568 280476 452570
rect 280153 452512 280158 452568
rect 280214 452512 280476 452568
rect 280153 452510 280476 452512
rect 280153 452507 280219 452510
rect 280470 452508 280476 452510
rect 280540 452508 280546 452572
rect 282085 452568 282132 452572
rect 282196 452570 282202 452572
rect 282085 452512 282090 452568
rect 282085 452508 282132 452512
rect 282196 452510 282242 452570
rect 282196 452508 282202 452510
rect 283046 452508 283052 452572
rect 283116 452570 283122 452572
rect 284201 452570 284267 452573
rect 283116 452568 284267 452570
rect 283116 452512 284206 452568
rect 284262 452512 284267 452568
rect 283116 452510 284267 452512
rect 283116 452508 283122 452510
rect 282085 452507 282151 452508
rect 284201 452507 284267 452510
rect 285581 452572 285647 452573
rect 285581 452568 285628 452572
rect 285692 452570 285698 452572
rect 285581 452512 285586 452568
rect 285581 452508 285628 452512
rect 285692 452510 285738 452570
rect 285692 452508 285698 452510
rect 288198 452508 288204 452572
rect 288268 452570 288274 452572
rect 288341 452570 288407 452573
rect 288268 452568 288407 452570
rect 288268 452512 288346 452568
rect 288402 452512 288407 452568
rect 288268 452510 288407 452512
rect 288268 452508 288274 452510
rect 285581 452507 285647 452508
rect 288341 452507 288407 452510
rect 290590 452508 290596 452572
rect 290660 452570 290666 452572
rect 291101 452570 291167 452573
rect 290660 452568 291167 452570
rect 290660 452512 291106 452568
rect 291162 452512 291167 452568
rect 290660 452510 291167 452512
rect 290660 452508 290666 452510
rect 291101 452507 291167 452510
rect 292573 452572 292639 452573
rect 293033 452572 293099 452573
rect 292573 452568 292620 452572
rect 292684 452570 292690 452572
rect 292982 452570 292988 452572
rect 292573 452512 292578 452568
rect 292573 452508 292620 452512
rect 292684 452510 292730 452570
rect 292942 452510 292988 452570
rect 293052 452568 293099 452572
rect 293094 452512 293099 452568
rect 292684 452508 292690 452510
rect 292982 452508 292988 452510
rect 293052 452508 293099 452512
rect 295558 452508 295564 452572
rect 295628 452570 295634 452572
rect 296621 452570 296687 452573
rect 295628 452568 296687 452570
rect 295628 452512 296626 452568
rect 296682 452512 296687 452568
rect 295628 452510 296687 452512
rect 295628 452508 295634 452510
rect 292573 452507 292639 452508
rect 293033 452507 293099 452508
rect 296621 452507 296687 452510
rect 298134 452508 298140 452572
rect 298204 452570 298210 452572
rect 299381 452570 299447 452573
rect 298204 452568 299447 452570
rect 298204 452512 299386 452568
rect 299442 452512 299447 452568
rect 298204 452510 299447 452512
rect 298204 452508 298210 452510
rect 299381 452507 299447 452510
rect 300342 452508 300348 452572
rect 300412 452570 300418 452572
rect 300761 452570 300827 452573
rect 300412 452568 300827 452570
rect 300412 452512 300766 452568
rect 300822 452512 300827 452568
rect 300412 452510 300827 452512
rect 300412 452508 300418 452510
rect 300761 452507 300827 452510
rect 301957 452572 302023 452573
rect 303061 452572 303127 452573
rect 304165 452572 304231 452573
rect 305269 452572 305335 452573
rect 306373 452572 306439 452573
rect 307845 452572 307911 452573
rect 308949 452572 309015 452573
rect 309869 452572 309935 452573
rect 313365 452572 313431 452573
rect 314653 452572 314719 452573
rect 301957 452568 302004 452572
rect 302068 452570 302074 452572
rect 301957 452512 301962 452568
rect 301957 452508 302004 452512
rect 302068 452510 302114 452570
rect 303061 452568 303108 452572
rect 303172 452570 303178 452572
rect 303061 452512 303066 452568
rect 302068 452508 302074 452510
rect 303061 452508 303108 452512
rect 303172 452510 303218 452570
rect 304165 452568 304212 452572
rect 304276 452570 304282 452572
rect 304165 452512 304170 452568
rect 303172 452508 303178 452510
rect 304165 452508 304212 452512
rect 304276 452510 304322 452570
rect 305269 452568 305316 452572
rect 305380 452570 305386 452572
rect 305269 452512 305274 452568
rect 304276 452508 304282 452510
rect 305269 452508 305316 452512
rect 305380 452510 305426 452570
rect 306373 452568 306420 452572
rect 306484 452570 306490 452572
rect 306373 452512 306378 452568
rect 305380 452508 305386 452510
rect 306373 452508 306420 452512
rect 306484 452510 306530 452570
rect 307845 452568 307892 452572
rect 307956 452570 307962 452572
rect 307845 452512 307850 452568
rect 306484 452508 306490 452510
rect 307845 452508 307892 452512
rect 307956 452510 308002 452570
rect 308949 452568 308996 452572
rect 309060 452570 309066 452572
rect 308949 452512 308954 452568
rect 307956 452508 307962 452510
rect 308949 452508 308996 452512
rect 309060 452510 309106 452570
rect 309869 452568 309916 452572
rect 309980 452570 309986 452572
rect 309869 452512 309874 452568
rect 309060 452508 309066 452510
rect 309869 452508 309916 452512
rect 309980 452510 310026 452570
rect 313365 452568 313412 452572
rect 313476 452570 313482 452572
rect 313365 452512 313370 452568
rect 309980 452508 309986 452510
rect 313365 452508 313412 452512
rect 313476 452510 313522 452570
rect 314653 452568 314700 452572
rect 314764 452570 314770 452572
rect 315982 452570 315988 452572
rect 314653 452512 314658 452568
rect 313476 452508 313482 452510
rect 314653 452508 314700 452512
rect 314764 452510 315988 452570
rect 314764 452508 314770 452510
rect 315982 452508 315988 452510
rect 316052 452570 316058 452572
rect 316902 452570 316908 452572
rect 316052 452510 316908 452570
rect 316052 452508 316058 452510
rect 316902 452508 316908 452510
rect 316972 452570 316978 452572
rect 318374 452570 318380 452572
rect 316972 452510 318380 452570
rect 316972 452508 316978 452510
rect 318374 452508 318380 452510
rect 318444 452508 318450 452572
rect 320173 452570 320239 452573
rect 320398 452570 320404 452572
rect 320173 452568 320404 452570
rect 320173 452512 320178 452568
rect 320234 452512 320404 452568
rect 320173 452510 320404 452512
rect 301957 452507 302023 452508
rect 303061 452507 303127 452508
rect 304165 452507 304231 452508
rect 305269 452507 305335 452508
rect 306373 452507 306439 452508
rect 307845 452507 307911 452508
rect 308949 452507 309015 452508
rect 309869 452507 309935 452508
rect 313365 452507 313431 452508
rect 314653 452507 314719 452508
rect 320173 452507 320239 452510
rect 320398 452508 320404 452510
rect 320468 452508 320474 452572
rect 425421 452570 425487 452573
rect 426014 452570 426020 452572
rect 425421 452568 426020 452570
rect 425421 452512 425426 452568
rect 425482 452512 426020 452568
rect 425421 452510 426020 452512
rect 425421 452507 425487 452510
rect 426014 452508 426020 452510
rect 426084 452508 426090 452572
rect 426893 452570 426959 452573
rect 427118 452570 427124 452572
rect 426893 452568 427124 452570
rect 426893 452512 426898 452568
rect 426954 452512 427124 452568
rect 426893 452510 427124 452512
rect 426893 452507 426959 452510
rect 427118 452508 427124 452510
rect 427188 452508 427194 452572
rect 428222 452508 428228 452572
rect 428292 452570 428298 452572
rect 428457 452570 428523 452573
rect 429510 452570 429516 452572
rect 428292 452568 429516 452570
rect 428292 452512 428462 452568
rect 428518 452512 429516 452568
rect 428292 452510 429516 452512
rect 428292 452508 428298 452510
rect 428457 452507 428523 452510
rect 429510 452508 429516 452510
rect 429580 452508 429586 452572
rect 432045 452570 432111 452573
rect 433006 452570 433012 452572
rect 432045 452568 433012 452570
rect 432045 452512 432050 452568
rect 432106 452512 433012 452568
rect 432045 452510 433012 452512
rect 432045 452507 432111 452510
rect 433006 452508 433012 452510
rect 433076 452508 433082 452572
rect 433701 452570 433767 452573
rect 434110 452570 434116 452572
rect 433701 452568 434116 452570
rect 433701 452512 433706 452568
rect 433762 452512 434116 452568
rect 433701 452510 434116 452512
rect 433701 452507 433767 452510
rect 434110 452508 434116 452510
rect 434180 452508 434186 452572
rect 434713 452570 434779 452573
rect 435398 452570 435404 452572
rect 434713 452568 435404 452570
rect 434713 452512 434718 452568
rect 434774 452512 435404 452568
rect 434713 452510 435404 452512
rect 434713 452507 434779 452510
rect 435398 452508 435404 452510
rect 435468 452508 435474 452572
rect 436277 452570 436343 452573
rect 436502 452570 436508 452572
rect 436277 452568 436508 452570
rect 436277 452512 436282 452568
rect 436338 452512 436508 452568
rect 436277 452510 436508 452512
rect 436277 452507 436343 452510
rect 436502 452508 436508 452510
rect 436572 452508 436578 452572
rect 450261 452570 450327 452573
rect 452837 452572 452903 452573
rect 466177 452572 466243 452573
rect 450670 452570 450676 452572
rect 450261 452568 450676 452570
rect 450261 452512 450266 452568
rect 450322 452512 450676 452568
rect 450261 452510 450676 452512
rect 450261 452507 450327 452510
rect 450670 452508 450676 452510
rect 450740 452508 450746 452572
rect 452837 452568 452884 452572
rect 452948 452570 452954 452572
rect 466126 452570 466132 452572
rect 452837 452512 452842 452568
rect 452837 452508 452884 452512
rect 452948 452510 452994 452570
rect 466086 452510 466132 452570
rect 466196 452568 466243 452572
rect 466238 452512 466243 452568
rect 452948 452508 452954 452510
rect 466126 452508 466132 452510
rect 466196 452508 466243 452512
rect 452837 452507 452903 452508
rect 466177 452507 466243 452508
rect 466545 452570 466611 452573
rect 467925 452572 467991 452573
rect 467046 452570 467052 452572
rect 466545 452568 467052 452570
rect 466545 452512 466550 452568
rect 466606 452512 467052 452568
rect 466545 452510 467052 452512
rect 466545 452507 466611 452510
rect 467046 452508 467052 452510
rect 467116 452508 467122 452572
rect 467925 452568 467972 452572
rect 468036 452570 468042 452572
rect 467925 452512 467930 452568
rect 467925 452508 467972 452512
rect 468036 452510 468082 452570
rect 468036 452508 468042 452510
rect 468518 452508 468524 452572
rect 468588 452570 468594 452572
rect 468661 452570 468727 452573
rect 468588 452568 468727 452570
rect 468588 452512 468666 452568
rect 468722 452512 468727 452568
rect 468588 452510 468727 452512
rect 468588 452508 468594 452510
rect 467925 452507 467991 452508
rect 468661 452507 468727 452510
rect 470910 452508 470916 452572
rect 470980 452570 470986 452572
rect 471881 452570 471947 452573
rect 473537 452572 473603 452573
rect 473486 452570 473492 452572
rect 470980 452568 471947 452570
rect 470980 452512 471886 452568
rect 471942 452512 471947 452568
rect 470980 452510 471947 452512
rect 473446 452510 473492 452570
rect 473556 452568 473603 452572
rect 473598 452512 473603 452568
rect 470980 452508 470986 452510
rect 471881 452507 471947 452510
rect 473486 452508 473492 452510
rect 473556 452508 473603 452512
rect 473537 452507 473603 452508
rect 476021 452572 476087 452573
rect 476021 452568 476068 452572
rect 476132 452570 476138 452572
rect 476021 452512 476026 452568
rect 476021 452508 476068 452512
rect 476132 452510 476178 452570
rect 476132 452508 476138 452510
rect 478270 452508 478276 452572
rect 478340 452570 478346 452572
rect 478413 452570 478479 452573
rect 481081 452572 481147 452573
rect 483473 452572 483539 452573
rect 481030 452570 481036 452572
rect 478340 452568 478479 452570
rect 478340 452512 478418 452568
rect 478474 452512 478479 452568
rect 478340 452510 478479 452512
rect 480990 452510 481036 452570
rect 481100 452568 481147 452572
rect 483422 452570 483428 452572
rect 481142 452512 481147 452568
rect 478340 452508 478346 452510
rect 476021 452507 476087 452508
rect 478413 452507 478479 452510
rect 481030 452508 481036 452510
rect 481100 452508 481147 452512
rect 483382 452510 483428 452570
rect 483492 452568 483539 452572
rect 483534 452512 483539 452568
rect 483422 452508 483428 452510
rect 483492 452508 483539 452512
rect 485998 452508 486004 452572
rect 486068 452570 486074 452572
rect 487061 452570 487127 452573
rect 488441 452572 488507 452573
rect 491017 452572 491083 452573
rect 493593 452572 493659 452573
rect 495985 452572 496051 452573
rect 488390 452570 488396 452572
rect 486068 452568 487127 452570
rect 486068 452512 487066 452568
rect 487122 452512 487127 452568
rect 486068 452510 487127 452512
rect 488350 452510 488396 452570
rect 488460 452568 488507 452572
rect 490966 452570 490972 452572
rect 488502 452512 488507 452568
rect 486068 452508 486074 452510
rect 481081 452507 481147 452508
rect 483473 452507 483539 452508
rect 487061 452507 487127 452510
rect 488390 452508 488396 452510
rect 488460 452508 488507 452512
rect 490926 452510 490972 452570
rect 491036 452568 491083 452572
rect 493542 452570 493548 452572
rect 491078 452512 491083 452568
rect 490966 452508 490972 452510
rect 491036 452508 491083 452512
rect 493502 452510 493548 452570
rect 493612 452568 493659 452572
rect 495934 452570 495940 452572
rect 493654 452512 493659 452568
rect 493542 452508 493548 452510
rect 493612 452508 493659 452512
rect 495894 452510 495940 452570
rect 496004 452568 496051 452572
rect 496046 452512 496051 452568
rect 495934 452508 495940 452510
rect 496004 452508 496051 452512
rect 498510 452508 498516 452572
rect 498580 452570 498586 452572
rect 499481 452570 499547 452573
rect 498580 452568 499547 452570
rect 498580 452512 499486 452568
rect 499542 452512 499547 452568
rect 498580 452510 499547 452512
rect 498580 452508 498586 452510
rect 488441 452507 488507 452508
rect 491017 452507 491083 452508
rect 493593 452507 493659 452508
rect 495985 452507 496051 452508
rect 499481 452507 499547 452510
rect 501086 452508 501092 452572
rect 501156 452570 501162 452572
rect 501229 452570 501295 452573
rect 503529 452572 503595 452573
rect 505921 452572 505987 452573
rect 503478 452570 503484 452572
rect 501156 452568 501295 452570
rect 501156 452512 501234 452568
rect 501290 452512 501295 452568
rect 501156 452510 501295 452512
rect 503438 452510 503484 452570
rect 503548 452568 503595 452572
rect 505870 452570 505876 452572
rect 503590 452512 503595 452568
rect 501156 452508 501162 452510
rect 501229 452507 501295 452510
rect 503478 452508 503484 452510
rect 503548 452508 503595 452512
rect 505830 452510 505876 452570
rect 505940 452568 505987 452572
rect 505982 452512 505987 452568
rect 505870 452508 505876 452510
rect 505940 452508 505987 452512
rect 508446 452508 508452 452572
rect 508516 452570 508522 452572
rect 509141 452570 509207 452573
rect 508516 452568 509207 452570
rect 508516 452512 509146 452568
rect 509202 452512 509207 452568
rect 508516 452510 509207 452512
rect 508516 452508 508522 452510
rect 503529 452507 503595 452508
rect 505921 452507 505987 452508
rect 509141 452507 509207 452510
rect 511022 452508 511028 452572
rect 511092 452570 511098 452572
rect 511901 452570 511967 452573
rect 511092 452568 511967 452570
rect 511092 452512 511906 452568
rect 511962 452512 511967 452568
rect 511092 452510 511967 452512
rect 511092 452508 511098 452510
rect 511901 452507 511967 452510
rect 513414 452508 513420 452572
rect 513484 452570 513490 452572
rect 514661 452570 514727 452573
rect 516041 452572 516107 452573
rect 515990 452570 515996 452572
rect 513484 452568 514727 452570
rect 513484 452512 514666 452568
rect 514722 452512 514727 452568
rect 513484 452510 514727 452512
rect 515950 452510 515996 452570
rect 516060 452568 516107 452572
rect 516102 452512 516107 452568
rect 513484 452508 513490 452510
rect 514661 452507 514727 452510
rect 515990 452508 515996 452510
rect 516060 452508 516107 452512
rect 516041 452507 516107 452508
rect 213361 452436 213427 452437
rect 213310 452434 213316 452436
rect 213234 452374 213316 452434
rect 213380 452434 213427 452436
rect 533286 452434 533292 452436
rect 213380 452432 533292 452434
rect 213422 452376 533292 452432
rect 213310 452372 213316 452374
rect 213380 452374 533292 452376
rect 213380 452372 213427 452374
rect 533286 452372 533292 452374
rect 533356 452372 533362 452436
rect 213361 452371 213427 452372
rect 283189 452300 283255 452301
rect 198958 452236 198964 452300
rect 199028 452298 199034 452300
rect 280838 452298 280844 452300
rect 199028 452238 280844 452298
rect 199028 452236 199034 452238
rect 280838 452236 280844 452238
rect 280908 452236 280914 452300
rect 283189 452296 283236 452300
rect 283300 452298 283306 452300
rect 287830 452298 287836 452300
rect 283189 452240 283194 452296
rect 283189 452236 283236 452240
rect 283300 452238 283346 452298
rect 287010 452238 287836 452298
rect 283300 452236 283306 452238
rect 283189 452235 283255 452236
rect 197302 452100 197308 452164
rect 197372 452162 197378 452164
rect 277158 452162 277164 452164
rect 197372 452102 277164 452162
rect 197372 452100 197378 452102
rect 277158 452100 277164 452102
rect 277228 452100 277234 452164
rect 281441 452162 281507 452165
rect 287010 452162 287070 452238
rect 287830 452236 287836 452238
rect 287900 452236 287906 452300
rect 300117 452298 300183 452301
rect 300710 452298 300716 452300
rect 300117 452296 300716 452298
rect 300117 452240 300122 452296
rect 300178 452240 300716 452296
rect 300117 452238 300716 452240
rect 300117 452235 300183 452238
rect 300710 452236 300716 452238
rect 300780 452236 300786 452300
rect 302918 452236 302924 452300
rect 302988 452298 302994 452300
rect 303521 452298 303587 452301
rect 302988 452296 303587 452298
rect 302988 452240 303526 452296
rect 303582 452240 303587 452296
rect 302988 452238 303587 452240
rect 302988 452236 302994 452238
rect 303521 452235 303587 452238
rect 305862 452236 305868 452300
rect 305932 452298 305938 452300
rect 306281 452298 306347 452301
rect 305932 452296 306347 452298
rect 305932 452240 306286 452296
rect 306342 452240 306347 452296
rect 305932 452238 306347 452240
rect 305932 452236 305938 452238
rect 306281 452235 306347 452238
rect 319437 452300 319503 452301
rect 319437 452296 319484 452300
rect 319548 452298 319554 452300
rect 319437 452240 319442 452296
rect 319437 452236 319484 452240
rect 319548 452238 319594 452298
rect 319548 452236 319554 452238
rect 438342 452236 438348 452300
rect 438412 452298 438418 452300
rect 438669 452298 438735 452301
rect 438412 452296 438735 452298
rect 438412 452240 438674 452296
rect 438730 452240 438735 452296
rect 438412 452238 438735 452240
rect 438412 452236 438418 452238
rect 319437 452235 319503 452236
rect 438669 452235 438735 452238
rect 454125 452298 454191 452301
rect 455270 452298 455276 452300
rect 454125 452296 455276 452298
rect 454125 452240 454130 452296
rect 454186 452240 455276 452296
rect 454125 452238 455276 452240
rect 454125 452235 454191 452238
rect 455270 452236 455276 452238
rect 455340 452236 455346 452300
rect 462313 452298 462379 452301
rect 463366 452298 463372 452300
rect 462313 452296 463372 452298
rect 462313 452240 462318 452296
rect 462374 452240 463372 452296
rect 462313 452238 463372 452240
rect 462313 452235 462379 452238
rect 463366 452236 463372 452238
rect 463436 452236 463442 452300
rect 468017 452298 468083 452301
rect 469070 452298 469076 452300
rect 468017 452296 469076 452298
rect 468017 452240 468022 452296
rect 468078 452240 469076 452296
rect 468017 452238 469076 452240
rect 468017 452235 468083 452238
rect 469070 452236 469076 452238
rect 469140 452236 469146 452300
rect 281441 452160 287070 452162
rect 281441 452104 281446 452160
rect 281502 452104 287070 452160
rect 281441 452102 287070 452104
rect 297357 452162 297423 452165
rect 405365 452162 405431 452165
rect 297357 452160 405431 452162
rect 297357 452104 297362 452160
rect 297418 452104 405370 452160
rect 405426 452104 405431 452160
rect 297357 452102 405431 452104
rect 281441 452099 281507 452102
rect 297357 452099 297423 452102
rect 405365 452099 405431 452102
rect 441613 452162 441679 452165
rect 442390 452162 442396 452164
rect 441613 452160 442396 452162
rect 441613 452104 441618 452160
rect 441674 452104 442396 452160
rect 441613 452102 442396 452104
rect 441613 452099 441679 452102
rect 442390 452100 442396 452102
rect 442460 452100 442466 452164
rect 442993 452162 443059 452165
rect 443494 452162 443500 452164
rect 442993 452160 443500 452162
rect 442993 452104 442998 452160
rect 443054 452104 443500 452160
rect 442993 452102 443500 452104
rect 442993 452099 443059 452102
rect 443494 452100 443500 452102
rect 443564 452100 443570 452164
rect 445753 452162 445819 452165
rect 445886 452162 445892 452164
rect 445753 452160 445892 452162
rect 445753 452104 445758 452160
rect 445814 452104 445892 452160
rect 445753 452102 445892 452104
rect 445753 452099 445819 452102
rect 445886 452100 445892 452102
rect 445956 452100 445962 452164
rect 446070 452100 446076 452164
rect 446140 452162 446146 452164
rect 447041 452162 447107 452165
rect 446140 452160 447107 452162
rect 446140 452104 447046 452160
rect 447102 452104 447107 452160
rect 446140 452102 447107 452104
rect 446140 452100 446146 452102
rect 447041 452099 447107 452102
rect 448605 452162 448671 452165
rect 449382 452162 449388 452164
rect 448605 452160 449388 452162
rect 448605 452104 448610 452160
rect 448666 452104 449388 452160
rect 448605 452102 449388 452104
rect 448605 452099 448671 452102
rect 449382 452100 449388 452102
rect 449452 452100 449458 452164
rect 451365 452162 451431 452165
rect 453665 452164 453731 452165
rect 451774 452162 451780 452164
rect 451365 452160 451780 452162
rect 451365 452104 451370 452160
rect 451426 452104 451780 452160
rect 451365 452102 451780 452104
rect 451365 452099 451431 452102
rect 451774 452100 451780 452102
rect 451844 452100 451850 452164
rect 453614 452162 453620 452164
rect 453574 452102 453620 452162
rect 453684 452160 453731 452164
rect 453726 452104 453731 452160
rect 453614 452100 453620 452102
rect 453684 452100 453731 452104
rect 456006 452100 456012 452164
rect 456076 452162 456082 452164
rect 456701 452162 456767 452165
rect 459737 452164 459803 452165
rect 459686 452162 459692 452164
rect 456076 452160 456767 452162
rect 456076 452104 456706 452160
rect 456762 452104 456767 452160
rect 456076 452102 456767 452104
rect 459646 452102 459692 452162
rect 459756 452160 459803 452164
rect 459798 452104 459803 452160
rect 456076 452100 456082 452102
rect 453665 452099 453731 452100
rect 456701 452099 456767 452102
rect 459686 452100 459692 452102
rect 459756 452100 459803 452104
rect 462262 452100 462268 452164
rect 462332 452162 462338 452164
rect 462405 452162 462471 452165
rect 463601 452164 463667 452165
rect 463550 452162 463556 452164
rect 462332 452160 462471 452162
rect 462332 452104 462410 452160
rect 462466 452104 462471 452160
rect 462332 452102 462471 452104
rect 463510 452102 463556 452162
rect 463620 452160 463667 452164
rect 463662 452104 463667 452160
rect 462332 452100 462338 452102
rect 459737 452099 459803 452100
rect 462405 452099 462471 452102
rect 463550 452100 463556 452102
rect 463620 452100 463667 452104
rect 463601 452099 463667 452100
rect 465073 452162 465139 452165
rect 465758 452162 465764 452164
rect 465073 452160 465764 452162
rect 465073 452104 465078 452160
rect 465134 452104 465764 452160
rect 465073 452102 465764 452104
rect 465073 452099 465139 452102
rect 465758 452100 465764 452102
rect 465828 452100 465834 452164
rect 198774 451964 198780 452028
rect 198844 452026 198850 452028
rect 294781 452026 294847 452029
rect 405549 452026 405615 452029
rect 198844 451966 258090 452026
rect 198844 451964 198850 451966
rect 45645 451890 45711 451893
rect 46790 451890 46796 451892
rect 45645 451888 46796 451890
rect 45645 451832 45650 451888
rect 45706 451832 46796 451888
rect 45645 451830 46796 451832
rect 45645 451827 45711 451830
rect 46790 451828 46796 451830
rect 46860 451828 46866 451892
rect 167269 451890 167335 451893
rect 167494 451890 167500 451892
rect 167269 451888 167500 451890
rect 167269 451832 167274 451888
rect 167330 451832 167500 451888
rect 167269 451830 167500 451832
rect 167269 451827 167335 451830
rect 167494 451828 167500 451830
rect 167564 451828 167570 451892
rect 258030 451890 258090 451966
rect 294781 452024 405615 452026
rect 294781 451968 294786 452024
rect 294842 451968 405554 452024
rect 405610 451968 405615 452024
rect 294781 451966 405615 451968
rect 294781 451963 294847 451966
rect 405549 451963 405615 451966
rect 278446 451890 278452 451892
rect 258030 451830 278452 451890
rect 278446 451828 278452 451830
rect 278516 451828 278522 451892
rect 293585 451890 293651 451893
rect 408217 451890 408283 451893
rect 293585 451888 408283 451890
rect 293585 451832 293590 451888
rect 293646 451832 408222 451888
rect 408278 451832 408283 451888
rect 293585 451830 408283 451832
rect 293585 451827 293651 451830
rect 408217 451827 408283 451830
rect 437657 451618 437723 451621
rect 438710 451618 438716 451620
rect 437657 451616 438716 451618
rect 437657 451560 437662 451616
rect 437718 451560 438716 451616
rect 437657 451558 438716 451560
rect 437657 451555 437723 451558
rect 438710 451556 438716 451558
rect 438780 451556 438786 451620
rect 440233 451618 440299 451621
rect 441286 451618 441292 451620
rect 440233 451616 441292 451618
rect 440233 451560 440238 451616
rect 440294 451560 441292 451616
rect 440233 451558 441292 451560
rect 440233 451555 440299 451558
rect 441286 451556 441292 451558
rect 441356 451556 441362 451620
rect 458398 451556 458404 451620
rect 458468 451618 458474 451620
rect 459461 451618 459527 451621
rect 458468 451616 459527 451618
rect 458468 451560 459466 451616
rect 459522 451560 459527 451616
rect 458468 451558 459527 451560
rect 458468 451556 458474 451558
rect 459461 451555 459527 451558
rect 213177 451482 213243 451485
rect 532734 451482 532740 451484
rect 213177 451480 532740 451482
rect 213177 451424 213182 451480
rect 213238 451424 532740 451480
rect 213177 451422 532740 451424
rect 213177 451419 213243 451422
rect 532734 451420 532740 451422
rect 532804 451420 532810 451484
rect 48037 451348 48103 451349
rect 48037 451346 48084 451348
rect 47992 451344 48084 451346
rect 47992 451288 48042 451344
rect 47992 451286 48084 451288
rect 48037 451284 48084 451286
rect 48148 451284 48154 451348
rect 248086 451284 248092 451348
rect 248156 451346 248162 451348
rect 248229 451346 248295 451349
rect 248156 451344 248295 451346
rect 248156 451288 248234 451344
rect 248290 451288 248295 451344
rect 248156 451286 248295 451288
rect 248156 451284 248162 451286
rect 48037 451283 48103 451284
rect 248229 451283 248295 451286
rect 250662 451284 250668 451348
rect 250732 451346 250738 451348
rect 251081 451346 251147 451349
rect 250732 451344 251147 451346
rect 250732 451288 251086 451344
rect 251142 451288 251147 451344
rect 250732 451286 251147 451288
rect 250732 451284 250738 451286
rect 251081 451283 251147 451286
rect 258022 451284 258028 451348
rect 258092 451346 258098 451348
rect 259361 451346 259427 451349
rect 258092 451344 259427 451346
rect 258092 451288 259366 451344
rect 259422 451288 259427 451344
rect 258092 451286 259427 451288
rect 258092 451284 258098 451286
rect 259361 451283 259427 451286
rect 308254 451284 308260 451348
rect 308324 451346 308330 451348
rect 309041 451346 309107 451349
rect 308324 451344 309107 451346
rect 308324 451288 309046 451344
rect 309102 451288 309107 451344
rect 308324 451286 309107 451288
rect 308324 451284 308330 451286
rect 309041 451283 309107 451286
rect 437565 451348 437631 451349
rect 437565 451344 437612 451348
rect 437676 451346 437682 451348
rect 438945 451346 439011 451349
rect 439998 451346 440004 451348
rect 437565 451288 437570 451344
rect 437565 451284 437612 451288
rect 437676 451286 437722 451346
rect 438945 451344 440004 451346
rect 438945 451288 438950 451344
rect 439006 451288 440004 451344
rect 438945 451286 440004 451288
rect 437676 451284 437682 451286
rect 437565 451283 437631 451284
rect 438945 451283 439011 451286
rect 439998 451284 440004 451286
rect 440068 451284 440074 451348
rect 440734 451284 440740 451348
rect 440804 451346 440810 451348
rect 441521 451346 441587 451349
rect 440804 451344 441587 451346
rect 440804 451288 441526 451344
rect 441582 451288 441587 451344
rect 440804 451286 441587 451288
rect 440804 451284 440810 451286
rect 441521 451283 441587 451286
rect 444465 451346 444531 451349
rect 444598 451346 444604 451348
rect 444465 451344 444604 451346
rect 444465 451288 444470 451344
rect 444526 451288 444604 451344
rect 444465 451286 444604 451288
rect 444465 451283 444531 451286
rect 444598 451284 444604 451286
rect 444668 451284 444674 451348
rect 445845 451346 445911 451349
rect 446990 451346 446996 451348
rect 445845 451344 446996 451346
rect 445845 451288 445850 451344
rect 445906 451288 446996 451344
rect 445845 451286 446996 451288
rect 445845 451283 445911 451286
rect 446990 451284 446996 451286
rect 447060 451284 447066 451348
rect 447225 451346 447291 451349
rect 448513 451348 448579 451349
rect 448094 451346 448100 451348
rect 447225 451344 448100 451346
rect 447225 451288 447230 451344
rect 447286 451288 448100 451344
rect 447225 451286 448100 451288
rect 447225 451283 447291 451286
rect 448094 451284 448100 451286
rect 448164 451284 448170 451348
rect 448462 451346 448468 451348
rect 448422 451286 448468 451346
rect 448532 451344 448579 451348
rect 448574 451288 448579 451344
rect 448462 451284 448468 451286
rect 448532 451284 448579 451288
rect 451038 451284 451044 451348
rect 451108 451346 451114 451348
rect 451181 451346 451247 451349
rect 451108 451344 451247 451346
rect 451108 451288 451186 451344
rect 451242 451288 451247 451344
rect 451108 451286 451247 451288
rect 451108 451284 451114 451286
rect 448513 451283 448579 451284
rect 451181 451283 451247 451286
rect 452745 451346 452811 451349
rect 453982 451346 453988 451348
rect 452745 451344 453988 451346
rect 452745 451288 452750 451344
rect 452806 451288 453988 451344
rect 452745 451286 453988 451288
rect 452745 451283 452811 451286
rect 453982 451284 453988 451286
rect 454052 451284 454058 451348
rect 455505 451346 455571 451349
rect 456374 451346 456380 451348
rect 455505 451344 456380 451346
rect 455505 451288 455510 451344
rect 455566 451288 456380 451344
rect 455505 451286 456380 451288
rect 455505 451283 455571 451286
rect 456374 451284 456380 451286
rect 456444 451284 456450 451348
rect 456885 451346 456951 451349
rect 457662 451346 457668 451348
rect 456885 451344 457668 451346
rect 456885 451288 456890 451344
rect 456946 451288 457668 451344
rect 456885 451286 457668 451288
rect 456885 451283 456951 451286
rect 457662 451284 457668 451286
rect 457732 451284 457738 451348
rect 458265 451346 458331 451349
rect 458582 451346 458588 451348
rect 458265 451344 458588 451346
rect 458265 451288 458270 451344
rect 458326 451288 458588 451344
rect 458265 451286 458588 451288
rect 458265 451283 458331 451286
rect 458582 451284 458588 451286
rect 458652 451284 458658 451348
rect 463785 451346 463851 451349
rect 464286 451346 464292 451348
rect 463785 451344 464292 451346
rect 463785 451288 463790 451344
rect 463846 451288 464292 451344
rect 463785 451286 464292 451288
rect 463785 451283 463851 451286
rect 464286 451284 464292 451286
rect 464356 451284 464362 451348
rect 170305 451210 170371 451213
rect 170438 451210 170444 451212
rect 170305 451208 170444 451210
rect 170305 451152 170310 451208
rect 170366 451152 170444 451208
rect 170305 451150 170444 451152
rect 170305 451147 170371 451150
rect 170438 451148 170444 451150
rect 170508 451148 170514 451212
rect 3417 450938 3483 450941
rect 341517 450938 341583 450941
rect 3417 450936 341583 450938
rect 3417 450880 3422 450936
rect 3478 450880 341522 450936
rect 341578 450880 341583 450936
rect 3417 450878 341583 450880
rect 3417 450875 3483 450878
rect 341517 450875 341583 450878
rect 28257 450802 28323 450805
rect 433149 450802 433215 450805
rect 28257 450800 433215 450802
rect 28257 450744 28262 450800
rect 28318 450744 433154 450800
rect 433210 450744 433215 450800
rect 28257 450742 433215 450744
rect 28257 450739 28323 450742
rect 433149 450739 433215 450742
rect 21357 450666 21423 450669
rect 438117 450666 438183 450669
rect 21357 450664 438183 450666
rect 21357 450608 21362 450664
rect 21418 450608 438122 450664
rect 438178 450608 438183 450664
rect 21357 450606 438183 450608
rect 21357 450603 21423 450606
rect 438117 450603 438183 450606
rect 23473 450530 23539 450533
rect 445661 450530 445727 450533
rect 23473 450528 445727 450530
rect 23473 450472 23478 450528
rect 23534 450472 445666 450528
rect 445722 450472 445727 450528
rect 23473 450470 445727 450472
rect 23473 450467 23539 450470
rect 445661 450467 445727 450470
rect 165429 449986 165495 449989
rect 167126 449986 167132 449988
rect 165429 449984 167132 449986
rect 165429 449928 165434 449984
rect 165490 449928 167132 449984
rect 165429 449926 167132 449928
rect 165429 449923 165495 449926
rect 167126 449924 167132 449926
rect 167196 449924 167202 449988
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 461025 449306 461091 449309
rect 461158 449306 461164 449308
rect 461025 449304 461164 449306
rect 461025 449248 461030 449304
rect 461086 449248 461164 449304
rect 461025 449246 461164 449248
rect 461025 449243 461091 449246
rect 461158 449244 461164 449246
rect 461228 449244 461234 449308
rect 460974 449108 460980 449172
rect 461044 449170 461050 449172
rect 462221 449170 462287 449173
rect 461044 449168 462287 449170
rect 461044 449112 462226 449168
rect 462282 449112 462287 449168
rect 461044 449110 462287 449112
rect 461044 449108 461050 449110
rect 462221 449107 462287 449110
rect 168598 448564 168604 448628
rect 168668 448626 168674 448628
rect 168833 448626 168899 448629
rect 168668 448624 168899 448626
rect 168668 448568 168838 448624
rect 168894 448568 168899 448624
rect 168668 448566 168899 448568
rect 168668 448564 168674 448566
rect 168833 448563 168899 448566
rect 197997 448490 198063 448493
rect 549621 448490 549687 448493
rect 197997 448488 549687 448490
rect 197997 448432 198002 448488
rect 198058 448432 549626 448488
rect 549682 448432 549687 448488
rect 197997 448430 549687 448432
rect 197997 448427 198063 448430
rect 549621 448427 549687 448430
rect 198089 448354 198155 448357
rect 549529 448354 549595 448357
rect 198089 448352 549595 448354
rect 198089 448296 198094 448352
rect 198150 448296 549534 448352
rect 549590 448296 549595 448352
rect 198089 448294 549595 448296
rect 198089 448291 198155 448294
rect 549529 448291 549595 448294
rect 198181 448218 198247 448221
rect 549437 448218 549503 448221
rect 198181 448216 549503 448218
rect 198181 448160 198186 448216
rect 198242 448160 549442 448216
rect 549498 448160 549503 448216
rect 198181 448158 549503 448160
rect 198181 448155 198247 448158
rect 549437 448155 549503 448158
rect 198273 448082 198339 448085
rect 549345 448082 549411 448085
rect 198273 448080 549411 448082
rect 198273 448024 198278 448080
rect 198334 448024 549350 448080
rect 549406 448024 549411 448080
rect 198273 448022 549411 448024
rect 198273 448019 198339 448022
rect 549345 448019 549411 448022
rect 174670 447884 174676 447948
rect 174740 447946 174746 447948
rect 204529 447946 204595 447949
rect 174740 447944 204595 447946
rect 174740 447888 204534 447944
rect 204590 447888 204595 447944
rect 174740 447886 204595 447888
rect 174740 447884 174746 447886
rect 204529 447883 204595 447886
rect 249517 447946 249583 447949
rect 338246 447946 338252 447948
rect 249517 447944 338252 447946
rect 249517 447888 249522 447944
rect 249578 447888 338252 447944
rect 249517 447886 338252 447888
rect 249517 447883 249583 447886
rect 338246 447884 338252 447886
rect 338316 447884 338322 447948
rect 240777 447810 240843 447813
rect 336958 447810 336964 447812
rect 240777 447808 336964 447810
rect 240777 447752 240782 447808
rect 240838 447752 336964 447808
rect 240777 447750 336964 447752
rect 240777 447747 240843 447750
rect 336958 447748 336964 447750
rect 337028 447748 337034 447812
rect 250805 447674 250871 447677
rect 336774 447674 336780 447676
rect 250805 447672 336780 447674
rect 250805 447616 250810 447672
rect 250866 447616 336780 447672
rect 250805 447614 336780 447616
rect 250805 447611 250871 447614
rect 336774 447612 336780 447614
rect 336844 447612 336850 447676
rect 193121 445362 193187 445365
rect 206829 445362 206895 445365
rect 193121 445360 206895 445362
rect 193121 445304 193126 445360
rect 193182 445304 206834 445360
rect 206890 445304 206895 445360
rect 193121 445302 206895 445304
rect 193121 445299 193187 445302
rect 206829 445299 206895 445302
rect 28717 445226 28783 445229
rect 194317 445226 194383 445229
rect 208025 445226 208091 445229
rect 28717 445224 30062 445226
rect 28717 445168 28722 445224
rect 28778 445168 30062 445224
rect 28717 445166 30062 445168
rect 194317 445224 208091 445226
rect 194317 445168 194322 445224
rect 194378 445168 208030 445224
rect 208086 445168 208091 445224
rect 194317 445166 208091 445168
rect 28717 445163 28783 445166
rect 194317 445163 194383 445166
rect 208025 445163 208091 445166
rect 192937 445090 193003 445093
rect 209313 445090 209379 445093
rect 192937 445088 209379 445090
rect 192937 445032 192942 445088
rect 192998 445032 209318 445088
rect 209374 445032 209379 445088
rect 192937 445030 209379 445032
rect 192937 445027 193003 445030
rect 209313 445027 209379 445030
rect 307385 445090 307451 445093
rect 406469 445090 406535 445093
rect 307385 445088 406535 445090
rect 307385 445032 307390 445088
rect 307446 445032 406474 445088
rect 406530 445032 406535 445088
rect 307385 445030 406535 445032
rect 307385 445027 307451 445030
rect 406469 445027 406535 445030
rect 181437 444954 181503 444957
rect 431861 444954 431927 444957
rect 181437 444952 431927 444954
rect 181437 444896 181442 444952
rect 181498 444896 431866 444952
rect 431922 444896 431927 444952
rect 181437 444894 431927 444896
rect 181437 444891 181503 444894
rect 431861 444891 431927 444894
rect 583520 444668 584960 444908
rect 248321 439514 248387 439517
rect 338062 439514 338068 439516
rect 248321 439512 338068 439514
rect 248321 439456 248326 439512
rect 248382 439456 338068 439512
rect 248321 439454 338068 439456
rect 248321 439451 248387 439454
rect 338062 439452 338068 439454
rect 338132 439452 338138 439516
rect 174486 438092 174492 438156
rect 174556 438154 174562 438156
rect 443177 438154 443243 438157
rect 174556 438152 443243 438154
rect 174556 438096 443182 438152
rect 443238 438096 443243 438152
rect 174556 438094 443243 438096
rect 174556 438092 174562 438094
rect 443177 438091 443243 438094
rect -960 436508 480 436748
rect 196566 432516 196572 432580
rect 196636 432578 196642 432580
rect 453205 432578 453271 432581
rect 196636 432576 453271 432578
rect 196636 432520 453210 432576
rect 453266 432520 453271 432576
rect 196636 432518 453271 432520
rect 196636 432516 196642 432518
rect 453205 432515 453271 432518
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect 341609 428092 341675 428093
rect 341558 428090 341564 428092
rect 341518 428030 341564 428090
rect 341628 428088 341675 428092
rect 341670 428032 341675 428088
rect 341558 428028 341564 428030
rect 341628 428028 341675 428032
rect 341609 428027 341675 428028
rect 170622 427620 170628 427684
rect 170692 427682 170698 427684
rect 172789 427682 172855 427685
rect 173709 427682 173775 427685
rect 170692 427680 173775 427682
rect 170692 427624 172794 427680
rect 172850 427624 173714 427680
rect 173770 427624 173775 427680
rect 170692 427622 173775 427624
rect 170692 427620 170698 427622
rect 172789 427619 172855 427622
rect 173709 427619 173775 427622
rect 199285 425778 199351 425781
rect 338430 425778 338436 425780
rect 199285 425776 338436 425778
rect 199285 425720 199290 425776
rect 199346 425720 338436 425776
rect 199285 425718 338436 425720
rect 199285 425715 199351 425718
rect 338430 425716 338436 425718
rect 338500 425716 338506 425780
rect 166942 425580 166948 425644
rect 167012 425642 167018 425644
rect 441613 425642 441679 425645
rect 167012 425640 441679 425642
rect 167012 425584 441618 425640
rect 441674 425584 441679 425640
rect 167012 425582 441679 425584
rect 167012 425580 167018 425582
rect 441613 425579 441679 425582
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 168189 423602 168255 423605
rect 170121 423604 170187 423605
rect 170070 423602 170076 423604
rect 168189 423600 170076 423602
rect 170140 423602 170187 423604
rect 170140 423600 170232 423602
rect 168189 423544 168194 423600
rect 168250 423544 170076 423600
rect 170182 423544 170232 423600
rect 168189 423542 170076 423544
rect 168189 423539 168255 423542
rect 170070 423540 170076 423542
rect 170140 423542 170232 423544
rect 170140 423540 170187 423542
rect 170121 423539 170187 423540
rect 198774 422860 198780 422924
rect 198844 422922 198850 422924
rect 549253 422922 549319 422925
rect 198844 422920 549319 422922
rect 198844 422864 549258 422920
rect 549314 422864 549319 422920
rect 198844 422862 549319 422864
rect 198844 422860 198850 422862
rect 549253 422859 549319 422862
rect 337142 421772 337148 421836
rect 337212 421834 337218 421836
rect 337377 421834 337443 421837
rect 337212 421832 337443 421834
rect 337212 421776 337382 421832
rect 337438 421776 337443 421832
rect 337212 421774 337443 421776
rect 337212 421772 337218 421774
rect 337377 421771 337443 421774
rect 338849 421834 338915 421837
rect 340045 421836 340111 421837
rect 338982 421834 338988 421836
rect 338849 421832 338988 421834
rect 338849 421776 338854 421832
rect 338910 421776 338988 421832
rect 338849 421774 338988 421776
rect 338849 421771 338915 421774
rect 338982 421772 338988 421774
rect 339052 421772 339058 421836
rect 340045 421832 340092 421836
rect 340156 421834 340162 421836
rect 340045 421776 340050 421832
rect 340045 421772 340092 421776
rect 340156 421774 340202 421834
rect 340156 421772 340162 421774
rect 340045 421771 340111 421772
rect 197813 421698 197879 421701
rect 390093 421698 390159 421701
rect 197813 421696 390159 421698
rect 197813 421640 197818 421696
rect 197874 421640 390098 421696
rect 390154 421640 390159 421696
rect 197813 421638 390159 421640
rect 197813 421635 197879 421638
rect 390093 421635 390159 421638
rect 200113 421562 200179 421565
rect 396349 421562 396415 421565
rect 200113 421560 396415 421562
rect 200113 421504 200118 421560
rect 200174 421504 396354 421560
rect 396410 421504 396415 421560
rect 200113 421502 396415 421504
rect 200113 421499 200179 421502
rect 396349 421499 396415 421502
rect 196709 421426 196775 421429
rect 395061 421426 395127 421429
rect 196709 421424 395127 421426
rect 196709 421368 196714 421424
rect 196770 421368 395066 421424
rect 395122 421368 395127 421424
rect 196709 421366 395127 421368
rect 196709 421363 196775 421366
rect 395061 421363 395127 421366
rect 171542 421228 171548 421292
rect 171612 421290 171618 421292
rect 401593 421290 401659 421293
rect 171612 421288 401659 421290
rect 171612 421232 401598 421288
rect 401654 421232 401659 421288
rect 171612 421230 401659 421232
rect 171612 421228 171618 421230
rect 401593 421227 401659 421230
rect 170254 421092 170260 421156
rect 170324 421154 170330 421156
rect 405181 421154 405247 421157
rect 170324 421152 405247 421154
rect 170324 421096 405186 421152
rect 405242 421096 405247 421152
rect 170324 421094 405247 421096
rect 170324 421092 170330 421094
rect 405181 421091 405247 421094
rect 167678 420956 167684 421020
rect 167748 421018 167754 421020
rect 168598 421018 168604 421020
rect 167748 420958 168604 421018
rect 167748 420956 167754 420958
rect 168598 420956 168604 420958
rect 168668 420956 168674 421020
rect 174670 420956 174676 421020
rect 174740 421018 174746 421020
rect 411437 421018 411503 421021
rect 174740 421016 411503 421018
rect 174740 420960 411442 421016
rect 411498 420960 411503 421016
rect 174740 420958 411503 420960
rect 174740 420956 174746 420958
rect 411437 420955 411503 420958
rect 174486 419596 174492 419660
rect 174556 419658 174562 419660
rect 391381 419658 391447 419661
rect 174556 419656 391447 419658
rect 174556 419600 391386 419656
rect 391442 419600 391447 419656
rect 174556 419598 391447 419600
rect 174556 419596 174562 419598
rect 391381 419595 391447 419598
rect 197353 419114 197419 419117
rect 197353 419112 200130 419114
rect 197353 419056 197358 419112
rect 197414 419056 200130 419112
rect 197353 419054 200130 419056
rect 197353 419051 197419 419054
rect 200070 418472 200130 419054
rect 580349 418298 580415 418301
rect 583520 418298 584960 418388
rect 580349 418296 584960 418298
rect 580349 418240 580354 418296
rect 580410 418240 584960 418296
rect 580349 418238 584960 418240
rect 580349 418235 580415 418238
rect 583520 418148 584960 418238
rect 196893 417210 196959 417213
rect 196893 417208 200032 417210
rect 196893 417152 196898 417208
rect 196954 417152 200032 417208
rect 196893 417150 200032 417152
rect 196893 417147 196959 417150
rect 197353 416666 197419 416669
rect 197353 416664 200130 416666
rect 197353 416608 197358 416664
rect 197414 416608 200130 416664
rect 197353 416606 200130 416608
rect 197353 416603 197419 416606
rect 200070 416024 200130 416606
rect 560201 415170 560267 415173
rect 556876 415168 560267 415170
rect 556876 415112 560206 415168
rect 560262 415112 560267 415168
rect 556876 415110 560267 415112
rect 560201 415107 560267 415110
rect 197353 415034 197419 415037
rect 197353 415032 200130 415034
rect 197353 414976 197358 415032
rect 197414 414976 200130 415032
rect 197353 414974 200130 414976
rect 197353 414971 197419 414974
rect 200070 414800 200130 414974
rect 197353 413538 197419 413541
rect 197353 413536 200032 413538
rect 197353 413480 197358 413536
rect 197414 413480 200032 413536
rect 197353 413478 200032 413480
rect 197353 413475 197419 413478
rect 197353 412314 197419 412317
rect 197353 412312 200032 412314
rect 197353 412256 197358 412312
rect 197414 412256 200032 412312
rect 197353 412254 200032 412256
rect 197353 412251 197419 412254
rect 197353 411090 197419 411093
rect 197353 411088 200032 411090
rect 197353 411032 197358 411088
rect 197414 411032 200032 411088
rect 197353 411030 200032 411032
rect 197353 411027 197419 411030
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 197353 409866 197419 409869
rect 197353 409864 200032 409866
rect 197353 409808 197358 409864
rect 197414 409808 200032 409864
rect 197353 409806 200032 409808
rect 197353 409803 197419 409806
rect 197445 408642 197511 408645
rect 197445 408640 200032 408642
rect 197445 408584 197450 408640
rect 197506 408584 200032 408640
rect 197445 408582 200032 408584
rect 197445 408579 197511 408582
rect 197353 407962 197419 407965
rect 197353 407960 200130 407962
rect 197353 407904 197358 407960
rect 197414 407904 200130 407960
rect 197353 407902 200130 407904
rect 197353 407899 197419 407902
rect 200070 407320 200130 407902
rect 560109 407146 560175 407149
rect 556876 407144 560175 407146
rect 556876 407088 560114 407144
rect 560170 407088 560175 407144
rect 556876 407086 560175 407088
rect 560109 407083 560175 407086
rect 197721 406058 197787 406061
rect 197721 406056 200032 406058
rect 197721 406000 197726 406056
rect 197782 406000 200032 406056
rect 197721 405998 200032 406000
rect 197721 405995 197787 405998
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 197353 404834 197419 404837
rect 197353 404832 200032 404834
rect 197353 404776 197358 404832
rect 197414 404776 200032 404832
rect 583520 404820 584960 404910
rect 197353 404774 200032 404776
rect 197353 404771 197419 404774
rect 197353 403610 197419 403613
rect 197353 403608 200032 403610
rect 197353 403552 197358 403608
rect 197414 403552 200032 403608
rect 197353 403550 200032 403552
rect 197353 403547 197419 403550
rect 168373 402930 168439 402933
rect 167134 402928 168439 402930
rect 167134 402924 168378 402928
rect 166612 402872 168378 402924
rect 168434 402872 168439 402928
rect 166612 402870 168439 402872
rect 166612 402864 167194 402870
rect 168373 402867 168439 402870
rect 196801 402386 196867 402389
rect 196801 402384 200032 402386
rect 196801 402328 196806 402384
rect 196862 402328 200032 402384
rect 196801 402326 200032 402328
rect 196801 402323 196867 402326
rect 169569 401978 169635 401981
rect 167134 401976 169635 401978
rect 167134 401972 169574 401976
rect 166612 401920 169574 401972
rect 169630 401920 169635 401976
rect 166612 401918 169635 401920
rect 166612 401912 167194 401918
rect 169569 401915 169635 401918
rect 168373 401706 168439 401709
rect 168925 401706 168991 401709
rect 168373 401704 168991 401706
rect 168373 401648 168378 401704
rect 168434 401648 168930 401704
rect 168986 401648 168991 401704
rect 168373 401646 168991 401648
rect 168373 401643 168439 401646
rect 168925 401643 168991 401646
rect 197353 401162 197419 401165
rect 197353 401160 200032 401162
rect 197353 401104 197358 401160
rect 197414 401104 200032 401160
rect 197353 401102 200032 401104
rect 197353 401099 197419 401102
rect 197353 399938 197419 399941
rect 197353 399936 200100 399938
rect 197353 399880 197358 399936
rect 197414 399880 200100 399936
rect 197353 399878 200100 399880
rect 197353 399875 197419 399878
rect 168465 399802 168531 399805
rect 168741 399802 168807 399805
rect 167134 399800 168807 399802
rect 167134 399796 168470 399800
rect 166612 399744 168470 399796
rect 168526 399744 168746 399800
rect 168802 399744 168807 399800
rect 166612 399742 168807 399744
rect 166612 399736 167194 399742
rect 168465 399739 168531 399742
rect 168741 399739 168807 399742
rect 560017 399122 560083 399125
rect 556876 399120 560083 399122
rect 556876 399064 560022 399120
rect 560078 399064 560083 399120
rect 556876 399062 560083 399064
rect 560017 399059 560083 399062
rect 168649 398850 168715 398853
rect 169661 398850 169727 398853
rect 166558 398848 169727 398850
rect 166558 398792 168654 398848
rect 168710 398792 169666 398848
rect 169722 398792 169727 398848
rect 166558 398790 169727 398792
rect 168649 398787 168715 398790
rect 169661 398787 169727 398790
rect 197353 398714 197419 398717
rect 197353 398712 200100 398714
rect 197353 398656 197358 398712
rect 197414 398656 200100 398712
rect 197353 398654 200100 398656
rect 197353 398651 197419 398654
rect -960 397490 480 397580
rect 3233 397490 3299 397493
rect -960 397488 3299 397490
rect -960 397432 3238 397488
rect 3294 397432 3299 397488
rect -960 397430 3299 397432
rect -960 397340 480 397430
rect 3233 397427 3299 397430
rect 197445 397490 197511 397493
rect 197445 397488 200032 397490
rect 197445 397432 197450 397488
rect 197506 397432 200032 397488
rect 197445 397430 200032 397432
rect 197445 397427 197511 397430
rect 168649 397082 168715 397085
rect 169477 397082 169543 397085
rect 167134 397080 169543 397082
rect 167134 397076 168654 397080
rect 166612 397024 168654 397076
rect 168710 397024 169482 397080
rect 169538 397024 169543 397080
rect 166612 397022 169543 397024
rect 166612 397016 167194 397022
rect 168649 397019 168715 397022
rect 169477 397019 169543 397022
rect 197353 396130 197419 396133
rect 197353 396128 200032 396130
rect 197353 396072 197358 396128
rect 197414 396072 200032 396128
rect 197353 396070 200032 396072
rect 197353 396067 197419 396070
rect 168833 395994 168899 395997
rect 169017 395994 169083 395997
rect 167134 395992 169083 395994
rect 167134 395988 168838 395992
rect 166612 395936 168838 395988
rect 168894 395936 169022 395992
rect 169078 395936 169083 395992
rect 166612 395934 169083 395936
rect 166612 395928 167194 395934
rect 168833 395931 168899 395934
rect 169017 395931 169083 395934
rect 197353 394906 197419 394909
rect 197353 394904 200032 394906
rect 197353 394848 197358 394904
rect 197414 394848 200032 394904
rect 197353 394846 200032 394848
rect 197353 394843 197419 394846
rect 169477 394226 169543 394229
rect 167134 394224 169543 394226
rect 167134 394220 169482 394224
rect 166612 394168 169482 394220
rect 169538 394168 169543 394224
rect 166612 394166 169543 394168
rect 166612 394160 167194 394166
rect 169477 394163 169543 394166
rect 197353 393682 197419 393685
rect 197353 393680 200032 393682
rect 197353 393624 197358 393680
rect 197414 393624 200032 393680
rect 197353 393622 200032 393624
rect 197353 393619 197419 393622
rect 197353 392458 197419 392461
rect 197353 392456 200032 392458
rect 197353 392400 197358 392456
rect 197414 392400 200032 392456
rect 197353 392398 200032 392400
rect 197353 392395 197419 392398
rect 583520 391628 584960 391868
rect 197353 391234 197419 391237
rect 560201 391234 560267 391237
rect 197353 391232 200032 391234
rect 197353 391176 197358 391232
rect 197414 391176 200032 391232
rect 197353 391174 200032 391176
rect 556876 391232 560267 391234
rect 556876 391176 560206 391232
rect 560262 391176 560267 391232
rect 556876 391174 560267 391176
rect 197353 391171 197419 391174
rect 560201 391171 560267 391174
rect 197353 390010 197419 390013
rect 197353 390008 200032 390010
rect 197353 389952 197358 390008
rect 197414 389952 200032 390008
rect 197353 389950 200032 389952
rect 197353 389947 197419 389950
rect 197353 388786 197419 388789
rect 197353 388784 200032 388786
rect 197353 388728 197358 388784
rect 197414 388728 200032 388784
rect 197353 388726 200032 388728
rect 197353 388723 197419 388726
rect 197353 387562 197419 387565
rect 197353 387560 200032 387562
rect 197353 387504 197358 387560
rect 197414 387504 200032 387560
rect 197353 387502 200032 387504
rect 197353 387499 197419 387502
rect 27153 386338 27219 386341
rect 27429 386338 27495 386341
rect 27153 386336 27495 386338
rect 27153 386280 27158 386336
rect 27214 386280 27434 386336
rect 27490 386280 27495 386336
rect 27153 386278 27495 386280
rect 27153 386275 27219 386278
rect 27429 386275 27495 386278
rect 197353 386338 197419 386341
rect 197353 386336 200032 386338
rect 197353 386280 197358 386336
rect 197414 386280 200032 386336
rect 197353 386278 200032 386280
rect 197353 386275 197419 386278
rect 27153 385386 27219 385389
rect 27153 385384 30062 385386
rect 27153 385328 27158 385384
rect 27214 385328 30062 385384
rect 27153 385326 30062 385328
rect 27153 385323 27219 385326
rect 197721 385114 197787 385117
rect 197721 385112 200032 385114
rect 197721 385056 197726 385112
rect 197782 385056 200032 385112
rect 197721 385054 200032 385056
rect 197721 385051 197787 385054
rect -960 384284 480 384524
rect 197353 384434 197419 384437
rect 197353 384432 200130 384434
rect 197353 384376 197358 384432
rect 197414 384376 200130 384432
rect 197353 384374 200130 384376
rect 197353 384371 197419 384374
rect 200070 383792 200130 384374
rect 27337 383754 27403 383757
rect 27337 383752 30062 383754
rect 27337 383696 27342 383752
rect 27398 383696 30062 383752
rect 27337 383694 30062 383696
rect 27337 383691 27403 383694
rect 197353 383210 197419 383213
rect 559189 383210 559255 383213
rect 197353 383208 200130 383210
rect 197353 383152 197358 383208
rect 197414 383152 200130 383208
rect 197353 383150 200130 383152
rect 556876 383208 559255 383210
rect 556876 383152 559194 383208
rect 559250 383152 559255 383208
rect 556876 383150 559255 383152
rect 197353 383147 197419 383150
rect 200070 382568 200130 383150
rect 559189 383147 559255 383150
rect 27061 382394 27127 382397
rect 27429 382394 27495 382397
rect 167729 382394 167795 382397
rect 168414 382394 168420 382396
rect 27061 382392 30062 382394
rect 27061 382336 27066 382392
rect 27122 382336 27434 382392
rect 27490 382336 30062 382392
rect 27061 382334 30062 382336
rect 167729 382392 168420 382394
rect 167729 382336 167734 382392
rect 167790 382336 168420 382392
rect 167729 382334 168420 382336
rect 27061 382331 27127 382334
rect 27429 382331 27495 382334
rect 167729 382331 167795 382334
rect 168414 382332 168420 382334
rect 168484 382332 168490 382396
rect 197353 381306 197419 381309
rect 197353 381304 200032 381306
rect 197353 381248 197358 381304
rect 197414 381248 200032 381304
rect 197353 381246 200032 381248
rect 197353 381243 197419 381246
rect 27521 380898 27587 380901
rect 27521 380896 30062 380898
rect 27521 380840 27526 380896
rect 27582 380840 30062 380896
rect 27521 380838 30062 380840
rect 27521 380835 27587 380838
rect 197353 380082 197419 380085
rect 197353 380080 200032 380082
rect 197353 380024 197358 380080
rect 197414 380024 200032 380080
rect 197353 380022 200032 380024
rect 197353 380019 197419 380022
rect 27061 379810 27127 379813
rect 27521 379810 27587 379813
rect 27061 379808 27587 379810
rect 27061 379752 27066 379808
rect 27122 379752 27526 379808
rect 27582 379752 27587 379808
rect 27061 379750 27587 379752
rect 27061 379747 27127 379750
rect 27521 379747 27587 379750
rect 27245 379674 27311 379677
rect 27521 379674 27587 379677
rect 27245 379672 30062 379674
rect 27245 379616 27250 379672
rect 27306 379616 27526 379672
rect 27582 379616 30062 379672
rect 27245 379614 30062 379616
rect 27245 379611 27311 379614
rect 27521 379611 27587 379614
rect 168230 379476 168236 379540
rect 168300 379538 168306 379540
rect 169201 379538 169267 379541
rect 168300 379536 169267 379538
rect 168300 379480 169206 379536
rect 169262 379480 169267 379536
rect 168300 379478 169267 379480
rect 168300 379476 168306 379478
rect 169201 379475 169267 379478
rect 197353 378858 197419 378861
rect 197353 378856 200032 378858
rect 197353 378800 197358 378856
rect 197414 378800 200032 378856
rect 197353 378798 200032 378800
rect 197353 378795 197419 378798
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 197353 377634 197419 377637
rect 197353 377632 200032 377634
rect 197353 377576 197358 377632
rect 197414 377576 200032 377632
rect 197353 377574 200032 377576
rect 197353 377571 197419 377574
rect 197353 376410 197419 376413
rect 197353 376408 200032 376410
rect 197353 376352 197358 376408
rect 197414 376352 200032 376408
rect 197353 376350 200032 376352
rect 197353 376347 197419 376350
rect 169385 376002 169451 376005
rect 167134 376000 169451 376002
rect 167134 375996 169390 376000
rect 166612 375944 169390 375996
rect 169446 375944 169451 376000
rect 166612 375942 169451 375944
rect 166612 375936 167194 375942
rect 169385 375939 169451 375942
rect 168373 375322 168439 375325
rect 169293 375322 169359 375325
rect 168373 375320 169359 375322
rect 168373 375264 168378 375320
rect 168434 375264 169298 375320
rect 169354 375264 169359 375320
rect 168373 375262 169359 375264
rect 168373 375259 168439 375262
rect 169293 375259 169359 375262
rect 197353 375186 197419 375189
rect 560201 375186 560267 375189
rect 197353 375184 200032 375186
rect 197353 375128 197358 375184
rect 197414 375128 200032 375184
rect 197353 375126 200032 375128
rect 556876 375184 560267 375186
rect 556876 375128 560206 375184
rect 560262 375128 560267 375184
rect 556876 375126 560267 375128
rect 197353 375123 197419 375126
rect 560201 375123 560267 375126
rect 168373 374370 168439 374373
rect 167134 374368 168439 374370
rect 167134 374364 168378 374368
rect 166612 374312 168378 374364
rect 168434 374312 168439 374368
rect 166612 374310 168439 374312
rect 166612 374304 167194 374310
rect 168373 374307 168439 374310
rect 168557 374098 168623 374101
rect 167134 374096 168623 374098
rect 167134 374092 168562 374096
rect 166612 374040 168562 374092
rect 168618 374040 168623 374096
rect 166612 374038 168623 374040
rect 166612 374032 167194 374038
rect 168557 374035 168623 374038
rect 197353 373962 197419 373965
rect 197353 373960 200032 373962
rect 197353 373904 197358 373960
rect 197414 373904 200032 373960
rect 197353 373902 200032 373904
rect 197353 373899 197419 373902
rect 197353 372602 197419 372605
rect 197353 372600 200032 372602
rect 197353 372544 197358 372600
rect 197414 372544 200032 372600
rect 197353 372542 200032 372544
rect 197353 372539 197419 372542
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 197445 371378 197511 371381
rect 197445 371376 200032 371378
rect 197445 371320 197450 371376
rect 197506 371320 200032 371376
rect 197445 371318 200032 371320
rect 197445 371315 197511 371318
rect 197353 370154 197419 370157
rect 197353 370152 200032 370154
rect 197353 370096 197358 370152
rect 197414 370096 200032 370152
rect 197353 370094 200032 370096
rect 197353 370091 197419 370094
rect 197353 368930 197419 368933
rect 197353 368928 200032 368930
rect 197353 368872 197358 368928
rect 197414 368872 200032 368928
rect 197353 368870 200032 368872
rect 197353 368867 197419 368870
rect 197353 368386 197419 368389
rect 197353 368384 200130 368386
rect 197353 368328 197358 368384
rect 197414 368328 200130 368384
rect 197353 368326 200130 368328
rect 197353 368323 197419 368326
rect 200070 367744 200130 368326
rect 559189 367298 559255 367301
rect 556876 367296 559255 367298
rect 556876 367240 559194 367296
rect 559250 367240 559255 367296
rect 556876 367238 559255 367240
rect 559189 367235 559255 367238
rect 197353 367026 197419 367029
rect 197353 367024 200130 367026
rect 197353 366968 197358 367024
rect 197414 366968 200130 367024
rect 197353 366966 200130 366968
rect 197353 366963 197419 366966
rect 200070 366520 200130 366966
rect 197353 365258 197419 365261
rect 197353 365256 200032 365258
rect 197353 365200 197358 365256
rect 197414 365200 200032 365256
rect 197353 365198 200032 365200
rect 197353 365195 197419 365198
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect 42885 364306 42951 364309
rect 43110 364306 43116 364308
rect 42885 364304 43116 364306
rect 42885 364248 42890 364304
rect 42946 364248 43116 364304
rect 42885 364246 43116 364248
rect 42885 364243 42951 364246
rect 43110 364244 43116 364246
rect 43180 364244 43186 364308
rect 112110 364244 112116 364308
rect 112180 364306 112186 364308
rect 112989 364306 113055 364309
rect 112180 364304 113055 364306
rect 112180 364248 112994 364304
rect 113050 364248 113055 364304
rect 112180 364246 113055 364248
rect 112180 364244 112186 364246
rect 112989 364243 113055 364246
rect 115422 364244 115428 364308
rect 115492 364306 115498 364308
rect 115749 364306 115815 364309
rect 132953 364308 133019 364309
rect 132902 364306 132908 364308
rect 115492 364304 115815 364306
rect 115492 364248 115754 364304
rect 115810 364248 115815 364304
rect 115492 364246 115815 364248
rect 132862 364246 132908 364306
rect 132972 364304 133019 364308
rect 133014 364248 133019 364304
rect 115492 364244 115498 364246
rect 115749 364243 115815 364246
rect 132902 364244 132908 364246
rect 132972 364244 133019 364248
rect 135294 364244 135300 364308
rect 135364 364306 135370 364308
rect 136541 364306 136607 364309
rect 135364 364304 136607 364306
rect 135364 364248 136546 364304
rect 136602 364248 136607 364304
rect 135364 364246 136607 364248
rect 135364 364244 135370 364246
rect 132953 364243 133019 364244
rect 136541 364243 136607 364246
rect 143349 364308 143415 364309
rect 143349 364304 143396 364308
rect 143460 364306 143466 364308
rect 143349 364248 143354 364304
rect 143349 364244 143396 364248
rect 143460 364246 143506 364306
rect 143460 364244 143466 364246
rect 144678 364244 144684 364308
rect 144748 364306 144754 364308
rect 145966 364306 145972 364308
rect 144748 364246 145972 364306
rect 144748 364244 144754 364246
rect 145966 364244 145972 364246
rect 146036 364244 146042 364308
rect 143349 364243 143415 364244
rect 42793 364170 42859 364173
rect 43478 364170 43484 364172
rect 42793 364168 43484 364170
rect 42793 364112 42798 364168
rect 42854 364112 43484 364168
rect 42793 364110 43484 364112
rect 42793 364107 42859 364110
rect 43478 364108 43484 364110
rect 43548 364108 43554 364172
rect 63166 364108 63172 364172
rect 63236 364170 63242 364172
rect 63401 364170 63467 364173
rect 63236 364168 63467 364170
rect 63236 364112 63406 364168
rect 63462 364112 63467 364168
rect 63236 364110 63467 364112
rect 63236 364108 63242 364110
rect 63401 364107 63467 364110
rect 65742 364108 65748 364172
rect 65812 364170 65818 364172
rect 66161 364170 66227 364173
rect 73153 364172 73219 364173
rect 73102 364170 73108 364172
rect 65812 364168 66227 364170
rect 65812 364112 66166 364168
rect 66222 364112 66227 364168
rect 65812 364110 66227 364112
rect 73062 364110 73108 364170
rect 73172 364168 73219 364172
rect 73214 364112 73219 364168
rect 65812 364108 65818 364110
rect 66161 364107 66227 364110
rect 73102 364108 73108 364110
rect 73172 364108 73219 364112
rect 75678 364108 75684 364172
rect 75748 364170 75754 364172
rect 75821 364170 75887 364173
rect 75748 364168 75887 364170
rect 75748 364112 75826 364168
rect 75882 364112 75887 364168
rect 75748 364110 75887 364112
rect 75748 364108 75754 364110
rect 73153 364107 73219 364108
rect 75821 364107 75887 364110
rect 83038 364108 83044 364172
rect 83108 364170 83114 364172
rect 84101 364170 84167 364173
rect 85665 364172 85731 364173
rect 85614 364170 85620 364172
rect 83108 364168 84167 364170
rect 83108 364112 84106 364168
rect 84162 364112 84167 364168
rect 83108 364110 84167 364112
rect 85574 364110 85620 364170
rect 85684 364168 85731 364172
rect 85726 364112 85731 364168
rect 83108 364108 83114 364110
rect 84101 364107 84167 364110
rect 85614 364108 85620 364110
rect 85684 364108 85731 364112
rect 93158 364108 93164 364172
rect 93228 364170 93234 364172
rect 93761 364170 93827 364173
rect 95601 364172 95667 364173
rect 103145 364172 103211 364173
rect 95550 364170 95556 364172
rect 93228 364168 93827 364170
rect 93228 364112 93766 364168
rect 93822 364112 93827 364168
rect 93228 364110 93827 364112
rect 95510 364110 95556 364170
rect 95620 364168 95667 364172
rect 103094 364170 103100 364172
rect 95662 364112 95667 364168
rect 93228 364108 93234 364110
rect 85665 364107 85731 364108
rect 93761 364107 93827 364110
rect 95550 364108 95556 364110
rect 95620 364108 95667 364112
rect 103054 364110 103100 364170
rect 103164 364168 103211 364172
rect 103206 364112 103211 364168
rect 103094 364108 103100 364110
rect 103164 364108 103211 364112
rect 105670 364108 105676 364172
rect 105740 364170 105746 364172
rect 106181 364170 106247 364173
rect 109585 364172 109651 364173
rect 113081 364172 113147 364173
rect 109534 364170 109540 364172
rect 105740 364168 106247 364170
rect 105740 364112 106186 364168
rect 106242 364112 106247 364168
rect 105740 364110 106247 364112
rect 109494 364110 109540 364170
rect 109604 364168 109651 364172
rect 113030 364170 113036 364172
rect 109646 364112 109651 364168
rect 105740 364108 105746 364110
rect 95601 364107 95667 364108
rect 103145 364107 103211 364108
rect 106181 364107 106247 364110
rect 109534 364108 109540 364110
rect 109604 364108 109651 364112
rect 112990 364110 113036 364170
rect 113100 364168 113147 364172
rect 113142 364112 113147 364168
rect 113030 364108 113036 364110
rect 113100 364108 113147 364112
rect 113214 364108 113220 364172
rect 113284 364170 113290 364172
rect 114461 364170 114527 364173
rect 113284 364168 114527 364170
rect 113284 364112 114466 364168
rect 114522 364112 114527 364168
rect 113284 364110 114527 364112
rect 113284 364108 113290 364110
rect 109585 364107 109651 364108
rect 113081 364107 113147 364108
rect 114461 364107 114527 364110
rect 115606 364108 115612 364172
rect 115676 364170 115682 364172
rect 115841 364170 115907 364173
rect 115676 364168 115907 364170
rect 115676 364112 115846 364168
rect 115902 364112 115907 364168
rect 115676 364110 115907 364112
rect 115676 364108 115682 364110
rect 115841 364107 115907 364110
rect 122966 364108 122972 364172
rect 123036 364170 123042 364172
rect 124029 364170 124095 364173
rect 125961 364172 126027 364173
rect 125910 364170 125916 364172
rect 123036 364168 124095 364170
rect 123036 364112 124034 364168
rect 124090 364112 124095 364168
rect 123036 364110 124095 364112
rect 125870 364110 125916 364170
rect 125980 364168 126027 364172
rect 126022 364112 126027 364168
rect 123036 364108 123042 364110
rect 124029 364107 124095 364110
rect 125910 364108 125916 364110
rect 125980 364108 126027 364112
rect 125961 364107 126027 364108
rect 129549 364172 129615 364173
rect 132033 364172 132099 364173
rect 133137 364172 133203 364173
rect 135897 364172 135963 364173
rect 129549 364168 129596 364172
rect 129660 364170 129666 364172
rect 131982 364170 131988 364172
rect 129549 364112 129554 364168
rect 129549 364108 129596 364112
rect 129660 364110 129706 364170
rect 131942 364110 131988 364170
rect 132052 364168 132099 364172
rect 133086 364170 133092 364172
rect 132094 364112 132099 364168
rect 129660 364108 129666 364110
rect 131982 364108 131988 364110
rect 132052 364108 132099 364112
rect 133046 364110 133092 364170
rect 133156 364168 133203 364172
rect 135846 364170 135852 364172
rect 133198 364112 133203 364168
rect 133086 364108 133092 364110
rect 133156 364108 133203 364112
rect 135806 364110 135852 364170
rect 135916 364168 135963 364172
rect 135958 364112 135963 364168
rect 135846 364108 135852 364110
rect 135916 364108 135963 364112
rect 142286 364108 142292 364172
rect 142356 364170 142362 364172
rect 143441 364170 143507 364173
rect 142356 364168 143507 364170
rect 142356 364112 143446 364168
rect 143502 364112 143507 364168
rect 142356 364110 143507 364112
rect 142356 364108 142362 364110
rect 129549 364107 129658 364108
rect 132033 364107 132099 364108
rect 133137 364107 133203 364108
rect 135897 364107 135963 364108
rect 143441 364107 143507 364110
rect 149462 364108 149468 364172
rect 149532 364170 149538 364172
rect 150341 364170 150407 364173
rect 167177 364172 167243 364173
rect 149532 364168 150407 364170
rect 149532 364112 150346 364168
rect 150402 364112 150407 364168
rect 149532 364110 150407 364112
rect 149532 364108 149538 364110
rect 150341 364107 150407 364110
rect 167126 364108 167132 364172
rect 167196 364170 167243 364172
rect 167196 364168 167288 364170
rect 167238 364112 167288 364168
rect 167196 364110 167288 364112
rect 167196 364108 167243 364110
rect 167177 364107 167243 364108
rect 120206 363972 120212 364036
rect 120276 364034 120282 364036
rect 127617 364034 127683 364037
rect 120276 364032 127683 364034
rect 120276 363976 127622 364032
rect 127678 363976 127683 364032
rect 120276 363974 127683 363976
rect 129598 364034 129658 364107
rect 170622 364034 170628 364036
rect 129598 363974 170628 364034
rect 120276 363972 120282 363974
rect 127617 363971 127683 363974
rect 170622 363972 170628 363974
rect 170692 363972 170698 364036
rect 197353 364034 197419 364037
rect 197353 364032 200032 364034
rect 197353 363976 197358 364032
rect 197414 363976 200032 364032
rect 197353 363974 200032 363976
rect 197353 363971 197419 363974
rect 122598 363836 122604 363900
rect 122668 363898 122674 363900
rect 122741 363898 122807 363901
rect 122668 363896 122807 363898
rect 122668 363840 122746 363896
rect 122802 363840 122807 363896
rect 122668 363838 122807 363840
rect 122668 363836 122674 363838
rect 122741 363835 122807 363838
rect 136541 363900 136607 363901
rect 136541 363896 136588 363900
rect 136652 363898 136658 363900
rect 166942 363898 166948 363900
rect 136541 363840 136546 363896
rect 136541 363836 136588 363840
rect 136652 363838 136698 363898
rect 142110 363838 166948 363898
rect 136652 363836 136658 363838
rect 136541 363835 136607 363836
rect 127198 363700 127204 363764
rect 127268 363762 127274 363764
rect 128261 363762 128327 363765
rect 127268 363760 128327 363762
rect 127268 363704 128266 363760
rect 128322 363704 128327 363760
rect 127268 363702 128327 363704
rect 127268 363700 127274 363702
rect 128261 363699 128327 363702
rect 135161 363762 135227 363765
rect 142110 363762 142170 363838
rect 166942 363836 166948 363838
rect 167012 363836 167018 363900
rect 135161 363760 142170 363762
rect 135161 363704 135166 363760
rect 135222 363704 142170 363760
rect 135161 363702 142170 363704
rect 135161 363699 135227 363702
rect 150566 363564 150572 363628
rect 150636 363626 150642 363628
rect 151169 363626 151235 363629
rect 150636 363624 151235 363626
rect 150636 363568 151174 363624
rect 151230 363568 151235 363624
rect 150636 363566 151235 363568
rect 150636 363564 150642 363566
rect 151169 363563 151235 363566
rect 123702 363428 123708 363492
rect 123772 363490 123778 363492
rect 124121 363490 124187 363493
rect 138289 363492 138355 363493
rect 138238 363490 138244 363492
rect 123772 363488 124187 363490
rect 123772 363432 124126 363488
rect 124182 363432 124187 363488
rect 123772 363430 124187 363432
rect 138198 363430 138244 363490
rect 138308 363488 138355 363492
rect 138350 363432 138355 363488
rect 123772 363428 123778 363430
rect 124121 363427 124187 363430
rect 138238 363428 138244 363430
rect 138308 363428 138355 363432
rect 138289 363427 138355 363428
rect 108062 363292 108068 363356
rect 108132 363354 108138 363356
rect 108849 363354 108915 363357
rect 108132 363352 108915 363354
rect 108132 363296 108854 363352
rect 108910 363296 108915 363352
rect 108132 363294 108915 363296
rect 108132 363292 108138 363294
rect 108849 363291 108915 363294
rect 118918 363292 118924 363356
rect 118988 363354 118994 363356
rect 119981 363354 120047 363357
rect 167126 363354 167132 363356
rect 118988 363352 167132 363354
rect 118988 363296 119986 363352
rect 120042 363296 167132 363352
rect 118988 363294 167132 363296
rect 118988 363292 118994 363294
rect 119981 363291 120047 363294
rect 167126 363292 167132 363294
rect 167196 363292 167202 363356
rect 110454 363156 110460 363220
rect 110524 363218 110530 363220
rect 111609 363218 111675 363221
rect 110524 363216 111675 363218
rect 110524 363160 111614 363216
rect 111670 363160 111675 363216
rect 110524 363158 111675 363160
rect 110524 363156 110530 363158
rect 111609 363155 111675 363158
rect 117814 363156 117820 363220
rect 117884 363218 117890 363220
rect 118509 363218 118575 363221
rect 117884 363216 118575 363218
rect 117884 363160 118514 363216
rect 118570 363160 118575 363216
rect 117884 363158 118575 363160
rect 117884 363156 117890 363158
rect 118509 363155 118575 363158
rect 120574 363156 120580 363220
rect 120644 363218 120650 363220
rect 121269 363218 121335 363221
rect 120644 363216 121335 363218
rect 120644 363160 121274 363216
rect 121330 363160 121335 363216
rect 120644 363158 121335 363160
rect 120644 363156 120650 363158
rect 121269 363155 121335 363158
rect 124806 363156 124812 363220
rect 124876 363218 124882 363220
rect 125501 363218 125567 363221
rect 124876 363216 125567 363218
rect 124876 363160 125506 363216
rect 125562 363160 125567 363216
rect 124876 363158 125567 363160
rect 124876 363156 124882 363158
rect 125501 363155 125567 363158
rect 130694 363156 130700 363220
rect 130764 363218 130770 363220
rect 130929 363218 130995 363221
rect 130764 363216 130995 363218
rect 130764 363160 130934 363216
rect 130990 363160 130995 363216
rect 130764 363158 130995 363160
rect 130764 363156 130770 363158
rect 130929 363155 130995 363158
rect 60641 363084 60707 363085
rect 60590 363082 60596 363084
rect 60550 363022 60596 363082
rect 60660 363080 60707 363084
rect 60702 363024 60707 363080
rect 60590 363020 60596 363022
rect 60660 363020 60707 363024
rect 68134 363020 68140 363084
rect 68204 363082 68210 363084
rect 68921 363082 68987 363085
rect 68204 363080 68987 363082
rect 68204 363024 68926 363080
rect 68982 363024 68987 363080
rect 68204 363022 68987 363024
rect 68204 363020 68210 363022
rect 60641 363019 60707 363020
rect 68921 363019 68987 363022
rect 70710 363020 70716 363084
rect 70780 363082 70786 363084
rect 71681 363082 71747 363085
rect 70780 363080 71747 363082
rect 70780 363024 71686 363080
rect 71742 363024 71747 363080
rect 70780 363022 71747 363024
rect 70780 363020 70786 363022
rect 71681 363019 71747 363022
rect 78070 363020 78076 363084
rect 78140 363082 78146 363084
rect 78581 363082 78647 363085
rect 78140 363080 78647 363082
rect 78140 363024 78586 363080
rect 78642 363024 78647 363080
rect 78140 363022 78647 363024
rect 78140 363020 78146 363022
rect 78581 363019 78647 363022
rect 80646 363020 80652 363084
rect 80716 363082 80722 363084
rect 81341 363082 81407 363085
rect 88241 363084 88307 363085
rect 88190 363082 88196 363084
rect 80716 363080 81407 363082
rect 80716 363024 81346 363080
rect 81402 363024 81407 363080
rect 80716 363022 81407 363024
rect 88150 363022 88196 363082
rect 88260 363080 88307 363084
rect 88302 363024 88307 363080
rect 80716 363020 80722 363022
rect 81341 363019 81407 363022
rect 88190 363020 88196 363022
rect 88260 363020 88307 363024
rect 90766 363020 90772 363084
rect 90836 363082 90842 363084
rect 91001 363082 91067 363085
rect 90836 363080 91067 363082
rect 90836 363024 91006 363080
rect 91062 363024 91067 363080
rect 90836 363022 91067 363024
rect 90836 363020 90842 363022
rect 88241 363019 88307 363020
rect 91001 363019 91067 363022
rect 98310 363020 98316 363084
rect 98380 363082 98386 363084
rect 99281 363082 99347 363085
rect 98380 363080 99347 363082
rect 98380 363024 99286 363080
rect 99342 363024 99347 363080
rect 98380 363022 99347 363024
rect 98380 363020 98386 363022
rect 99281 363019 99347 363022
rect 100518 363020 100524 363084
rect 100588 363082 100594 363084
rect 100661 363082 100727 363085
rect 100588 363080 100727 363082
rect 100588 363024 100666 363080
rect 100722 363024 100727 363080
rect 100588 363022 100727 363024
rect 100588 363020 100594 363022
rect 100661 363019 100727 363022
rect 107326 363020 107332 363084
rect 107396 363082 107402 363084
rect 107561 363082 107627 363085
rect 107396 363080 107627 363082
rect 107396 363024 107566 363080
rect 107622 363024 107627 363080
rect 107396 363022 107627 363024
rect 107396 363020 107402 363022
rect 107561 363019 107627 363022
rect 108430 363020 108436 363084
rect 108500 363082 108506 363084
rect 108941 363082 109007 363085
rect 108500 363080 109007 363082
rect 108500 363024 108946 363080
rect 109002 363024 109007 363080
rect 108500 363022 109007 363024
rect 108500 363020 108506 363022
rect 108941 363019 109007 363022
rect 110822 363020 110828 363084
rect 110892 363082 110898 363084
rect 111701 363082 111767 363085
rect 114369 363084 114435 363085
rect 114318 363082 114324 363084
rect 110892 363080 111767 363082
rect 110892 363024 111706 363080
rect 111762 363024 111767 363080
rect 110892 363022 111767 363024
rect 114278 363022 114324 363082
rect 114388 363080 114435 363084
rect 114430 363024 114435 363080
rect 110892 363020 110898 363022
rect 111701 363019 111767 363022
rect 114318 363020 114324 363022
rect 114388 363020 114435 363024
rect 116710 363020 116716 363084
rect 116780 363082 116786 363084
rect 117221 363082 117287 363085
rect 116780 363080 117287 363082
rect 116780 363024 117226 363080
rect 117282 363024 117287 363080
rect 116780 363022 117287 363024
rect 116780 363020 116786 363022
rect 114369 363019 114435 363020
rect 117221 363019 117287 363022
rect 118366 363020 118372 363084
rect 118436 363082 118442 363084
rect 118601 363082 118667 363085
rect 118436 363080 118667 363082
rect 118436 363024 118606 363080
rect 118662 363024 118667 363080
rect 118436 363022 118667 363024
rect 118436 363020 118442 363022
rect 118601 363019 118667 363022
rect 121177 363082 121243 363085
rect 125409 363084 125475 363085
rect 128169 363084 128235 363085
rect 121310 363082 121316 363084
rect 121177 363080 121316 363082
rect 121177 363024 121182 363080
rect 121238 363024 121316 363080
rect 121177 363022 121316 363024
rect 121177 363019 121243 363022
rect 121310 363020 121316 363022
rect 121380 363020 121386 363084
rect 125358 363082 125364 363084
rect 125318 363022 125364 363082
rect 125428 363080 125475 363084
rect 128118 363082 128124 363084
rect 125470 363024 125475 363080
rect 125358 363020 125364 363022
rect 125428 363020 125475 363024
rect 128078 363022 128124 363082
rect 128188 363080 128235 363084
rect 128230 363024 128235 363080
rect 128118 363020 128124 363022
rect 128188 363020 128235 363024
rect 128486 363020 128492 363084
rect 128556 363082 128562 363084
rect 129641 363082 129707 363085
rect 128556 363080 129707 363082
rect 128556 363024 129646 363080
rect 129702 363024 129707 363080
rect 128556 363022 129707 363024
rect 128556 363020 128562 363022
rect 125409 363019 125475 363020
rect 128169 363019 128235 363020
rect 129641 363019 129707 363022
rect 130510 363020 130516 363084
rect 130580 363082 130586 363084
rect 131021 363082 131087 363085
rect 130580 363080 131087 363082
rect 130580 363024 131026 363080
rect 131082 363024 131087 363080
rect 130580 363022 131087 363024
rect 130580 363020 130586 363022
rect 131021 363019 131087 363022
rect 134190 363020 134196 363084
rect 134260 363082 134266 363084
rect 135161 363082 135227 363085
rect 137921 363084 137987 363085
rect 137870 363082 137876 363084
rect 134260 363080 135227 363082
rect 134260 363024 135166 363080
rect 135222 363024 135227 363080
rect 134260 363022 135227 363024
rect 137830 363022 137876 363082
rect 137940 363080 137987 363084
rect 137982 363024 137987 363080
rect 134260 363020 134266 363022
rect 135161 363019 135227 363022
rect 137870 363020 137876 363022
rect 137940 363020 137987 363024
rect 138974 363020 138980 363084
rect 139044 363082 139050 363084
rect 139209 363082 139275 363085
rect 139044 363080 139275 363082
rect 139044 363024 139214 363080
rect 139270 363024 139275 363080
rect 139044 363022 139275 363024
rect 139044 363020 139050 363022
rect 137921 363019 137987 363020
rect 139209 363019 139275 363022
rect 140078 363020 140084 363084
rect 140148 363082 140154 363084
rect 140313 363082 140379 363085
rect 140148 363080 140379 363082
rect 140148 363024 140318 363080
rect 140374 363024 140379 363080
rect 140148 363022 140379 363024
rect 140148 363020 140154 363022
rect 140313 363019 140379 363022
rect 141182 363020 141188 363084
rect 141252 363082 141258 363084
rect 142061 363082 142127 363085
rect 141252 363080 142127 363082
rect 141252 363024 142066 363080
rect 142122 363024 142127 363080
rect 141252 363022 142127 363024
rect 141252 363020 141258 363022
rect 142061 363019 142127 363022
rect 148358 363020 148364 363084
rect 148428 363082 148434 363084
rect 148961 363082 149027 363085
rect 148428 363080 149027 363082
rect 148428 363024 148966 363080
rect 149022 363024 149027 363080
rect 148428 363022 149027 363024
rect 148428 363020 148434 363022
rect 148961 363019 149027 363022
rect 197353 362810 197419 362813
rect 197353 362808 200032 362810
rect 197353 362752 197358 362808
rect 197414 362752 200032 362808
rect 197353 362750 200032 362752
rect 197353 362747 197419 362750
rect 170438 361660 170444 361724
rect 170508 361722 170514 361724
rect 170765 361722 170831 361725
rect 170508 361720 170831 361722
rect 170508 361664 170770 361720
rect 170826 361664 170831 361720
rect 170508 361662 170831 361664
rect 170508 361660 170514 361662
rect 170765 361659 170831 361662
rect 197353 361450 197419 361453
rect 197353 361448 200032 361450
rect 197353 361392 197358 361448
rect 197414 361392 200032 361448
rect 197353 361390 200032 361392
rect 197353 361387 197419 361390
rect 197445 360226 197511 360229
rect 197445 360224 200032 360226
rect 197445 360168 197450 360224
rect 197506 360168 200032 360224
rect 197445 360166 200032 360168
rect 197445 360163 197511 360166
rect 197353 359682 197419 359685
rect 197353 359680 200130 359682
rect 197353 359624 197358 359680
rect 197414 359624 200130 359680
rect 197353 359622 200130 359624
rect 197353 359619 197419 359622
rect 200070 359040 200130 359622
rect 560201 359274 560267 359277
rect 556876 359272 560267 359274
rect 556876 359216 560206 359272
rect 560262 359216 560267 359272
rect 556876 359214 560267 359216
rect 560201 359211 560267 359214
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 197353 357778 197419 357781
rect 197353 357776 200032 357778
rect 197353 357720 197358 357776
rect 197414 357720 200032 357776
rect 197353 357718 200032 357720
rect 197353 357715 197419 357718
rect 197353 356554 197419 356557
rect 197353 356552 200032 356554
rect 197353 356496 197358 356552
rect 197414 356496 200032 356552
rect 197353 356494 200032 356496
rect 197353 356491 197419 356494
rect 197353 355330 197419 355333
rect 197353 355328 200032 355330
rect 197353 355272 197358 355328
rect 197414 355272 200032 355328
rect 197353 355270 200032 355272
rect 197353 355267 197419 355270
rect 197353 354106 197419 354109
rect 197353 354104 200032 354106
rect 197353 354048 197358 354104
rect 197414 354048 200032 354104
rect 197353 354046 200032 354048
rect 197353 354043 197419 354046
rect 107561 353290 107627 353293
rect 168598 353290 168604 353292
rect 107561 353288 168604 353290
rect 107561 353232 107566 353288
rect 107622 353232 168604 353288
rect 107561 353230 168604 353232
rect 107561 353227 107627 353230
rect 168598 353228 168604 353230
rect 168668 353228 168674 353292
rect 197353 352882 197419 352885
rect 197353 352880 200032 352882
rect 197353 352824 197358 352880
rect 197414 352824 200032 352880
rect 197353 352822 200032 352824
rect 197353 352819 197419 352822
rect 168598 352548 168604 352612
rect 168668 352610 168674 352612
rect 180149 352610 180215 352613
rect 168668 352608 180215 352610
rect 168668 352552 180154 352608
rect 180210 352552 180215 352608
rect 168668 352550 180215 352552
rect 168668 352548 168674 352550
rect 180149 352547 180215 352550
rect 578877 351930 578943 351933
rect 583520 351930 584960 352020
rect 578877 351928 584960 351930
rect 578877 351872 578882 351928
rect 578938 351872 584960 351928
rect 578877 351870 584960 351872
rect 578877 351867 578943 351870
rect 583520 351780 584960 351870
rect 197353 351658 197419 351661
rect 197353 351656 200100 351658
rect 197353 351600 197358 351656
rect 197414 351600 200100 351656
rect 197353 351598 200100 351600
rect 197353 351595 197419 351598
rect 559649 351250 559715 351253
rect 556876 351248 559715 351250
rect 556876 351192 559654 351248
rect 559710 351192 559715 351248
rect 556876 351190 559715 351192
rect 559649 351187 559715 351190
rect 197353 350434 197419 350437
rect 197353 350432 200100 350434
rect 197353 350376 197358 350432
rect 197414 350376 200100 350432
rect 197353 350374 200100 350376
rect 197353 350371 197419 350374
rect 197445 349074 197511 349077
rect 197445 349072 200032 349074
rect 197445 349016 197450 349072
rect 197506 349016 200032 349072
rect 197445 349014 200032 349016
rect 197445 349011 197511 349014
rect 197353 347850 197419 347853
rect 197353 347848 200032 347850
rect 197353 347792 197358 347848
rect 197414 347792 200032 347848
rect 197353 347790 200032 347792
rect 197353 347787 197419 347790
rect 197353 346626 197419 346629
rect 197353 346624 200032 346626
rect 197353 346568 197358 346624
rect 197414 346568 200032 346624
rect 197353 346566 200032 346568
rect 197353 346563 197419 346566
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 197353 345402 197419 345405
rect 197353 345400 200032 345402
rect 197353 345344 197358 345400
rect 197414 345344 200032 345400
rect 197353 345342 200032 345344
rect 197353 345339 197419 345342
rect 197353 344858 197419 344861
rect 197353 344856 200130 344858
rect 197353 344800 197358 344856
rect 197414 344800 200130 344856
rect 197353 344798 200130 344800
rect 197353 344795 197419 344798
rect 200070 344216 200130 344798
rect 111701 343634 111767 343637
rect 111701 343632 161490 343634
rect 111701 343576 111706 343632
rect 111762 343576 161490 343632
rect 111701 343574 161490 343576
rect 111701 343571 111767 343574
rect 161430 342954 161490 343574
rect 197353 343498 197419 343501
rect 197353 343496 200130 343498
rect 197353 343440 197358 343496
rect 197414 343440 200130 343496
rect 197353 343438 200130 343440
rect 197353 343435 197419 343438
rect 200070 342992 200130 343438
rect 560201 343362 560267 343365
rect 556876 343360 560267 343362
rect 556876 343304 560206 343360
rect 560262 343304 560267 343360
rect 556876 343302 560267 343304
rect 560201 343299 560267 343302
rect 172646 342954 172652 342956
rect 161430 342894 172652 342954
rect 172646 342892 172652 342894
rect 172716 342954 172722 342956
rect 192477 342954 192543 342957
rect 172716 342952 192543 342954
rect 172716 342896 192482 342952
rect 192538 342896 192543 342952
rect 172716 342894 192543 342896
rect 172716 342892 172722 342894
rect 192477 342891 192543 342894
rect 197353 341730 197419 341733
rect 197353 341728 200032 341730
rect 197353 341672 197358 341728
rect 197414 341672 200032 341728
rect 197353 341670 200032 341672
rect 197353 341667 197419 341670
rect 46933 340778 46999 340781
rect 48078 340778 48084 340780
rect 46933 340776 48084 340778
rect 46933 340720 46938 340776
rect 46994 340720 48084 340776
rect 46933 340718 48084 340720
rect 46933 340715 46999 340718
rect 48078 340716 48084 340718
rect 48148 340716 48154 340780
rect 197353 340506 197419 340509
rect 197353 340504 200032 340506
rect 197353 340448 197358 340504
rect 197414 340448 200032 340504
rect 197353 340446 200032 340448
rect 197353 340443 197419 340446
rect 46197 340234 46263 340237
rect 46790 340234 46796 340236
rect 46197 340232 46796 340234
rect 46197 340176 46202 340232
rect 46258 340176 46796 340232
rect 46197 340174 46796 340176
rect 46197 340171 46263 340174
rect 46790 340172 46796 340174
rect 46860 340172 46866 340236
rect 3693 340098 3759 340101
rect 174670 340098 174676 340100
rect 3693 340096 174676 340098
rect 3693 340040 3698 340096
rect 3754 340040 174676 340096
rect 3693 340038 174676 340040
rect 3693 340035 3759 340038
rect 174670 340036 174676 340038
rect 174740 340036 174746 340100
rect 35157 339556 35223 339557
rect 35157 339552 35204 339556
rect 35268 339554 35274 339556
rect 35157 339496 35162 339552
rect 35157 339492 35204 339496
rect 35268 339494 35314 339554
rect 35268 339492 35274 339494
rect 35157 339491 35223 339492
rect 197353 339282 197419 339285
rect 197353 339280 200032 339282
rect 197353 339224 197358 339280
rect 197414 339224 200032 339280
rect 197353 339222 200032 339224
rect 197353 339219 197419 339222
rect 583520 338452 584960 338692
rect 197353 337922 197419 337925
rect 197353 337920 200032 337922
rect 197353 337864 197358 337920
rect 197414 337864 200032 337920
rect 197353 337862 200032 337864
rect 197353 337859 197419 337862
rect 197445 336698 197511 336701
rect 197445 336696 200032 336698
rect 197445 336640 197450 336696
rect 197506 336640 200032 336696
rect 197445 336638 200032 336640
rect 197445 336635 197511 336638
rect 197353 336154 197419 336157
rect 197353 336152 200130 336154
rect 197353 336096 197358 336152
rect 197414 336096 200130 336152
rect 197353 336094 200130 336096
rect 197353 336091 197419 336094
rect 200070 335512 200130 336094
rect 560201 335338 560267 335341
rect 556876 335336 560267 335338
rect 556876 335280 560206 335336
rect 560262 335280 560267 335336
rect 556876 335278 560267 335280
rect 560201 335275 560267 335278
rect 197353 334250 197419 334253
rect 197353 334248 200032 334250
rect 197353 334192 197358 334248
rect 197414 334192 200032 334248
rect 197353 334190 200032 334192
rect 197353 334187 197419 334190
rect 28533 333162 28599 333165
rect 29318 333162 30032 333220
rect 28533 333160 30032 333162
rect 28533 333104 28538 333160
rect 28594 333104 29378 333160
rect 28533 333102 29378 333104
rect 28533 333099 28599 333102
rect 197353 333026 197419 333029
rect 197353 333024 200032 333026
rect 197353 332968 197358 333024
rect 197414 332968 200032 333024
rect 197353 332966 200032 332968
rect 197353 332963 197419 332966
rect -960 332196 480 332436
rect 197353 331802 197419 331805
rect 197353 331800 200032 331802
rect 197353 331744 197358 331800
rect 197414 331744 200032 331800
rect 197353 331742 200032 331744
rect 197353 331739 197419 331742
rect 197353 330578 197419 330581
rect 197353 330576 200032 330578
rect 197353 330520 197358 330576
rect 197414 330520 200032 330576
rect 197353 330518 200032 330520
rect 197353 330515 197419 330518
rect 197353 329354 197419 329357
rect 197353 329352 200032 329354
rect 197353 329296 197358 329352
rect 197414 329296 200032 329352
rect 197353 329294 200032 329296
rect 197353 329291 197419 329294
rect 197353 328402 197419 328405
rect 197353 328400 200130 328402
rect 197353 328344 197358 328400
rect 197414 328344 200130 328400
rect 197353 328342 200130 328344
rect 197353 328339 197419 328342
rect 200070 328168 200130 328342
rect 559925 327314 559991 327317
rect 556876 327312 559991 327314
rect 556876 327256 559930 327312
rect 559986 327256 559991 327312
rect 556876 327254 559991 327256
rect 559925 327251 559991 327254
rect 197353 327042 197419 327045
rect 197353 327040 200130 327042
rect 197353 326984 197358 327040
rect 197414 326984 200130 327040
rect 197353 326982 200130 326984
rect 197353 326979 197419 326982
rect 200070 326808 200130 326982
rect 197353 325546 197419 325549
rect 197353 325544 200032 325546
rect 197353 325488 197358 325544
rect 197414 325488 200032 325544
rect 197353 325486 200032 325488
rect 197353 325483 197419 325486
rect 580073 325274 580139 325277
rect 583520 325274 584960 325364
rect 580073 325272 584960 325274
rect 580073 325216 580078 325272
rect 580134 325216 584960 325272
rect 580073 325214 584960 325216
rect 580073 325211 580139 325214
rect 583520 325124 584960 325214
rect 197353 324322 197419 324325
rect 197353 324320 200032 324322
rect 197353 324264 197358 324320
rect 197414 324264 200032 324320
rect 197353 324262 200032 324264
rect 197353 324259 197419 324262
rect 197445 323098 197511 323101
rect 197445 323096 200032 323098
rect 197445 323040 197450 323096
rect 197506 323040 200032 323096
rect 197445 323038 200032 323040
rect 197445 323035 197511 323038
rect 197353 321874 197419 321877
rect 197353 321872 200032 321874
rect 197353 321816 197358 321872
rect 197414 321816 200032 321872
rect 197353 321814 200032 321816
rect 197353 321811 197419 321814
rect 197353 320650 197419 320653
rect 197353 320648 200032 320650
rect 197353 320592 197358 320648
rect 197414 320592 200032 320648
rect 197353 320590 200032 320592
rect 197353 320587 197419 320590
rect 197353 319426 197419 319429
rect 559373 319426 559439 319429
rect 197353 319424 200032 319426
rect -960 319290 480 319380
rect 197353 319368 197358 319424
rect 197414 319368 200032 319424
rect 197353 319366 200032 319368
rect 556876 319424 559439 319426
rect 556876 319368 559378 319424
rect 559434 319368 559439 319424
rect 556876 319366 559439 319368
rect 197353 319363 197419 319366
rect 559373 319363 559439 319366
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 197353 318202 197419 318205
rect 197353 318200 200032 318202
rect 197353 318144 197358 318200
rect 197414 318144 200032 318200
rect 197353 318142 200032 318144
rect 197353 318139 197419 318142
rect 197353 316978 197419 316981
rect 197353 316976 200032 316978
rect 197353 316920 197358 316976
rect 197414 316920 200032 316976
rect 197353 316918 200032 316920
rect 197353 316915 197419 316918
rect 197353 315754 197419 315757
rect 197353 315752 200032 315754
rect 197353 315696 197358 315752
rect 197414 315696 200032 315752
rect 197353 315694 200032 315696
rect 197353 315691 197419 315694
rect 197353 314394 197419 314397
rect 197353 314392 200032 314394
rect 197353 314336 197358 314392
rect 197414 314336 200032 314392
rect 197353 314334 200032 314336
rect 197353 314331 197419 314334
rect 197353 313170 197419 313173
rect 197353 313168 200032 313170
rect 197353 313112 197358 313168
rect 197414 313112 200032 313168
rect 197353 313110 200032 313112
rect 197353 313107 197419 313110
rect 197445 312626 197511 312629
rect 197445 312624 200130 312626
rect 197445 312568 197450 312624
rect 197506 312568 200130 312624
rect 197445 312566 200130 312568
rect 197445 312563 197511 312566
rect 200070 311984 200130 312566
rect 580441 312082 580507 312085
rect 583520 312082 584960 312172
rect 580441 312080 584960 312082
rect 580441 312024 580446 312080
rect 580502 312024 584960 312080
rect 580441 312022 584960 312024
rect 580441 312019 580507 312022
rect 583520 311932 584960 312022
rect 197353 311402 197419 311405
rect 560201 311402 560267 311405
rect 197353 311400 200130 311402
rect 197353 311344 197358 311400
rect 197414 311344 200130 311400
rect 197353 311342 200130 311344
rect 556876 311400 560267 311402
rect 556876 311344 560206 311400
rect 560262 311344 560267 311400
rect 556876 311342 560267 311344
rect 197353 311339 197419 311342
rect 200070 310760 200130 311342
rect 560201 311339 560267 311342
rect 197353 309498 197419 309501
rect 197353 309496 200032 309498
rect 197353 309440 197358 309496
rect 197414 309440 200032 309496
rect 197353 309438 200032 309440
rect 197353 309435 197419 309438
rect 197353 308274 197419 308277
rect 197353 308272 200032 308274
rect 197353 308216 197358 308272
rect 197414 308216 200032 308272
rect 197353 308214 200032 308216
rect 197353 308211 197419 308214
rect 197721 307050 197787 307053
rect 197721 307048 200032 307050
rect 197721 306992 197726 307048
rect 197782 306992 200032 307048
rect 197721 306990 200032 306992
rect 197721 306987 197787 306990
rect -960 306234 480 306324
rect 3969 306234 4035 306237
rect -960 306232 4035 306234
rect -960 306176 3974 306232
rect 4030 306176 4035 306232
rect -960 306174 4035 306176
rect -960 306084 480 306174
rect 3969 306171 4035 306174
rect 197353 305826 197419 305829
rect 197353 305824 200032 305826
rect 197353 305768 197358 305824
rect 197414 305768 200032 305824
rect 197353 305766 200032 305768
rect 197353 305763 197419 305766
rect 197353 304602 197419 304605
rect 197353 304600 200032 304602
rect 197353 304544 197358 304600
rect 197414 304544 200032 304600
rect 197353 304542 200032 304544
rect 197353 304539 197419 304542
rect 197353 303514 197419 303517
rect 197353 303512 200130 303514
rect 197353 303456 197358 303512
rect 197414 303456 200130 303512
rect 197353 303454 200130 303456
rect 197353 303451 197419 303454
rect 200070 303280 200130 303454
rect 559281 303378 559347 303381
rect 556876 303376 559347 303378
rect 556876 303320 559286 303376
rect 559342 303320 559347 303376
rect 556876 303318 559347 303320
rect 559281 303315 559347 303318
rect 197353 302018 197419 302021
rect 197353 302016 200032 302018
rect 197353 301960 197358 302016
rect 197414 301960 200032 302016
rect 197353 301958 200032 301960
rect 197353 301955 197419 301958
rect 197353 300794 197419 300797
rect 197353 300792 200032 300794
rect 197353 300736 197358 300792
rect 197414 300736 200032 300792
rect 197353 300734 200032 300736
rect 197353 300731 197419 300734
rect 197353 299570 197419 299573
rect 197353 299568 200032 299570
rect 197353 299512 197358 299568
rect 197414 299512 200032 299568
rect 197353 299510 200032 299512
rect 197353 299507 197419 299510
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 197353 298346 197419 298349
rect 197353 298344 200032 298346
rect 197353 298288 197358 298344
rect 197414 298288 200032 298344
rect 197353 298286 200032 298288
rect 197353 298283 197419 298286
rect 197353 297122 197419 297125
rect 197353 297120 200032 297122
rect 197353 297064 197358 297120
rect 197414 297064 200032 297120
rect 197353 297062 200032 297064
rect 197353 297059 197419 297062
rect 197353 295490 197419 295493
rect 200070 295490 200130 295864
rect 197353 295488 200130 295490
rect 197353 295432 197358 295488
rect 197414 295432 200130 295488
rect 197353 295430 200130 295432
rect 197353 295427 197419 295430
rect 559005 295354 559071 295357
rect 556876 295352 559071 295354
rect 556876 295296 559010 295352
rect 559066 295296 559071 295352
rect 556876 295294 559071 295296
rect 559005 295291 559071 295294
rect 197353 294402 197419 294405
rect 200070 294402 200130 294640
rect 197353 294400 200130 294402
rect 197353 294344 197358 294400
rect 197414 294344 200130 294400
rect 197353 294342 200130 294344
rect 197353 294339 197419 294342
rect 197353 293450 197419 293453
rect 197353 293448 200032 293450
rect 197353 293392 197358 293448
rect 197414 293392 200032 293448
rect 197353 293390 200032 293392
rect 197353 293387 197419 293390
rect -960 293178 480 293268
rect 3877 293178 3943 293181
rect -960 293176 3943 293178
rect -960 293120 3882 293176
rect 3938 293120 3943 293176
rect -960 293118 3943 293120
rect -960 293028 480 293118
rect 3877 293115 3943 293118
rect 197353 292090 197419 292093
rect 197353 292088 200032 292090
rect 197353 292032 197358 292088
rect 197414 292032 200032 292088
rect 197353 292030 200032 292032
rect 197353 292027 197419 292030
rect 166612 290866 167194 290924
rect 168925 290866 168991 290869
rect 166612 290864 168991 290866
rect 167134 290808 168930 290864
rect 168986 290808 168991 290864
rect 167134 290806 168991 290808
rect 168925 290803 168991 290806
rect 197353 290866 197419 290869
rect 197353 290864 200032 290866
rect 197353 290808 197358 290864
rect 197414 290808 200032 290864
rect 197353 290806 200032 290808
rect 197353 290803 197419 290806
rect 166612 289914 167194 289972
rect 169569 289914 169635 289917
rect 166612 289912 169635 289914
rect 167134 289856 169574 289912
rect 169630 289856 169635 289912
rect 167134 289854 169635 289856
rect 169569 289851 169635 289854
rect 197353 289642 197419 289645
rect 197353 289640 200032 289642
rect 197353 289584 197358 289640
rect 197414 289584 200032 289640
rect 197353 289582 200032 289584
rect 197353 289579 197419 289582
rect 168741 288418 168807 288421
rect 169017 288418 169083 288421
rect 168741 288416 169083 288418
rect 168741 288360 168746 288416
rect 168802 288360 169022 288416
rect 169078 288360 169083 288416
rect 168741 288358 169083 288360
rect 168741 288355 168807 288358
rect 169017 288355 169083 288358
rect 197445 288418 197511 288421
rect 197445 288416 200032 288418
rect 197445 288360 197450 288416
rect 197506 288360 200032 288416
rect 197445 288358 200032 288360
rect 197445 288355 197511 288358
rect 166612 287738 167194 287796
rect 169017 287738 169083 287741
rect 166612 287736 169083 287738
rect 167134 287680 169022 287736
rect 169078 287680 169083 287736
rect 167134 287678 169083 287680
rect 169017 287675 169083 287678
rect 560201 287466 560267 287469
rect 556876 287464 560267 287466
rect 556876 287408 560206 287464
rect 560262 287408 560267 287464
rect 556876 287406 560267 287408
rect 560201 287403 560267 287406
rect 197353 287194 197419 287197
rect 197353 287192 200100 287194
rect 197353 287136 197358 287192
rect 197414 287136 200100 287192
rect 197353 287134 200100 287136
rect 197353 287131 197419 287134
rect 166612 286786 167194 286844
rect 169661 286786 169727 286789
rect 166612 286784 169727 286786
rect 167134 286728 169666 286784
rect 169722 286728 169727 286784
rect 167134 286726 169727 286728
rect 169661 286723 169727 286726
rect 197353 285970 197419 285973
rect 197353 285968 200032 285970
rect 197353 285912 197358 285968
rect 197414 285912 200032 285968
rect 197353 285910 200032 285912
rect 197353 285907 197419 285910
rect 168741 285698 168807 285701
rect 169661 285698 169727 285701
rect 168741 285696 169727 285698
rect 168741 285640 168746 285696
rect 168802 285640 169666 285696
rect 169722 285640 169727 285696
rect 168741 285638 169727 285640
rect 168741 285635 168807 285638
rect 169661 285635 169727 285638
rect 583520 285276 584960 285516
rect 166612 285018 167194 285076
rect 168649 285018 168715 285021
rect 166612 285016 168715 285018
rect 167134 284960 168654 285016
rect 168710 284960 168715 285016
rect 167134 284958 168715 284960
rect 168649 284955 168715 284958
rect 197353 284746 197419 284749
rect 197353 284744 200032 284746
rect 197353 284688 197358 284744
rect 197414 284688 200032 284744
rect 197353 284686 200032 284688
rect 197353 284683 197419 284686
rect 166612 283930 167194 283988
rect 168833 283930 168899 283933
rect 166612 283928 168899 283930
rect 167134 283872 168838 283928
rect 168894 283872 168899 283928
rect 167134 283870 168899 283872
rect 168833 283867 168899 283870
rect 197353 283522 197419 283525
rect 197353 283520 200032 283522
rect 197353 283464 197358 283520
rect 197414 283464 200032 283520
rect 197353 283462 200032 283464
rect 197353 283459 197419 283462
rect 197353 282298 197419 282301
rect 197353 282296 200032 282298
rect 197353 282240 197358 282296
rect 197414 282240 200032 282296
rect 197353 282238 200032 282240
rect 197353 282235 197419 282238
rect 166612 282162 167194 282220
rect 169109 282162 169175 282165
rect 166612 282160 169175 282162
rect 167134 282104 169114 282160
rect 169170 282104 169175 282160
rect 167134 282102 169175 282104
rect 169109 282099 169175 282102
rect 197353 281074 197419 281077
rect 197353 281072 200032 281074
rect 197353 281016 197358 281072
rect 197414 281016 200032 281072
rect 197353 281014 200032 281016
rect 197353 281011 197419 281014
rect -960 279972 480 280212
rect 197353 279170 197419 279173
rect 200070 279170 200130 279680
rect 559925 279442 559991 279445
rect 556876 279440 559991 279442
rect 556876 279384 559930 279440
rect 559986 279384 559991 279440
rect 556876 279382 559991 279384
rect 559925 279379 559991 279382
rect 197353 279168 200130 279170
rect 197353 279112 197358 279168
rect 197414 279112 200130 279168
rect 197353 279110 200130 279112
rect 197353 279107 197419 279110
rect 197353 278490 197419 278493
rect 197353 278488 200032 278490
rect 197353 278432 197358 278488
rect 197414 278432 200032 278488
rect 197353 278430 200032 278432
rect 197353 278427 197419 278430
rect 197445 277266 197511 277269
rect 197445 277264 200032 277266
rect 197445 277208 197450 277264
rect 197506 277208 200032 277264
rect 197445 277206 200032 277208
rect 197445 277203 197511 277206
rect 197353 276042 197419 276045
rect 197353 276040 200032 276042
rect 197353 275984 197358 276040
rect 197414 275984 200032 276040
rect 197353 275982 200032 275984
rect 197353 275979 197419 275982
rect 197353 274818 197419 274821
rect 197353 274816 200032 274818
rect 197353 274760 197358 274816
rect 197414 274760 200032 274816
rect 197353 274758 200032 274760
rect 197353 274755 197419 274758
rect 197353 273594 197419 273597
rect 197353 273592 200032 273594
rect 197353 273536 197358 273592
rect 197414 273536 200032 273592
rect 197353 273534 200032 273536
rect 197353 273531 197419 273534
rect 27153 273322 27219 273325
rect 29318 273322 30032 273380
rect 27153 273320 30032 273322
rect 27153 273264 27158 273320
rect 27214 273264 29378 273320
rect 27153 273262 29378 273264
rect 27153 273259 27219 273262
rect 197353 272370 197419 272373
rect 197353 272368 200032 272370
rect 197353 272312 197358 272368
rect 197414 272312 200032 272368
rect 197353 272310 200032 272312
rect 197353 272307 197419 272310
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect 27337 271690 27403 271693
rect 29318 271690 30032 271748
rect 27337 271688 30032 271690
rect 27337 271632 27342 271688
rect 27398 271632 29378 271688
rect 27337 271630 29378 271632
rect 27337 271627 27403 271630
rect 559557 271418 559623 271421
rect 556876 271416 559623 271418
rect 556876 271360 559562 271416
rect 559618 271360 559623 271416
rect 556876 271358 559623 271360
rect 559557 271355 559623 271358
rect 197353 270602 197419 270605
rect 200070 270602 200130 271112
rect 197353 270600 200130 270602
rect 197353 270544 197358 270600
rect 197414 270544 200130 270600
rect 197353 270542 200130 270544
rect 197353 270539 197419 270542
rect 27429 270330 27495 270333
rect 29318 270330 30032 270388
rect 27429 270328 30032 270330
rect 27429 270272 27434 270328
rect 27490 270272 29378 270328
rect 27429 270270 29378 270272
rect 27429 270267 27495 270270
rect 197813 269922 197879 269925
rect 197813 269920 200032 269922
rect 197813 269864 197818 269920
rect 197874 269864 200032 269920
rect 197813 269862 200032 269864
rect 197813 269859 197879 269862
rect 27061 269106 27127 269109
rect 27245 269106 27311 269109
rect 27061 269104 29378 269106
rect 27061 269048 27066 269104
rect 27122 269048 27250 269104
rect 27306 269048 29378 269104
rect 27061 269046 29378 269048
rect 27061 269043 27127 269046
rect 27245 269043 27311 269046
rect 29318 268892 29378 269046
rect 29318 268832 30032 268892
rect 197353 268562 197419 268565
rect 197353 268560 200032 268562
rect 197353 268504 197358 268560
rect 197414 268504 200032 268560
rect 197353 268502 200032 268504
rect 197353 268499 197419 268502
rect 27521 267610 27587 267613
rect 29318 267610 30032 267668
rect 27521 267608 30032 267610
rect 27521 267552 27526 267608
rect 27582 267552 29378 267608
rect 27521 267550 29378 267552
rect 27521 267547 27587 267550
rect 197353 267338 197419 267341
rect 197353 267336 200032 267338
rect -960 267202 480 267292
rect 197353 267280 197358 267336
rect 197414 267280 200032 267336
rect 197353 267278 200032 267280
rect 197353 267275 197419 267278
rect 3785 267202 3851 267205
rect -960 267200 3851 267202
rect -960 267144 3790 267200
rect 3846 267144 3851 267200
rect -960 267142 3851 267144
rect -960 267052 480 267142
rect 3785 267139 3851 267142
rect 197353 266114 197419 266117
rect 197353 266112 200032 266114
rect 197353 266056 197358 266112
rect 197414 266056 200032 266112
rect 197353 266054 200032 266056
rect 197353 266051 197419 266054
rect 197445 264890 197511 264893
rect 197445 264888 200032 264890
rect 197445 264832 197450 264888
rect 197506 264832 200032 264888
rect 197445 264830 200032 264832
rect 197445 264827 197511 264830
rect 169201 264074 169267 264077
rect 167134 264072 169267 264074
rect 167134 264016 169206 264072
rect 169262 264016 169267 264072
rect 167134 264014 169267 264016
rect 167134 263996 167194 264014
rect 169201 264011 169267 264014
rect 166612 263936 167194 263996
rect 197353 263666 197419 263669
rect 197353 263664 200100 263666
rect 197353 263608 197358 263664
rect 197414 263608 200100 263664
rect 197353 263606 200100 263608
rect 197353 263603 197419 263606
rect 560201 263530 560267 263533
rect 556876 263528 560267 263530
rect 556876 263472 560206 263528
rect 560262 263472 560267 263528
rect 556876 263470 560267 263472
rect 560201 263467 560267 263470
rect 197353 262442 197419 262445
rect 197353 262440 200032 262442
rect 197353 262384 197358 262440
rect 197414 262384 200032 262440
rect 197353 262382 200032 262384
rect 197353 262379 197419 262382
rect 166612 262306 167194 262364
rect 168373 262306 168439 262309
rect 166612 262304 168439 262306
rect 167134 262248 168378 262304
rect 168434 262248 168439 262304
rect 167134 262246 168439 262248
rect 168373 262243 168439 262246
rect 166612 262034 167194 262092
rect 168557 262034 168623 262037
rect 166612 262032 168623 262034
rect 167134 261976 168562 262032
rect 168618 261976 168623 262032
rect 167134 261974 168623 261976
rect 168557 261971 168623 261974
rect 197353 261218 197419 261221
rect 197353 261216 200032 261218
rect 197353 261160 197358 261216
rect 197414 261160 200032 261216
rect 197353 261158 200032 261160
rect 197353 261155 197419 261158
rect 168046 259524 168052 259588
rect 168116 259586 168122 259588
rect 199377 259586 199443 259589
rect 200002 259586 200062 259964
rect 168116 259584 200062 259586
rect 168116 259528 199382 259584
rect 199438 259528 200062 259584
rect 168116 259526 200062 259528
rect 168116 259524 168122 259526
rect 199377 259523 199443 259526
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 197353 258770 197419 258773
rect 199469 258770 199535 258773
rect 197353 258768 200032 258770
rect 197353 258712 197358 258768
rect 197414 258712 199474 258768
rect 199530 258712 200032 258768
rect 583520 258756 584960 258846
rect 197353 258710 200032 258712
rect 197353 258707 197419 258710
rect 199469 258707 199535 258710
rect 197905 257410 197971 257413
rect 197905 257408 200032 257410
rect 197905 257352 197910 257408
rect 197966 257352 200032 257408
rect 197905 257350 200032 257352
rect 197905 257347 197971 257350
rect 197997 256186 198063 256189
rect 197997 256184 200100 256186
rect 197997 256128 198002 256184
rect 198058 256128 200100 256184
rect 197997 256126 200100 256128
rect 197997 256123 198063 256126
rect 560017 255506 560083 255509
rect 556876 255504 560083 255506
rect 556876 255448 560022 255504
rect 560078 255448 560083 255504
rect 556876 255446 560083 255448
rect 560017 255443 560083 255446
rect 197537 254826 197603 254829
rect 198089 254826 198155 254829
rect 200070 254826 200130 254928
rect 197537 254824 200130 254826
rect 197537 254768 197542 254824
rect 197598 254768 198094 254824
rect 198150 254768 200130 254824
rect 197537 254766 200130 254768
rect 197537 254763 197603 254766
rect 198089 254763 198155 254766
rect -960 254146 480 254236
rect 3693 254146 3759 254149
rect -960 254144 3759 254146
rect -960 254088 3698 254144
rect 3754 254088 3759 254144
rect -960 254086 3759 254088
rect -960 253996 480 254086
rect 3693 254083 3759 254086
rect 27337 253874 27403 253877
rect 198181 253874 198247 253877
rect 27337 253872 199578 253874
rect 27337 253816 27342 253872
rect 27398 253816 198186 253872
rect 198242 253816 199578 253872
rect 27337 253814 199578 253816
rect 27337 253811 27403 253814
rect 198181 253811 198247 253814
rect 60641 253740 60707 253741
rect 65701 253740 65767 253741
rect 70669 253740 70735 253741
rect 75545 253740 75611 253741
rect 98269 253740 98335 253741
rect 115657 253740 115723 253741
rect 118325 253740 118391 253741
rect 60600 253738 60606 253740
rect 60550 253678 60606 253738
rect 60670 253736 60707 253740
rect 65632 253738 65638 253740
rect 60702 253680 60707 253736
rect 60600 253676 60606 253678
rect 60670 253676 60707 253680
rect 65610 253678 65638 253738
rect 65632 253676 65638 253678
rect 65702 253736 65767 253740
rect 70664 253738 70670 253740
rect 65702 253680 65706 253736
rect 65762 253680 65767 253736
rect 65702 253676 65767 253680
rect 70578 253678 70670 253738
rect 70664 253676 70670 253678
rect 70734 253676 70740 253740
rect 75545 253736 75566 253740
rect 75630 253738 75636 253740
rect 75545 253680 75550 253736
rect 75545 253676 75566 253680
rect 75630 253678 75702 253738
rect 98269 253736 98278 253740
rect 98342 253738 98348 253740
rect 115606 253738 115612 253740
rect 98269 253680 98274 253736
rect 75630 253676 75636 253678
rect 98269 253676 98278 253680
rect 98342 253678 98426 253738
rect 115566 253678 115612 253738
rect 115676 253736 115723 253740
rect 118264 253738 118270 253740
rect 115718 253680 115723 253736
rect 98342 253676 98348 253678
rect 115606 253676 115612 253678
rect 115676 253676 115723 253680
rect 118234 253678 118270 253738
rect 118334 253736 118391 253740
rect 118386 253680 118391 253736
rect 118264 253676 118270 253678
rect 118334 253676 118391 253680
rect 60641 253675 60707 253676
rect 65701 253675 65767 253676
rect 70669 253675 70735 253676
rect 75545 253675 75611 253676
rect 98269 253675 98335 253676
rect 115657 253675 115723 253676
rect 118325 253675 118391 253676
rect 123017 253740 123083 253741
rect 125501 253740 125567 253741
rect 128077 253740 128143 253741
rect 123017 253736 123030 253740
rect 123094 253738 123100 253740
rect 125472 253738 125478 253740
rect 123017 253680 123022 253736
rect 123017 253676 123030 253680
rect 123094 253678 123174 253738
rect 125410 253678 125478 253738
rect 125542 253736 125567 253740
rect 128056 253738 128062 253740
rect 125562 253680 125567 253736
rect 123094 253676 123100 253678
rect 125472 253676 125478 253678
rect 125542 253676 125567 253680
rect 127986 253678 128062 253738
rect 128126 253736 128143 253740
rect 128138 253680 128143 253736
rect 199518 253740 199578 253814
rect 199518 253680 200062 253740
rect 128056 253676 128062 253678
rect 128126 253676 128143 253680
rect 123017 253675 123083 253676
rect 125501 253675 125567 253676
rect 128077 253675 128143 253676
rect 43345 253604 43411 253605
rect 130561 253604 130627 253605
rect 43328 253602 43334 253604
rect 43254 253542 43334 253602
rect 43398 253600 43411 253604
rect 130510 253602 130516 253604
rect 43406 253544 43411 253600
rect 43328 253540 43334 253542
rect 43398 253540 43411 253544
rect 130470 253542 130516 253602
rect 130580 253600 130627 253604
rect 130622 253544 130627 253600
rect 130510 253540 130516 253542
rect 130580 253540 130627 253544
rect 43345 253539 43411 253540
rect 130561 253539 130627 253540
rect 136449 253604 136515 253605
rect 136449 253600 136494 253604
rect 136558 253602 136564 253604
rect 136449 253544 136454 253600
rect 136449 253540 136494 253544
rect 136558 253542 136606 253602
rect 136558 253540 136564 253542
rect 136449 253539 136515 253540
rect 132953 253468 133019 253469
rect 132902 253466 132908 253468
rect 132862 253406 132908 253466
rect 132972 253464 133019 253468
rect 133014 253408 133019 253464
rect 132902 253404 132908 253406
rect 132972 253404 133019 253408
rect 132953 253403 133019 253404
rect 27153 252650 27219 252653
rect 166993 252650 167059 252653
rect 27153 252648 167059 252650
rect 27153 252592 27158 252648
rect 27214 252592 166998 252648
rect 167054 252592 167059 252648
rect 27153 252590 167059 252592
rect 27153 252587 27219 252590
rect 166993 252587 167059 252590
rect 26969 252514 27035 252517
rect 27429 252514 27495 252517
rect 26969 252512 27495 252514
rect 26969 252456 26974 252512
rect 27030 252456 27434 252512
rect 27490 252456 27495 252512
rect 26969 252454 27495 252456
rect 26969 252451 27035 252454
rect 27429 252451 27495 252454
rect 63166 252452 63172 252516
rect 63236 252514 63242 252516
rect 63401 252514 63467 252517
rect 68185 252516 68251 252517
rect 73153 252516 73219 252517
rect 78121 252516 78187 252517
rect 68134 252514 68140 252516
rect 63236 252512 63467 252514
rect 63236 252456 63406 252512
rect 63462 252456 63467 252512
rect 63236 252454 63467 252456
rect 68094 252454 68140 252514
rect 68204 252512 68251 252516
rect 73102 252514 73108 252516
rect 68246 252456 68251 252512
rect 63236 252452 63242 252454
rect 63401 252451 63467 252454
rect 68134 252452 68140 252454
rect 68204 252452 68251 252456
rect 73062 252454 73108 252514
rect 73172 252512 73219 252516
rect 78070 252514 78076 252516
rect 73214 252456 73219 252512
rect 73102 252452 73108 252454
rect 73172 252452 73219 252456
rect 78030 252454 78076 252514
rect 78140 252512 78187 252516
rect 78182 252456 78187 252512
rect 78070 252452 78076 252454
rect 78140 252452 78187 252456
rect 80646 252452 80652 252516
rect 80716 252514 80722 252516
rect 81249 252514 81315 252517
rect 80716 252512 81315 252514
rect 80716 252456 81254 252512
rect 81310 252456 81315 252512
rect 80716 252454 81315 252456
rect 80716 252452 80722 252454
rect 68185 252451 68251 252452
rect 73153 252451 73219 252452
rect 78121 252451 78187 252452
rect 81249 252451 81315 252454
rect 83038 252452 83044 252516
rect 83108 252514 83114 252516
rect 83549 252514 83615 252517
rect 85665 252516 85731 252517
rect 88241 252516 88307 252517
rect 90817 252516 90883 252517
rect 93209 252516 93275 252517
rect 95601 252516 95667 252517
rect 100569 252516 100635 252517
rect 103145 252516 103211 252517
rect 85614 252514 85620 252516
rect 83108 252512 83615 252514
rect 83108 252456 83554 252512
rect 83610 252456 83615 252512
rect 83108 252454 83615 252456
rect 85574 252454 85620 252514
rect 85684 252512 85731 252516
rect 88190 252514 88196 252516
rect 85726 252456 85731 252512
rect 83108 252452 83114 252454
rect 83549 252451 83615 252454
rect 85614 252452 85620 252454
rect 85684 252452 85731 252456
rect 88150 252454 88196 252514
rect 88260 252512 88307 252516
rect 90766 252514 90772 252516
rect 88302 252456 88307 252512
rect 88190 252452 88196 252454
rect 88260 252452 88307 252456
rect 90726 252454 90772 252514
rect 90836 252512 90883 252516
rect 93158 252514 93164 252516
rect 90878 252456 90883 252512
rect 90766 252452 90772 252454
rect 90836 252452 90883 252456
rect 93118 252454 93164 252514
rect 93228 252512 93275 252516
rect 95550 252514 95556 252516
rect 93270 252456 93275 252512
rect 93158 252452 93164 252454
rect 93228 252452 93275 252456
rect 95510 252454 95556 252514
rect 95620 252512 95667 252516
rect 100518 252514 100524 252516
rect 95662 252456 95667 252512
rect 95550 252452 95556 252454
rect 95620 252452 95667 252456
rect 100478 252454 100524 252514
rect 100588 252512 100635 252516
rect 103094 252514 103100 252516
rect 100630 252456 100635 252512
rect 100518 252452 100524 252454
rect 100588 252452 100635 252456
rect 103054 252454 103100 252514
rect 103164 252512 103211 252516
rect 103206 252456 103211 252512
rect 103094 252452 103100 252454
rect 103164 252452 103211 252456
rect 105670 252452 105676 252516
rect 105740 252514 105746 252516
rect 106089 252514 106155 252517
rect 105740 252512 106155 252514
rect 105740 252456 106094 252512
rect 106150 252456 106155 252512
rect 105740 252454 106155 252456
rect 105740 252452 105746 252454
rect 85665 252451 85731 252452
rect 88241 252451 88307 252452
rect 90817 252451 90883 252452
rect 93209 252451 93275 252452
rect 95601 252451 95667 252452
rect 100569 252451 100635 252452
rect 103145 252451 103211 252452
rect 106089 252451 106155 252454
rect 108062 252452 108068 252516
rect 108132 252514 108138 252516
rect 108481 252514 108547 252517
rect 110505 252516 110571 252517
rect 113081 252516 113147 252517
rect 110454 252514 110460 252516
rect 108132 252512 108547 252514
rect 108132 252456 108486 252512
rect 108542 252456 108547 252512
rect 108132 252454 108547 252456
rect 110414 252454 110460 252514
rect 110524 252512 110571 252516
rect 113030 252514 113036 252516
rect 110566 252456 110571 252512
rect 108132 252452 108138 252454
rect 108481 252451 108547 252454
rect 110454 252452 110460 252454
rect 110524 252452 110571 252456
rect 112990 252454 113036 252514
rect 113100 252512 113147 252516
rect 113142 252456 113147 252512
rect 113030 252452 113036 252454
rect 113100 252452 113147 252456
rect 115422 252452 115428 252516
rect 115492 252514 115498 252516
rect 115841 252514 115907 252517
rect 115492 252512 115907 252514
rect 115492 252456 115846 252512
rect 115902 252456 115907 252512
rect 115492 252454 115907 252456
rect 115492 252452 115498 252454
rect 110505 252451 110571 252452
rect 113081 252451 113147 252452
rect 115841 252451 115907 252454
rect 120574 252452 120580 252516
rect 120644 252514 120650 252516
rect 120901 252514 120967 252517
rect 120644 252512 120967 252514
rect 120644 252456 120906 252512
rect 120962 252456 120967 252512
rect 120644 252454 120967 252456
rect 120644 252452 120650 252454
rect 120901 252451 120967 252454
rect 135846 252452 135852 252516
rect 135916 252514 135922 252516
rect 135989 252514 136055 252517
rect 135916 252512 136055 252514
rect 135916 252456 135994 252512
rect 136050 252456 136055 252512
rect 135916 252454 136055 252456
rect 135916 252452 135922 252454
rect 135989 252451 136055 252454
rect 143349 252516 143415 252517
rect 148317 252516 148383 252517
rect 143349 252512 143396 252516
rect 143460 252514 143466 252516
rect 143349 252456 143354 252512
rect 143349 252452 143396 252456
rect 143460 252454 143506 252514
rect 143460 252452 143466 252454
rect 144862 252452 144868 252516
rect 144932 252514 144938 252516
rect 145966 252514 145972 252516
rect 144932 252454 145972 252514
rect 144932 252452 144938 252454
rect 145966 252452 145972 252454
rect 146036 252514 146042 252516
rect 147070 252514 147076 252516
rect 146036 252454 147076 252514
rect 146036 252452 146042 252454
rect 147070 252452 147076 252454
rect 147140 252514 147146 252516
rect 148317 252514 148364 252516
rect 147140 252512 148364 252514
rect 148428 252514 148434 252516
rect 147140 252456 148322 252512
rect 147140 252454 148364 252456
rect 147140 252452 147146 252454
rect 148317 252452 148364 252454
rect 148428 252454 148474 252514
rect 148428 252452 148434 252454
rect 150566 252452 150572 252516
rect 150636 252514 150642 252516
rect 151077 252514 151143 252517
rect 150636 252512 151143 252514
rect 150636 252456 151082 252512
rect 151138 252456 151143 252512
rect 150636 252454 151143 252456
rect 150636 252452 150642 252454
rect 143349 252451 143415 252452
rect 148317 252451 148383 252452
rect 151077 252451 151143 252454
rect 197445 252514 197511 252517
rect 198273 252514 198339 252517
rect 197445 252512 200032 252514
rect 197445 252456 197450 252512
rect 197506 252456 198278 252512
rect 198334 252456 200032 252512
rect 197445 252454 200032 252456
rect 197445 252451 197511 252454
rect 198273 252451 198339 252454
rect 28625 252378 28691 252381
rect 43110 252378 43116 252380
rect 28625 252376 43116 252378
rect 28625 252320 28630 252376
rect 28686 252320 43116 252376
rect 28625 252318 43116 252320
rect 28625 252315 28691 252318
rect 43110 252316 43116 252318
rect 43180 252378 43186 252380
rect 43180 252318 45570 252378
rect 43180 252316 43186 252318
rect 45510 252242 45570 252318
rect 109534 252316 109540 252380
rect 109604 252378 109610 252380
rect 110321 252378 110387 252381
rect 109604 252376 110387 252378
rect 109604 252320 110326 252376
rect 110382 252320 110387 252376
rect 109604 252318 110387 252320
rect 109604 252316 109610 252318
rect 110321 252315 110387 252318
rect 110822 252316 110828 252380
rect 110892 252378 110898 252380
rect 111701 252378 111767 252381
rect 110892 252376 111767 252378
rect 110892 252320 111706 252376
rect 111762 252320 111767 252376
rect 110892 252318 111767 252320
rect 110892 252316 110898 252318
rect 111701 252315 111767 252318
rect 112110 252316 112116 252380
rect 112180 252378 112186 252380
rect 112989 252378 113055 252381
rect 112180 252376 113055 252378
rect 112180 252320 112994 252376
rect 113050 252320 113055 252376
rect 112180 252318 113055 252320
rect 112180 252316 112186 252318
rect 112989 252315 113055 252318
rect 113214 252316 113220 252380
rect 113284 252378 113290 252380
rect 114461 252378 114527 252381
rect 113284 252376 114527 252378
rect 113284 252320 114466 252376
rect 114522 252320 114527 252376
rect 113284 252318 114527 252320
rect 113284 252316 113290 252318
rect 114461 252315 114527 252318
rect 125910 252316 125916 252380
rect 125980 252378 125986 252380
rect 126881 252378 126947 252381
rect 125980 252376 126947 252378
rect 125980 252320 126886 252376
rect 126942 252320 126947 252376
rect 125980 252318 126947 252320
rect 125980 252316 125986 252318
rect 126881 252315 126947 252318
rect 129549 252380 129615 252381
rect 132033 252380 132099 252381
rect 129549 252376 129596 252380
rect 129660 252378 129666 252380
rect 131982 252378 131988 252380
rect 129549 252320 129554 252376
rect 129549 252316 129596 252320
rect 129660 252318 129706 252378
rect 131942 252318 131988 252378
rect 132052 252376 132099 252380
rect 132094 252320 132099 252376
rect 129660 252316 129666 252318
rect 131982 252316 131988 252318
rect 132052 252316 132099 252320
rect 133086 252316 133092 252380
rect 133156 252378 133162 252380
rect 133781 252378 133847 252381
rect 138289 252380 138355 252381
rect 138238 252378 138244 252380
rect 133156 252376 133847 252378
rect 133156 252320 133786 252376
rect 133842 252320 133847 252376
rect 133156 252318 133847 252320
rect 138198 252318 138244 252378
rect 138308 252376 138355 252380
rect 138350 252320 138355 252376
rect 133156 252316 133162 252318
rect 129549 252315 129615 252316
rect 132033 252315 132099 252316
rect 133781 252315 133847 252318
rect 138238 252316 138244 252318
rect 138308 252316 138355 252320
rect 142286 252316 142292 252380
rect 142356 252378 142362 252380
rect 143441 252378 143507 252381
rect 142356 252376 143507 252378
rect 142356 252320 143446 252376
rect 143502 252320 143507 252376
rect 142356 252318 143507 252320
rect 142356 252316 142362 252318
rect 138289 252315 138355 252316
rect 143441 252315 143507 252318
rect 168046 252242 168052 252244
rect 45510 252182 168052 252242
rect 168046 252180 168052 252182
rect 168116 252180 168122 252244
rect 150014 252044 150020 252108
rect 150084 252106 150090 252108
rect 167085 252106 167151 252109
rect 150084 252104 167151 252106
rect 150084 252048 167090 252104
rect 167146 252048 167151 252104
rect 150084 252046 167151 252048
rect 150084 252044 150090 252046
rect 167085 252043 167151 252046
rect 114369 251972 114435 251973
rect 114318 251970 114324 251972
rect 114278 251910 114324 251970
rect 114388 251968 114435 251972
rect 114430 251912 114435 251968
rect 114318 251908 114324 251910
rect 114388 251908 114435 251912
rect 141182 251908 141188 251972
rect 141252 251970 141258 251972
rect 142061 251970 142127 251973
rect 141252 251968 142127 251970
rect 141252 251912 142066 251968
rect 142122 251912 142127 251968
rect 141252 251910 142127 251912
rect 141252 251908 141258 251910
rect 114369 251907 114435 251908
rect 142061 251907 142127 251910
rect 120206 251636 120212 251700
rect 120276 251698 120282 251700
rect 121177 251698 121243 251701
rect 120276 251696 121243 251698
rect 120276 251640 121182 251696
rect 121238 251640 121243 251696
rect 120276 251638 121243 251640
rect 120276 251636 120282 251638
rect 121177 251635 121243 251638
rect 135294 251636 135300 251700
rect 135364 251698 135370 251700
rect 136357 251698 136423 251701
rect 135364 251696 136423 251698
rect 135364 251640 136362 251696
rect 136418 251640 136423 251696
rect 135364 251638 136423 251640
rect 135364 251636 135370 251638
rect 136357 251635 136423 251638
rect 26969 251562 27035 251565
rect 197537 251562 197603 251565
rect 26969 251560 197603 251562
rect 26969 251504 26974 251560
rect 27030 251504 197542 251560
rect 197598 251504 197603 251560
rect 26969 251502 197603 251504
rect 26969 251499 27035 251502
rect 197537 251499 197603 251502
rect 43345 251426 43411 251429
rect 169845 251426 169911 251429
rect 43345 251424 169911 251426
rect 43345 251368 43350 251424
rect 43406 251368 169850 251424
rect 169906 251368 169911 251424
rect 43345 251366 169911 251368
rect 43345 251363 43411 251366
rect 169845 251363 169911 251366
rect 107326 251228 107332 251292
rect 107396 251290 107402 251292
rect 107561 251290 107627 251293
rect 107396 251288 107627 251290
rect 107396 251232 107566 251288
rect 107622 251232 107627 251288
rect 107396 251230 107627 251232
rect 107396 251228 107402 251230
rect 107561 251227 107627 251230
rect 108430 251228 108436 251292
rect 108500 251290 108506 251292
rect 108941 251290 109007 251293
rect 108500 251288 109007 251290
rect 108500 251232 108946 251288
rect 109002 251232 109007 251288
rect 108500 251230 109007 251232
rect 108500 251228 108506 251230
rect 108941 251227 109007 251230
rect 116710 251228 116716 251292
rect 116780 251290 116786 251292
rect 117221 251290 117287 251293
rect 116780 251288 117287 251290
rect 116780 251232 117226 251288
rect 117282 251232 117287 251288
rect 116780 251230 117287 251232
rect 116780 251228 116786 251230
rect 117221 251227 117287 251230
rect 117814 251228 117820 251292
rect 117884 251290 117890 251292
rect 118601 251290 118667 251293
rect 117884 251288 118667 251290
rect 117884 251232 118606 251288
rect 118662 251232 118667 251288
rect 117884 251230 118667 251232
rect 117884 251228 117890 251230
rect 118601 251227 118667 251230
rect 118918 251228 118924 251292
rect 118988 251290 118994 251292
rect 119981 251290 120047 251293
rect 118988 251288 120047 251290
rect 118988 251232 119986 251288
rect 120042 251232 120047 251288
rect 118988 251230 120047 251232
rect 118988 251228 118994 251230
rect 119981 251227 120047 251230
rect 121269 251292 121335 251293
rect 121269 251288 121316 251292
rect 121380 251290 121386 251292
rect 121269 251232 121274 251288
rect 121269 251228 121316 251232
rect 121380 251230 121426 251290
rect 121380 251228 121386 251230
rect 122598 251228 122604 251292
rect 122668 251290 122674 251292
rect 122741 251290 122807 251293
rect 122668 251288 122807 251290
rect 122668 251232 122746 251288
rect 122802 251232 122807 251288
rect 122668 251230 122807 251232
rect 122668 251228 122674 251230
rect 121269 251227 121335 251228
rect 122741 251227 122807 251230
rect 123702 251228 123708 251292
rect 123772 251290 123778 251292
rect 124121 251290 124187 251293
rect 123772 251288 124187 251290
rect 123772 251232 124126 251288
rect 124182 251232 124187 251288
rect 123772 251230 124187 251232
rect 123772 251228 123778 251230
rect 124121 251227 124187 251230
rect 124806 251228 124812 251292
rect 124876 251290 124882 251292
rect 125501 251290 125567 251293
rect 124876 251288 125567 251290
rect 124876 251232 125506 251288
rect 125562 251232 125567 251288
rect 124876 251230 125567 251232
rect 124876 251228 124882 251230
rect 125501 251227 125567 251230
rect 127198 251228 127204 251292
rect 127268 251290 127274 251292
rect 128261 251290 128327 251293
rect 127268 251288 128327 251290
rect 127268 251232 128266 251288
rect 128322 251232 128327 251288
rect 127268 251230 128327 251232
rect 127268 251228 127274 251230
rect 128261 251227 128327 251230
rect 128486 251228 128492 251292
rect 128556 251290 128562 251292
rect 129641 251290 129707 251293
rect 128556 251288 129707 251290
rect 128556 251232 129646 251288
rect 129702 251232 129707 251288
rect 128556 251230 129707 251232
rect 128556 251228 128562 251230
rect 129641 251227 129707 251230
rect 130694 251228 130700 251292
rect 130764 251290 130770 251292
rect 131021 251290 131087 251293
rect 130764 251288 131087 251290
rect 130764 251232 131026 251288
rect 131082 251232 131087 251288
rect 130764 251230 131087 251232
rect 130764 251228 130770 251230
rect 131021 251227 131087 251230
rect 134190 251228 134196 251292
rect 134260 251290 134266 251292
rect 135161 251290 135227 251293
rect 137921 251292 137987 251293
rect 137870 251290 137876 251292
rect 134260 251288 135227 251290
rect 134260 251232 135166 251288
rect 135222 251232 135227 251288
rect 134260 251230 135227 251232
rect 137830 251230 137876 251290
rect 137940 251288 137987 251292
rect 137982 251232 137987 251288
rect 134260 251228 134266 251230
rect 135161 251227 135227 251230
rect 137870 251228 137876 251230
rect 137940 251228 137987 251232
rect 138974 251228 138980 251292
rect 139044 251290 139050 251292
rect 139209 251290 139275 251293
rect 139044 251288 139275 251290
rect 139044 251232 139214 251288
rect 139270 251232 139275 251288
rect 139044 251230 139275 251232
rect 139044 251228 139050 251230
rect 137921 251227 137987 251228
rect 139209 251227 139275 251230
rect 140078 251228 140084 251292
rect 140148 251290 140154 251292
rect 140681 251290 140747 251293
rect 140148 251288 140747 251290
rect 140148 251232 140686 251288
rect 140742 251232 140747 251288
rect 140148 251230 140747 251232
rect 140148 251228 140154 251230
rect 140681 251227 140747 251230
rect 197353 251290 197419 251293
rect 197353 251288 200032 251290
rect 197353 251232 197358 251288
rect 197414 251232 200032 251288
rect 197353 251230 200032 251232
rect 197353 251227 197419 251230
rect 50337 250474 50403 250477
rect 198590 250474 198596 250476
rect 50337 250472 198596 250474
rect 50337 250416 50342 250472
rect 50398 250416 198596 250472
rect 50337 250414 198596 250416
rect 50337 250411 50403 250414
rect 198590 250412 198596 250414
rect 198660 250474 198666 250476
rect 198660 250414 200062 250474
rect 198660 250412 198666 250414
rect 200002 250036 200062 250414
rect 197261 248842 197327 248845
rect 197261 248840 200032 248842
rect 197261 248784 197266 248840
rect 197322 248784 200032 248840
rect 197261 248782 200032 248784
rect 197261 248779 197327 248782
rect 198774 247964 198780 248028
rect 198844 248026 198850 248028
rect 198844 247966 200130 248026
rect 198844 247964 198850 247966
rect 200070 247656 200130 247966
rect 560201 247482 560267 247485
rect 556876 247480 560267 247482
rect 556876 247424 560206 247480
rect 560262 247424 560267 247480
rect 556876 247422 560267 247424
rect 560201 247419 560267 247422
rect 197353 246394 197419 246397
rect 197353 246392 200032 246394
rect 197353 246336 197358 246392
rect 197414 246336 200032 246392
rect 197353 246334 200032 246336
rect 197353 246331 197419 246334
rect 167494 245652 167500 245716
rect 167564 245714 167570 245716
rect 167637 245714 167703 245717
rect 167564 245712 167703 245714
rect 167564 245656 167642 245712
rect 167698 245656 167703 245712
rect 167564 245654 167703 245656
rect 167564 245652 167570 245654
rect 167637 245651 167703 245654
rect 580257 245578 580323 245581
rect 583520 245578 584960 245668
rect 580257 245576 584960 245578
rect 580257 245520 580262 245576
rect 580318 245520 584960 245576
rect 580257 245518 584960 245520
rect 580257 245515 580323 245518
rect 583520 245428 584960 245518
rect 197353 245034 197419 245037
rect 197353 245032 200032 245034
rect 197353 244976 197358 245032
rect 197414 244976 200032 245032
rect 197353 244974 200032 244976
rect 197353 244971 197419 244974
rect 197353 243810 197419 243813
rect 197353 243808 200032 243810
rect 197353 243752 197358 243808
rect 197414 243752 200032 243808
rect 197353 243750 200032 243752
rect 197353 243747 197419 243750
rect 197353 242586 197419 242589
rect 197353 242584 200032 242586
rect 197353 242528 197358 242584
rect 197414 242528 200032 242584
rect 197353 242526 200032 242528
rect 197353 242523 197419 242526
rect 197537 241362 197603 241365
rect 197537 241360 200032 241362
rect 197537 241304 197542 241360
rect 197598 241304 200032 241360
rect 197537 241302 200032 241304
rect 197537 241299 197603 241302
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 197445 239594 197511 239597
rect 200070 239594 200130 240104
rect 560201 239594 560267 239597
rect 197445 239592 200130 239594
rect 197445 239536 197450 239592
rect 197506 239536 200130 239592
rect 197445 239534 200130 239536
rect 556876 239592 560267 239594
rect 556876 239536 560206 239592
rect 560262 239536 560267 239592
rect 556876 239534 560267 239536
rect 197445 239531 197511 239534
rect 560201 239531 560267 239534
rect 197353 238914 197419 238917
rect 197353 238912 200100 238914
rect 197353 238856 197358 238912
rect 197414 238856 200100 238912
rect 197353 238854 200100 238856
rect 197353 238851 197419 238854
rect 168189 238644 168255 238645
rect 168189 238640 168236 238644
rect 168300 238642 168306 238644
rect 168189 238584 168194 238640
rect 168189 238580 168236 238584
rect 168300 238582 168346 238642
rect 168300 238580 168306 238582
rect 168189 238579 168255 238580
rect 199285 237690 199351 237693
rect 199285 237688 200032 237690
rect 199285 237632 199290 237688
rect 199346 237632 200032 237688
rect 199285 237630 200032 237632
rect 199285 237627 199351 237630
rect 197353 236466 197419 236469
rect 197353 236464 200032 236466
rect 197353 236408 197358 236464
rect 197414 236408 200032 236464
rect 197353 236406 200032 236408
rect 197353 236403 197419 236406
rect 197721 235242 197787 235245
rect 197721 235240 200032 235242
rect 197721 235184 197726 235240
rect 197782 235184 200032 235240
rect 197721 235182 200032 235184
rect 197721 235179 197787 235182
rect 197353 233882 197419 233885
rect 197353 233880 200032 233882
rect 197353 233824 197358 233880
rect 197414 233824 200032 233880
rect 197353 233822 200032 233824
rect 197353 233819 197419 233822
rect 197353 232658 197419 232661
rect 197813 232658 197879 232661
rect 197353 232656 200032 232658
rect 197353 232600 197358 232656
rect 197414 232600 197818 232656
rect 197874 232600 200032 232656
rect 197353 232598 200032 232600
rect 197353 232595 197419 232598
rect 197813 232595 197879 232598
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect 197353 231706 197419 231709
rect 197353 231704 200130 231706
rect 197353 231648 197358 231704
rect 197414 231648 200130 231704
rect 197353 231646 200130 231648
rect 197353 231643 197419 231646
rect 200070 231472 200130 231646
rect 559189 231570 559255 231573
rect 556876 231568 559255 231570
rect 556876 231512 559194 231568
rect 559250 231512 559255 231568
rect 556876 231510 559255 231512
rect 559189 231507 559255 231510
rect 197537 230210 197603 230213
rect 199193 230210 199259 230213
rect 197537 230208 200032 230210
rect 197537 230152 197542 230208
rect 197598 230152 199198 230208
rect 199254 230152 200032 230208
rect 197537 230150 200032 230152
rect 197537 230147 197603 230150
rect 199193 230147 199259 230150
rect 168557 228986 168623 228989
rect 168966 228986 168972 228988
rect 168557 228984 168972 228986
rect 168557 228928 168562 228984
rect 168618 228928 168972 228984
rect 168557 228926 168972 228928
rect 168557 228923 168623 228926
rect 168966 228924 168972 228926
rect 169036 228924 169042 228988
rect 198365 228986 198431 228989
rect 198365 228984 200032 228986
rect 198365 228928 198370 228984
rect 198426 228928 200032 228984
rect 198365 228926 200032 228928
rect 198365 228923 198431 228926
rect -960 227884 480 228124
rect 35157 227764 35223 227765
rect 46749 227764 46815 227765
rect 35157 227760 35204 227764
rect 35268 227762 35274 227764
rect 35157 227704 35162 227760
rect 35157 227700 35204 227704
rect 35268 227702 35314 227762
rect 46749 227760 46796 227764
rect 46860 227762 46866 227764
rect 47577 227762 47643 227765
rect 48078 227762 48084 227764
rect 46749 227704 46754 227760
rect 35268 227700 35274 227702
rect 46749 227700 46796 227704
rect 46860 227702 46906 227762
rect 47577 227760 48084 227762
rect 47577 227704 47582 227760
rect 47638 227704 48084 227760
rect 47577 227702 48084 227704
rect 46860 227700 46866 227702
rect 35157 227699 35223 227700
rect 46749 227699 46815 227700
rect 47577 227699 47643 227702
rect 48078 227700 48084 227702
rect 48148 227700 48154 227764
rect 199101 227762 199167 227765
rect 199101 227760 200032 227762
rect 199101 227704 199106 227760
rect 199162 227704 200032 227760
rect 199101 227702 200032 227704
rect 199101 227699 199167 227702
rect 3969 227082 4035 227085
rect 170254 227082 170260 227084
rect 3969 227080 170260 227082
rect 3969 227024 3974 227080
rect 4030 227024 170260 227080
rect 3969 227022 170260 227024
rect 3969 227019 4035 227022
rect 170254 227020 170260 227022
rect 170324 227020 170330 227084
rect 3785 226946 3851 226949
rect 171542 226946 171548 226948
rect 3785 226944 171548 226946
rect 3785 226888 3790 226944
rect 3846 226888 171548 226944
rect 3785 226886 171548 226888
rect 3785 226883 3851 226886
rect 171542 226884 171548 226886
rect 171612 226884 171618 226948
rect 197537 226538 197603 226541
rect 198549 226538 198615 226541
rect 197537 226536 200032 226538
rect 197537 226480 197542 226536
rect 197598 226480 198554 226536
rect 198610 226480 200032 226536
rect 197537 226478 200032 226480
rect 197537 226475 197603 226478
rect 198549 226475 198615 226478
rect 198457 225314 198523 225317
rect 198457 225312 200032 225314
rect 198457 225256 198462 225312
rect 198518 225256 200032 225312
rect 198457 225254 200032 225256
rect 198457 225251 198523 225254
rect 197353 224090 197419 224093
rect 198641 224090 198707 224093
rect 197353 224088 200100 224090
rect 197353 224032 197358 224088
rect 197414 224032 198646 224088
rect 198702 224032 200100 224088
rect 197353 224030 200100 224032
rect 197353 224027 197419 224030
rect 198641 224027 198707 224030
rect 560201 223546 560267 223549
rect 556876 223544 560267 223546
rect 556876 223488 560206 223544
rect 560262 223488 560267 223544
rect 556876 223486 560267 223488
rect 560201 223483 560267 223486
rect 199561 222934 199627 222937
rect 199561 222932 200100 222934
rect 199561 222876 199566 222932
rect 199622 222876 200100 222932
rect 199561 222874 200100 222876
rect 199561 222871 199627 222874
rect 198917 221506 198983 221509
rect 198917 221504 200032 221506
rect 198917 221448 198922 221504
rect 198978 221448 200032 221504
rect 198917 221446 200032 221448
rect 198917 221443 198983 221446
rect 28441 221234 28507 221237
rect 28441 221232 29378 221234
rect 28441 221176 28446 221232
rect 28502 221220 29378 221232
rect 28502 221176 30032 221220
rect 28441 221174 30032 221176
rect 28441 221171 28507 221174
rect 29318 221160 30032 221174
rect 197353 220282 197419 220285
rect 198733 220282 198799 220285
rect 197353 220280 200032 220282
rect 197353 220224 197358 220280
rect 197414 220224 198738 220280
rect 198794 220224 200032 220280
rect 197353 220222 200032 220224
rect 197353 220219 197419 220222
rect 198733 220219 198799 220222
rect 197905 219058 197971 219061
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 197905 219056 200032 219058
rect 197905 219000 197910 219056
rect 197966 219000 200032 219056
rect 197905 218998 200032 219000
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 197905 218995 197971 218998
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect 197353 217834 197419 217837
rect 197353 217832 200032 217834
rect 197353 217776 197358 217832
rect 197414 217776 200032 217832
rect 197353 217774 200032 217776
rect 197353 217771 197419 217774
rect 197353 216610 197419 216613
rect 197353 216608 200032 216610
rect 197353 216552 197358 216608
rect 197414 216552 200032 216608
rect 197353 216550 200032 216552
rect 197353 216547 197419 216550
rect 559189 215658 559255 215661
rect 556876 215656 559255 215658
rect 556876 215600 559194 215656
rect 559250 215600 559255 215656
rect 556876 215598 559255 215600
rect 559189 215595 559255 215598
rect 198089 215386 198155 215389
rect 198089 215384 200100 215386
rect 198089 215328 198094 215384
rect 198150 215328 200100 215384
rect 198089 215326 200100 215328
rect 198089 215323 198155 215326
rect -960 214978 480 215068
rect 3969 214978 4035 214981
rect -960 214976 4035 214978
rect -960 214920 3974 214976
rect 4030 214920 4035 214976
rect -960 214918 4035 214920
rect -960 214828 480 214918
rect 3969 214915 4035 214918
rect 197353 214162 197419 214165
rect 197353 214160 200032 214162
rect 197353 214104 197358 214160
rect 197414 214104 200032 214160
rect 197353 214102 200032 214104
rect 197353 214099 197419 214102
rect 197353 212938 197419 212941
rect 197353 212936 200032 212938
rect 197353 212880 197358 212936
rect 197414 212880 200032 212936
rect 197353 212878 200032 212880
rect 197353 212875 197419 212878
rect 197629 211714 197695 211717
rect 197629 211712 200032 211714
rect 197629 211656 197634 211712
rect 197690 211656 200032 211712
rect 197629 211654 200032 211656
rect 197629 211651 197695 211654
rect 197353 210354 197419 210357
rect 197353 210352 200032 210354
rect 197353 210296 197358 210352
rect 197414 210296 200032 210352
rect 197353 210294 200032 210296
rect 197353 210291 197419 210294
rect 197721 209130 197787 209133
rect 197721 209128 200032 209130
rect 197721 209072 197726 209128
rect 197782 209072 200032 209128
rect 197721 209070 200032 209072
rect 197721 209067 197787 209070
rect 197353 208314 197419 208317
rect 197353 208312 200130 208314
rect 197353 208256 197358 208312
rect 197414 208256 200130 208312
rect 197353 208254 200130 208256
rect 197353 208251 197419 208254
rect 200070 207944 200130 208254
rect 560201 207634 560267 207637
rect 556876 207632 560267 207634
rect 556876 207576 560206 207632
rect 560262 207576 560267 207632
rect 556876 207574 560267 207576
rect 560201 207571 560267 207574
rect 197353 206682 197419 206685
rect 197353 206680 200032 206682
rect 197353 206624 197358 206680
rect 197414 206624 200032 206680
rect 197353 206622 200032 206624
rect 197353 206619 197419 206622
rect 580257 205730 580323 205733
rect 583520 205730 584960 205820
rect 580257 205728 584960 205730
rect 580257 205672 580262 205728
rect 580318 205672 584960 205728
rect 580257 205670 584960 205672
rect 580257 205667 580323 205670
rect 583520 205580 584960 205670
rect 197353 205458 197419 205461
rect 197353 205456 200032 205458
rect 197353 205400 197358 205456
rect 197414 205400 200032 205456
rect 197353 205398 200032 205400
rect 197353 205395 197419 205398
rect 197353 204234 197419 204237
rect 197353 204232 200032 204234
rect 197353 204176 197358 204232
rect 197414 204176 200032 204232
rect 197353 204174 200032 204176
rect 197353 204171 197419 204174
rect 197721 203010 197787 203013
rect 197721 203008 200032 203010
rect 197721 202952 197726 203008
rect 197782 202952 200032 203008
rect 197721 202950 200032 202952
rect 197721 202947 197787 202950
rect -960 201922 480 202012
rect 3601 201922 3667 201925
rect -960 201920 3667 201922
rect -960 201864 3606 201920
rect 3662 201864 3667 201920
rect -960 201862 3667 201864
rect -960 201772 480 201862
rect 3601 201859 3667 201862
rect 197353 201786 197419 201789
rect 197353 201784 200032 201786
rect 197353 201728 197358 201784
rect 197414 201728 200032 201784
rect 197353 201726 200032 201728
rect 197353 201723 197419 201726
rect 197353 200562 197419 200565
rect 197353 200560 200032 200562
rect 197353 200504 197358 200560
rect 197414 200504 200032 200560
rect 197353 200502 200032 200504
rect 197353 200499 197419 200502
rect 559557 199610 559623 199613
rect 556876 199608 559623 199610
rect 556876 199552 559562 199608
rect 559618 199552 559623 199608
rect 556876 199550 559623 199552
rect 559557 199547 559623 199550
rect 197353 199202 197419 199205
rect 197353 199200 200100 199202
rect 197353 199144 197358 199200
rect 197414 199144 200100 199200
rect 197353 199142 200100 199144
rect 197353 199139 197419 199142
rect 197353 197978 197419 197981
rect 197353 197976 200032 197978
rect 197353 197920 197358 197976
rect 197414 197920 200032 197976
rect 197353 197918 200032 197920
rect 197353 197915 197419 197918
rect 197353 196754 197419 196757
rect 197353 196752 200032 196754
rect 197353 196696 197358 196752
rect 197414 196696 200032 196752
rect 197353 196694 200032 196696
rect 197353 196691 197419 196694
rect 197353 195530 197419 195533
rect 197353 195528 200032 195530
rect 197353 195472 197358 195528
rect 197414 195472 200032 195528
rect 197353 195470 200032 195472
rect 197353 195467 197419 195470
rect 197353 194306 197419 194309
rect 197353 194304 200032 194306
rect 197353 194248 197358 194304
rect 197414 194248 200032 194304
rect 197353 194246 200032 194248
rect 197353 194243 197419 194246
rect 197353 193082 197419 193085
rect 197353 193080 200032 193082
rect 197353 193024 197358 193080
rect 197414 193024 200032 193080
rect 197353 193022 200032 193024
rect 197353 193019 197419 193022
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 197721 192402 197787 192405
rect 197721 192400 200130 192402
rect 197721 192344 197726 192400
rect 197782 192344 200130 192400
rect 583520 192388 584960 192478
rect 197721 192342 200130 192344
rect 197721 192339 197787 192342
rect 200070 191896 200130 192342
rect 560201 191722 560267 191725
rect 556876 191720 560267 191722
rect 556876 191664 560206 191720
rect 560262 191664 560267 191720
rect 556876 191662 560267 191664
rect 560201 191659 560267 191662
rect 197353 190634 197419 190637
rect 197353 190632 200032 190634
rect 197353 190576 197358 190632
rect 197414 190576 200032 190632
rect 197353 190574 200032 190576
rect 197353 190571 197419 190574
rect 197353 189410 197419 189413
rect 197353 189408 200032 189410
rect 197353 189352 197358 189408
rect 197414 189352 200032 189408
rect 197353 189350 200032 189352
rect 197353 189347 197419 189350
rect -960 188866 480 188956
rect 3877 188866 3943 188869
rect -960 188864 3943 188866
rect -960 188808 3882 188864
rect 3938 188808 3943 188864
rect -960 188806 3943 188808
rect -960 188716 480 188806
rect 3877 188803 3943 188806
rect 197353 188186 197419 188189
rect 197353 188184 200032 188186
rect 197353 188128 197358 188184
rect 197414 188128 200032 188184
rect 197353 188126 200032 188128
rect 197353 188123 197419 188126
rect 197353 186826 197419 186829
rect 197353 186824 200032 186826
rect 197353 186768 197358 186824
rect 197414 186768 200032 186824
rect 197353 186766 200032 186768
rect 197353 186763 197419 186766
rect 197353 185602 197419 185605
rect 197353 185600 200032 185602
rect 197353 185544 197358 185600
rect 197414 185544 200032 185600
rect 197353 185542 200032 185544
rect 197353 185539 197419 185542
rect 197353 184242 197419 184245
rect 200070 184242 200130 184344
rect 197353 184240 200130 184242
rect 197353 184184 197358 184240
rect 197414 184184 200130 184240
rect 197353 184182 200130 184184
rect 197353 184179 197419 184182
rect 560017 183698 560083 183701
rect 556876 183696 560083 183698
rect 556876 183640 560022 183696
rect 560078 183640 560083 183696
rect 556876 183638 560083 183640
rect 560017 183635 560083 183638
rect 197353 182882 197419 182885
rect 200070 182882 200130 183120
rect 197353 182880 200130 182882
rect 197353 182824 197358 182880
rect 197414 182824 200130 182880
rect 197353 182822 200130 182824
rect 197353 182819 197419 182822
rect 197353 181930 197419 181933
rect 197353 181928 200032 181930
rect 197353 181872 197358 181928
rect 197414 181872 200032 181928
rect 197353 181870 200032 181872
rect 197353 181867 197419 181870
rect 197353 180706 197419 180709
rect 197353 180704 200032 180706
rect 197353 180648 197358 180704
rect 197414 180648 200032 180704
rect 197353 180646 200032 180648
rect 197353 180643 197419 180646
rect 197353 179482 197419 179485
rect 197353 179480 200032 179482
rect 197353 179424 197358 179480
rect 197414 179424 200032 179480
rect 197353 179422 200032 179424
rect 197353 179419 197419 179422
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 168925 178938 168991 178941
rect 167134 178936 168991 178938
rect 167134 178924 168930 178936
rect 166612 178880 168930 178924
rect 168986 178880 168991 178936
rect 166612 178878 168991 178880
rect 166612 178864 167194 178878
rect 168925 178875 168991 178878
rect 197905 178258 197971 178261
rect 197905 178256 200032 178258
rect 197905 178200 197910 178256
rect 197966 178200 200032 178256
rect 197905 178198 200032 178200
rect 197905 178195 197971 178198
rect 169293 177986 169359 177989
rect 167134 177984 169359 177986
rect 167134 177972 169298 177984
rect 166612 177928 169298 177972
rect 169354 177928 169359 177984
rect 166612 177926 169359 177928
rect 166612 177912 167194 177926
rect 169293 177923 169359 177926
rect 197353 177034 197419 177037
rect 197353 177032 200032 177034
rect 197353 176976 197358 177032
rect 197414 176976 200032 177032
rect 197353 176974 200032 176976
rect 197353 176971 197419 176974
rect -960 175796 480 176036
rect 168925 175810 168991 175813
rect 167134 175808 168991 175810
rect 167134 175796 168930 175808
rect 166612 175752 168930 175796
rect 168986 175752 168991 175808
rect 166612 175750 168991 175752
rect 166612 175736 167194 175750
rect 168925 175747 168991 175750
rect 197353 175674 197419 175677
rect 560201 175674 560267 175677
rect 197353 175672 200032 175674
rect 197353 175616 197358 175672
rect 197414 175616 200032 175672
rect 197353 175614 200032 175616
rect 556876 175672 560267 175674
rect 556876 175616 560206 175672
rect 560262 175616 560267 175672
rect 556876 175614 560267 175616
rect 197353 175611 197419 175614
rect 560201 175611 560267 175614
rect 168833 174858 168899 174861
rect 167134 174856 168899 174858
rect 167134 174844 168838 174856
rect 166612 174800 168838 174844
rect 168894 174800 168899 174856
rect 166612 174798 168899 174800
rect 166612 174784 167194 174798
rect 168833 174795 168899 174798
rect 197353 174450 197419 174453
rect 197353 174448 200032 174450
rect 197353 174392 197358 174448
rect 197414 174392 200032 174448
rect 197353 174390 200032 174392
rect 197353 174387 197419 174390
rect 197353 173226 197419 173229
rect 197353 173224 200032 173226
rect 197353 173168 197358 173224
rect 197414 173168 200032 173224
rect 197353 173166 200032 173168
rect 197353 173163 197419 173166
rect 168741 173090 168807 173093
rect 167134 173088 168807 173090
rect 167134 173076 168746 173088
rect 166612 173032 168746 173076
rect 168802 173032 168807 173088
rect 166612 173030 168807 173032
rect 166612 173016 167194 173030
rect 168741 173027 168807 173030
rect 168925 172002 168991 172005
rect 167134 172000 168991 172002
rect 167134 171988 168930 172000
rect 166612 171944 168930 171988
rect 168986 171944 168991 172000
rect 166612 171942 168991 171944
rect 166612 171928 167194 171942
rect 168925 171939 168991 171942
rect 197353 172002 197419 172005
rect 197353 172000 200032 172002
rect 197353 171944 197358 172000
rect 197414 171944 200032 172000
rect 197353 171942 200032 171944
rect 197353 171939 197419 171942
rect 197353 170778 197419 170781
rect 197353 170776 200032 170778
rect 197353 170720 197358 170776
rect 197414 170720 200032 170776
rect 197353 170718 200032 170720
rect 197353 170715 197419 170718
rect 169109 170234 169175 170237
rect 167134 170232 169175 170234
rect 167134 170220 169114 170232
rect 166612 170176 169114 170220
rect 169170 170176 169175 170232
rect 166612 170174 169175 170176
rect 166612 170160 167194 170174
rect 169109 170171 169175 170174
rect 197353 169554 197419 169557
rect 197353 169552 200032 169554
rect 197353 169496 197358 169552
rect 197414 169496 200032 169552
rect 197353 169494 200032 169496
rect 197353 169491 197419 169494
rect 197353 167786 197419 167789
rect 200070 167786 200130 168296
rect 197353 167784 200130 167786
rect 197353 167728 197358 167784
rect 197414 167728 200130 167784
rect 197353 167726 200130 167728
rect 197353 167723 197419 167726
rect 197537 167650 197603 167653
rect 559005 167650 559071 167653
rect 197537 167648 200130 167650
rect 197537 167592 197542 167648
rect 197598 167592 200130 167648
rect 197537 167590 200130 167592
rect 556876 167648 559071 167650
rect 556876 167592 559010 167648
rect 559066 167592 559071 167648
rect 556876 167590 559071 167592
rect 197537 167587 197603 167590
rect 200070 167144 200130 167590
rect 559005 167587 559071 167590
rect 197353 165882 197419 165885
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 197353 165880 200032 165882
rect 197353 165824 197358 165880
rect 197414 165824 200032 165880
rect 197353 165822 200032 165824
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 197353 165819 197419 165822
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 197353 164522 197419 164525
rect 197353 164520 200032 164522
rect 197353 164464 197358 164520
rect 197414 164464 200032 164520
rect 197353 164462 200032 164464
rect 197353 164459 197419 164462
rect 197353 163298 197419 163301
rect 197353 163296 200032 163298
rect 197353 163240 197358 163296
rect 197414 163240 200032 163296
rect 197353 163238 200032 163240
rect 197353 163235 197419 163238
rect -960 162890 480 162980
rect 3785 162890 3851 162893
rect -960 162888 3851 162890
rect -960 162832 3790 162888
rect 3846 162832 3851 162888
rect -960 162830 3851 162832
rect -960 162740 480 162830
rect 3785 162827 3851 162830
rect 197353 162074 197419 162077
rect 197353 162072 200032 162074
rect 197353 162016 197358 162072
rect 197414 162016 200032 162072
rect 197353 162014 200032 162016
rect 197353 162011 197419 162014
rect 27153 161394 27219 161397
rect 27153 161392 29378 161394
rect 27153 161336 27158 161392
rect 27214 161380 29378 161392
rect 27214 161336 30032 161380
rect 27153 161334 30032 161336
rect 27153 161331 27219 161334
rect 29318 161320 30032 161334
rect 197353 160850 197419 160853
rect 197353 160848 200032 160850
rect 197353 160792 197358 160848
rect 197414 160792 200032 160848
rect 197353 160790 200032 160792
rect 197353 160787 197419 160790
rect 27153 160170 27219 160173
rect 27429 160170 27495 160173
rect 27153 160168 27495 160170
rect 27153 160112 27158 160168
rect 27214 160112 27434 160168
rect 27490 160112 27495 160168
rect 27153 160110 27495 160112
rect 27153 160107 27219 160110
rect 27429 160107 27495 160110
rect 27337 159762 27403 159765
rect 559557 159762 559623 159765
rect 27337 159760 29378 159762
rect 27337 159704 27342 159760
rect 27398 159748 29378 159760
rect 556876 159760 559623 159762
rect 27398 159704 30032 159748
rect 27337 159702 30032 159704
rect 556876 159704 559562 159760
rect 559618 159704 559623 159760
rect 556876 159702 559623 159704
rect 27337 159699 27403 159702
rect 29318 159688 30032 159702
rect 559557 159699 559623 159702
rect 197353 159490 197419 159493
rect 200070 159490 200130 159592
rect 197353 159488 200130 159490
rect 197353 159432 197358 159488
rect 197414 159432 200130 159488
rect 197353 159430 200130 159432
rect 197353 159427 197419 159430
rect 26969 158402 27035 158405
rect 27245 158402 27311 158405
rect 197353 158402 197419 158405
rect 26969 158400 29378 158402
rect 26969 158344 26974 158400
rect 27030 158344 27250 158400
rect 27306 158388 29378 158400
rect 197353 158400 200032 158402
rect 27306 158344 30032 158388
rect 26969 158342 30032 158344
rect 26969 158339 27035 158342
rect 27245 158339 27311 158342
rect 29318 158328 30032 158342
rect 197353 158344 197358 158400
rect 197414 158344 200032 158400
rect 197353 158342 200032 158344
rect 197353 158339 197419 158342
rect 197353 157178 197419 157181
rect 197353 157176 200032 157178
rect 197353 157120 197358 157176
rect 197414 157120 200032 157176
rect 197353 157118 200032 157120
rect 197353 157115 197419 157118
rect 27061 156906 27127 156909
rect 27061 156904 29378 156906
rect 27061 156848 27066 156904
rect 27122 156892 29378 156904
rect 27122 156848 30032 156892
rect 27061 156846 30032 156848
rect 27061 156843 27127 156846
rect 29318 156832 30032 156846
rect 197353 155954 197419 155957
rect 197353 155952 200032 155954
rect 197353 155896 197358 155952
rect 197414 155896 200032 155952
rect 197353 155894 200032 155896
rect 197353 155891 197419 155894
rect 27153 155682 27219 155685
rect 27521 155682 27587 155685
rect 27153 155680 29378 155682
rect 27153 155624 27158 155680
rect 27214 155624 27526 155680
rect 27582 155668 29378 155680
rect 27582 155624 30032 155668
rect 27153 155622 30032 155624
rect 27153 155619 27219 155622
rect 27521 155619 27587 155622
rect 29318 155608 30032 155622
rect 197537 154730 197603 154733
rect 197537 154728 200032 154730
rect 197537 154672 197542 154728
rect 197598 154672 200032 154728
rect 197537 154670 200032 154672
rect 197537 154667 197603 154670
rect 197353 153506 197419 153509
rect 197353 153504 200032 153506
rect 197353 153448 197358 153504
rect 197414 153448 200032 153504
rect 197353 153446 200032 153448
rect 197353 153443 197419 153446
rect 168373 153098 168439 153101
rect 169109 153098 169175 153101
rect 168373 153096 169175 153098
rect 168373 153040 168378 153096
rect 168434 153040 169114 153096
rect 169170 153040 169175 153096
rect 168373 153038 169175 153040
rect 168373 153035 168439 153038
rect 169109 153035 169175 153038
rect 197353 152826 197419 152829
rect 197353 152824 200130 152826
rect 197353 152768 197358 152824
rect 197414 152768 200130 152824
rect 197353 152766 200130 152768
rect 197353 152763 197419 152766
rect 200070 152184 200130 152766
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect 168373 152010 168439 152013
rect 167134 152008 168439 152010
rect 167134 151996 168378 152008
rect 166612 151952 168378 151996
rect 168434 151952 168439 152008
rect 166612 151950 168439 151952
rect 166612 151936 167194 151950
rect 168373 151947 168439 151950
rect 559557 151738 559623 151741
rect 556876 151736 559623 151738
rect 556876 151680 559562 151736
rect 559618 151680 559623 151736
rect 556876 151678 559623 151680
rect 559557 151675 559623 151678
rect 197353 150514 197419 150517
rect 200070 150514 200130 150888
rect 197353 150512 200130 150514
rect 197353 150456 197358 150512
rect 197414 150456 200130 150512
rect 197353 150454 200130 150456
rect 197353 150451 197419 150454
rect 168557 150378 168623 150381
rect 167134 150376 168623 150378
rect 167134 150364 168562 150376
rect 166612 150320 168562 150364
rect 168618 150320 168623 150376
rect 166612 150318 168623 150320
rect 166612 150304 167194 150318
rect 168557 150315 168623 150318
rect 168465 150106 168531 150109
rect 168741 150106 168807 150109
rect 167134 150104 168807 150106
rect 167134 150092 168470 150104
rect 166612 150048 168470 150092
rect 168526 150048 168746 150104
rect 168802 150048 168807 150104
rect 166612 150046 168807 150048
rect 166612 150032 167194 150046
rect 168465 150043 168531 150046
rect 168741 150043 168807 150046
rect -960 149834 480 149924
rect 3693 149834 3759 149837
rect -960 149832 3759 149834
rect -960 149776 3698 149832
rect 3754 149776 3759 149832
rect -960 149774 3759 149776
rect -960 149684 480 149774
rect 3693 149771 3759 149774
rect 197353 149698 197419 149701
rect 197353 149696 200032 149698
rect 197353 149640 197358 149696
rect 197414 149640 200032 149696
rect 197353 149638 200032 149640
rect 197353 149635 197419 149638
rect 197537 148474 197603 148477
rect 197537 148472 200032 148474
rect 197537 148416 197542 148472
rect 197598 148416 200032 148472
rect 197537 148414 200032 148416
rect 197537 148411 197603 148414
rect 197353 147250 197419 147253
rect 197353 147248 200032 147250
rect 197353 147192 197358 147248
rect 197414 147192 200032 147248
rect 197353 147190 200032 147192
rect 197353 147187 197419 147190
rect 197353 146026 197419 146029
rect 197353 146024 200032 146026
rect 197353 145968 197358 146024
rect 197414 145968 200032 146024
rect 197353 145966 200032 145968
rect 197353 145963 197419 145966
rect 197353 144802 197419 144805
rect 197353 144800 200032 144802
rect 197353 144744 197358 144800
rect 197414 144744 200032 144800
rect 197353 144742 200032 144744
rect 197353 144739 197419 144742
rect 560017 143714 560083 143717
rect 556876 143712 560083 143714
rect 556876 143656 560022 143712
rect 560078 143656 560083 143712
rect 556876 143654 560083 143656
rect 560017 143651 560083 143654
rect 197353 143578 197419 143581
rect 197353 143576 200100 143578
rect 197353 143520 197358 143576
rect 197414 143520 200100 143576
rect 197353 143518 200100 143520
rect 197353 143515 197419 143518
rect 197353 142354 197419 142357
rect 197353 142352 200032 142354
rect 197353 142296 197358 142352
rect 197414 142296 200032 142352
rect 197353 142294 200032 142296
rect 197353 142291 197419 142294
rect 122741 141810 122807 141813
rect 133137 141812 133203 141813
rect 123024 141810 123030 141812
rect 122696 141808 123030 141810
rect 122696 141752 122746 141808
rect 122802 141752 123030 141808
rect 122696 141750 123030 141752
rect 122741 141747 122807 141750
rect 123024 141748 123030 141750
rect 123094 141748 123100 141812
rect 133088 141810 133094 141812
rect 133046 141750 133094 141810
rect 133158 141808 133203 141812
rect 133198 141752 133203 141808
rect 133088 141748 133094 141750
rect 133158 141748 133203 141752
rect 133137 141747 133203 141748
rect 108481 141676 108547 141677
rect 112161 141676 112227 141677
rect 123753 141676 123819 141677
rect 128537 141676 128603 141677
rect 134241 141676 134307 141677
rect 136541 141676 136607 141677
rect 140037 141676 140103 141677
rect 142337 141676 142403 141677
rect 108472 141674 108478 141676
rect 108390 141614 108478 141674
rect 108472 141612 108478 141614
rect 108542 141612 108548 141676
rect 112144 141674 112150 141676
rect 112070 141614 112150 141674
rect 112214 141672 112227 141676
rect 123704 141674 123710 141676
rect 112222 141616 112227 141672
rect 112144 141612 112150 141614
rect 112214 141612 112227 141616
rect 123662 141614 123710 141674
rect 123774 141672 123819 141676
rect 128464 141674 128470 141676
rect 123814 141616 123819 141672
rect 123704 141612 123710 141614
rect 123774 141612 123819 141616
rect 128446 141614 128470 141674
rect 128464 141612 128470 141614
rect 128534 141672 128603 141676
rect 134176 141674 134182 141676
rect 128534 141616 128542 141672
rect 128598 141616 128603 141672
rect 128534 141612 128603 141616
rect 134150 141614 134182 141674
rect 134176 141612 134182 141614
rect 134246 141672 134307 141676
rect 136488 141674 136494 141676
rect 134302 141616 134307 141672
rect 134246 141612 134307 141616
rect 136450 141614 136494 141674
rect 136558 141672 136607 141676
rect 140024 141674 140030 141676
rect 136602 141616 136607 141672
rect 136488 141612 136494 141614
rect 136558 141612 136607 141616
rect 139946 141614 140030 141674
rect 140094 141672 140103 141676
rect 140098 141616 140103 141672
rect 140024 141612 140030 141614
rect 140094 141612 140103 141616
rect 142336 141612 142342 141676
rect 142406 141674 142412 141676
rect 142406 141614 142494 141674
rect 142406 141612 142412 141614
rect 108481 141611 108547 141612
rect 112161 141611 112227 141612
rect 123753 141611 123819 141612
rect 128537 141611 128603 141612
rect 134241 141611 134307 141612
rect 136541 141611 136607 141612
rect 140037 141611 140103 141612
rect 142337 141611 142403 141612
rect 197261 140994 197327 140997
rect 197261 140992 200032 140994
rect 197261 140936 197266 140992
rect 197322 140936 200032 140992
rect 197261 140934 200032 140936
rect 197261 140931 197327 140934
rect 109585 140724 109651 140725
rect 113265 140724 113331 140725
rect 116761 140724 116827 140725
rect 118969 140724 119035 140725
rect 125961 140724 126027 140725
rect 132033 140724 132099 140725
rect 135345 140724 135411 140725
rect 137921 140724 137987 140725
rect 139025 140724 139091 140725
rect 141233 140724 141299 140725
rect 143441 140724 143507 140725
rect 149513 140724 149579 140725
rect 109534 140722 109540 140724
rect 109494 140662 109540 140722
rect 109604 140720 109651 140724
rect 113214 140722 113220 140724
rect 109646 140664 109651 140720
rect 109534 140660 109540 140662
rect 109604 140660 109651 140664
rect 113174 140662 113220 140722
rect 113284 140720 113331 140724
rect 116710 140722 116716 140724
rect 113326 140664 113331 140720
rect 113214 140660 113220 140662
rect 113284 140660 113331 140664
rect 116670 140662 116716 140722
rect 116780 140720 116827 140724
rect 118918 140722 118924 140724
rect 116822 140664 116827 140720
rect 116710 140660 116716 140662
rect 116780 140660 116827 140664
rect 118878 140662 118924 140722
rect 118988 140720 119035 140724
rect 125910 140722 125916 140724
rect 119030 140664 119035 140720
rect 118918 140660 118924 140662
rect 118988 140660 119035 140664
rect 125870 140662 125916 140722
rect 125980 140720 126027 140724
rect 131982 140722 131988 140724
rect 126022 140664 126027 140720
rect 125910 140660 125916 140662
rect 125980 140660 126027 140664
rect 131942 140662 131988 140722
rect 132052 140720 132099 140724
rect 135294 140722 135300 140724
rect 132094 140664 132099 140720
rect 131982 140660 131988 140662
rect 132052 140660 132099 140664
rect 135254 140662 135300 140722
rect 135364 140720 135411 140724
rect 137870 140722 137876 140724
rect 135406 140664 135411 140720
rect 135294 140660 135300 140662
rect 135364 140660 135411 140664
rect 137830 140662 137876 140722
rect 137940 140720 137987 140724
rect 138974 140722 138980 140724
rect 137982 140664 137987 140720
rect 137870 140660 137876 140662
rect 137940 140660 137987 140664
rect 138934 140662 138980 140722
rect 139044 140720 139091 140724
rect 141182 140722 141188 140724
rect 139086 140664 139091 140720
rect 138974 140660 138980 140662
rect 139044 140660 139091 140664
rect 141142 140662 141188 140722
rect 141252 140720 141299 140724
rect 143390 140722 143396 140724
rect 141294 140664 141299 140720
rect 141182 140660 141188 140662
rect 141252 140660 141299 140664
rect 143350 140662 143396 140722
rect 143460 140720 143507 140724
rect 149462 140722 149468 140724
rect 143502 140664 143507 140720
rect 143390 140660 143396 140662
rect 143460 140660 143507 140664
rect 149422 140662 149468 140722
rect 149532 140720 149579 140724
rect 149574 140664 149579 140720
rect 149462 140660 149468 140662
rect 149532 140660 149579 140664
rect 109585 140659 109651 140660
rect 113265 140659 113331 140660
rect 116761 140659 116827 140660
rect 118969 140659 119035 140660
rect 125961 140659 126027 140660
rect 132033 140659 132099 140660
rect 135345 140659 135411 140660
rect 137921 140659 137987 140660
rect 139025 140659 139091 140660
rect 141233 140659 141299 140660
rect 143441 140659 143507 140660
rect 149513 140659 149579 140660
rect 43069 140180 43135 140181
rect 63217 140180 63283 140181
rect 65793 140180 65859 140181
rect 115473 140180 115539 140181
rect 43069 140176 43116 140180
rect 43180 140178 43186 140180
rect 63166 140178 63172 140180
rect 43069 140120 43074 140176
rect 43069 140116 43116 140120
rect 43180 140118 43226 140178
rect 63126 140118 63172 140178
rect 63236 140176 63283 140180
rect 65742 140178 65748 140180
rect 63278 140120 63283 140176
rect 43180 140116 43186 140118
rect 63166 140116 63172 140118
rect 63236 140116 63283 140120
rect 65702 140118 65748 140178
rect 65812 140176 65859 140180
rect 115422 140178 115428 140180
rect 65854 140120 65859 140176
rect 65742 140116 65748 140118
rect 65812 140116 65859 140120
rect 115382 140118 115428 140178
rect 115492 140176 115539 140180
rect 115534 140120 115539 140176
rect 115422 140116 115428 140118
rect 115492 140116 115539 140120
rect 115606 140116 115612 140180
rect 115676 140178 115682 140180
rect 115841 140178 115907 140181
rect 129641 140180 129707 140181
rect 129590 140178 129596 140180
rect 115676 140176 115907 140178
rect 115676 140120 115846 140176
rect 115902 140120 115907 140176
rect 115676 140118 115907 140120
rect 129550 140118 129596 140178
rect 129660 140176 129707 140180
rect 129702 140120 129707 140176
rect 115676 140116 115682 140118
rect 43069 140115 43135 140116
rect 63217 140115 63283 140116
rect 65793 140115 65859 140116
rect 115473 140115 115539 140116
rect 115841 140115 115907 140118
rect 129590 140116 129596 140118
rect 129660 140116 129707 140120
rect 129641 140115 129707 140116
rect 197353 139770 197419 139773
rect 197353 139768 200032 139770
rect 197353 139712 197358 139768
rect 197414 139712 200032 139768
rect 197353 139710 200032 139712
rect 197353 139707 197419 139710
rect 43437 139362 43503 139365
rect 60641 139364 60707 139365
rect 107377 139364 107443 139365
rect 110873 139364 110939 139365
rect 114369 139364 114435 139365
rect 117865 139364 117931 139365
rect 43662 139362 43668 139364
rect 43437 139360 43668 139362
rect 43437 139304 43442 139360
rect 43498 139304 43668 139360
rect 43437 139302 43668 139304
rect 43437 139299 43503 139302
rect 43662 139300 43668 139302
rect 43732 139300 43738 139364
rect 60590 139362 60596 139364
rect 60550 139302 60596 139362
rect 60660 139360 60707 139364
rect 107326 139362 107332 139364
rect 60702 139304 60707 139360
rect 60590 139300 60596 139302
rect 60660 139300 60707 139304
rect 107286 139302 107332 139362
rect 107396 139360 107443 139364
rect 110822 139362 110828 139364
rect 107438 139304 107443 139360
rect 107326 139300 107332 139302
rect 107396 139300 107443 139304
rect 110782 139302 110828 139362
rect 110892 139360 110939 139364
rect 114318 139362 114324 139364
rect 110934 139304 110939 139360
rect 110822 139300 110828 139302
rect 110892 139300 110939 139304
rect 114278 139302 114324 139362
rect 114388 139360 114435 139364
rect 117814 139362 117820 139364
rect 114430 139304 114435 139360
rect 114318 139300 114324 139302
rect 114388 139300 114435 139304
rect 117774 139302 117820 139362
rect 117884 139360 117931 139364
rect 117926 139304 117931 139360
rect 117814 139300 117820 139302
rect 117884 139300 117931 139304
rect 120206 139300 120212 139364
rect 120276 139362 120282 139364
rect 120349 139362 120415 139365
rect 121361 139364 121427 139365
rect 122649 139364 122715 139365
rect 121310 139362 121316 139364
rect 120276 139360 120415 139362
rect 120276 139304 120354 139360
rect 120410 139304 120415 139360
rect 120276 139302 120415 139304
rect 121270 139302 121316 139362
rect 121380 139360 121427 139364
rect 122598 139362 122604 139364
rect 121422 139304 121427 139360
rect 120276 139300 120282 139302
rect 60641 139299 60707 139300
rect 107377 139299 107443 139300
rect 110873 139299 110939 139300
rect 114369 139299 114435 139300
rect 117865 139299 117931 139300
rect 120349 139299 120415 139302
rect 121310 139300 121316 139302
rect 121380 139300 121427 139304
rect 122558 139302 122604 139362
rect 122668 139360 122715 139364
rect 122710 139304 122715 139360
rect 122598 139300 122604 139302
rect 122668 139300 122715 139304
rect 124806 139300 124812 139364
rect 124876 139362 124882 139364
rect 125225 139362 125291 139365
rect 124876 139360 125291 139362
rect 124876 139304 125230 139360
rect 125286 139304 125291 139360
rect 124876 139302 125291 139304
rect 124876 139300 124882 139302
rect 121361 139299 121427 139300
rect 122649 139299 122715 139300
rect 125225 139299 125291 139302
rect 127198 139300 127204 139364
rect 127268 139362 127274 139364
rect 127709 139362 127775 139365
rect 130745 139364 130811 139365
rect 148409 139364 148475 139365
rect 130694 139362 130700 139364
rect 127268 139360 127775 139362
rect 127268 139304 127714 139360
rect 127770 139304 127775 139360
rect 127268 139302 127775 139304
rect 130654 139302 130700 139362
rect 130764 139360 130811 139364
rect 148358 139362 148364 139364
rect 130806 139304 130811 139360
rect 127268 139300 127274 139302
rect 127709 139299 127775 139302
rect 130694 139300 130700 139302
rect 130764 139300 130811 139304
rect 148318 139302 148364 139362
rect 148428 139360 148475 139364
rect 148470 139304 148475 139360
rect 148358 139300 148364 139302
rect 148428 139300 148475 139304
rect 150566 139300 150572 139364
rect 150636 139362 150642 139364
rect 151077 139362 151143 139365
rect 150636 139360 151143 139362
rect 150636 139304 151082 139360
rect 151138 139304 151143 139360
rect 150636 139302 151143 139304
rect 150636 139300 150642 139302
rect 130745 139299 130811 139300
rect 148409 139299 148475 139300
rect 151077 139299 151143 139302
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 136214 139028 136220 139092
rect 136284 139090 136290 139092
rect 136449 139090 136515 139093
rect 136284 139088 136515 139090
rect 136284 139032 136454 139088
rect 136510 139032 136515 139088
rect 136284 139030 136515 139032
rect 136284 139028 136290 139030
rect 136449 139027 136515 139030
rect 68134 138620 68140 138684
rect 68204 138682 68210 138684
rect 68921 138682 68987 138685
rect 68204 138680 68987 138682
rect 68204 138624 68926 138680
rect 68982 138624 68987 138680
rect 68204 138622 68987 138624
rect 68204 138620 68210 138622
rect 68921 138619 68987 138622
rect 122741 138682 122807 138685
rect 124121 138682 124187 138685
rect 122741 138680 124187 138682
rect 122741 138624 122746 138680
rect 122802 138624 124126 138680
rect 124182 138624 124187 138680
rect 122741 138622 124187 138624
rect 122741 138619 122807 138622
rect 124121 138619 124187 138622
rect 197445 138546 197511 138549
rect 197445 138544 200032 138546
rect 197445 138488 197450 138544
rect 197506 138488 200032 138544
rect 197445 138486 200032 138488
rect 197445 138483 197511 138486
rect 70710 138076 70716 138140
rect 70780 138138 70786 138140
rect 71037 138138 71103 138141
rect 70780 138136 71103 138138
rect 70780 138080 71042 138136
rect 71098 138080 71103 138136
rect 70780 138078 71103 138080
rect 70780 138076 70786 138078
rect 71037 138075 71103 138078
rect 73654 138076 73660 138140
rect 73724 138138 73730 138140
rect 74441 138138 74507 138141
rect 73724 138136 74507 138138
rect 73724 138080 74446 138136
rect 74502 138080 74507 138136
rect 73724 138078 74507 138080
rect 73724 138076 73730 138078
rect 74441 138075 74507 138078
rect 75310 138076 75316 138140
rect 75380 138138 75386 138140
rect 75821 138138 75887 138141
rect 75380 138136 75887 138138
rect 75380 138080 75826 138136
rect 75882 138080 75887 138136
rect 75380 138078 75887 138080
rect 75380 138076 75386 138078
rect 75821 138075 75887 138078
rect 78070 138076 78076 138140
rect 78140 138138 78146 138140
rect 78581 138138 78647 138141
rect 78140 138136 78647 138138
rect 78140 138080 78586 138136
rect 78642 138080 78647 138136
rect 78140 138078 78647 138080
rect 78140 138076 78146 138078
rect 78581 138075 78647 138078
rect 80646 138076 80652 138140
rect 80716 138138 80722 138140
rect 81341 138138 81407 138141
rect 80716 138136 81407 138138
rect 80716 138080 81346 138136
rect 81402 138080 81407 138136
rect 80716 138078 81407 138080
rect 80716 138076 80722 138078
rect 81341 138075 81407 138078
rect 83774 138076 83780 138140
rect 83844 138138 83850 138140
rect 84101 138138 84167 138141
rect 83844 138136 84167 138138
rect 83844 138080 84106 138136
rect 84162 138080 84167 138136
rect 83844 138078 84167 138080
rect 83844 138076 83850 138078
rect 84101 138075 84167 138078
rect 86350 138076 86356 138140
rect 86420 138138 86426 138140
rect 86861 138138 86927 138141
rect 88241 138140 88307 138141
rect 88190 138138 88196 138140
rect 86420 138136 86927 138138
rect 86420 138080 86866 138136
rect 86922 138080 86927 138136
rect 86420 138078 86927 138080
rect 88150 138078 88196 138138
rect 88260 138136 88307 138140
rect 88302 138080 88307 138136
rect 86420 138076 86426 138078
rect 86861 138075 86927 138078
rect 88190 138076 88196 138078
rect 88260 138076 88307 138080
rect 90766 138076 90772 138140
rect 90836 138138 90842 138140
rect 91001 138138 91067 138141
rect 93761 138140 93827 138141
rect 93710 138138 93716 138140
rect 90836 138136 91067 138138
rect 90836 138080 91006 138136
rect 91062 138080 91067 138136
rect 90836 138078 91067 138080
rect 93670 138078 93716 138138
rect 93780 138136 93827 138140
rect 93822 138080 93827 138136
rect 90836 138076 90842 138078
rect 88241 138075 88307 138076
rect 91001 138075 91067 138078
rect 93710 138076 93716 138078
rect 93780 138076 93827 138080
rect 96286 138076 96292 138140
rect 96356 138138 96362 138140
rect 96521 138138 96587 138141
rect 96356 138136 96587 138138
rect 96356 138080 96526 138136
rect 96582 138080 96587 138136
rect 96356 138078 96587 138080
rect 96356 138076 96362 138078
rect 93761 138075 93827 138076
rect 96521 138075 96587 138078
rect 98310 138076 98316 138140
rect 98380 138138 98386 138140
rect 99281 138138 99347 138141
rect 98380 138136 99347 138138
rect 98380 138080 99286 138136
rect 99342 138080 99347 138136
rect 98380 138078 99347 138080
rect 98380 138076 98386 138078
rect 99281 138075 99347 138078
rect 100518 138076 100524 138140
rect 100588 138138 100594 138140
rect 100661 138138 100727 138141
rect 100588 138136 100727 138138
rect 100588 138080 100666 138136
rect 100722 138080 100727 138136
rect 100588 138078 100727 138080
rect 100588 138076 100594 138078
rect 100661 138075 100727 138078
rect 102726 138076 102732 138140
rect 102796 138138 102802 138140
rect 103421 138138 103487 138141
rect 102796 138136 103487 138138
rect 102796 138080 103426 138136
rect 103482 138080 103487 138136
rect 102796 138078 103487 138080
rect 102796 138076 102802 138078
rect 103421 138075 103487 138078
rect 105302 138076 105308 138140
rect 105372 138138 105378 138140
rect 106181 138138 106247 138141
rect 105372 138136 106247 138138
rect 105372 138080 106186 138136
rect 106242 138080 106247 138136
rect 105372 138078 106247 138080
rect 105372 138076 105378 138078
rect 106181 138075 106247 138078
rect 108062 138076 108068 138140
rect 108132 138138 108138 138140
rect 108941 138138 109007 138141
rect 108132 138136 109007 138138
rect 108132 138080 108946 138136
rect 109002 138080 109007 138136
rect 108132 138078 109007 138080
rect 108132 138076 108138 138078
rect 108941 138075 109007 138078
rect 110454 138076 110460 138140
rect 110524 138138 110530 138140
rect 111701 138138 111767 138141
rect 110524 138136 111767 138138
rect 110524 138080 111706 138136
rect 111762 138080 111767 138136
rect 110524 138078 111767 138080
rect 110524 138076 110530 138078
rect 111701 138075 111767 138078
rect 112662 138076 112668 138140
rect 112732 138138 112738 138140
rect 113081 138138 113147 138141
rect 118417 138140 118483 138141
rect 118366 138138 118372 138140
rect 112732 138136 113147 138138
rect 112732 138080 113086 138136
rect 113142 138080 113147 138136
rect 112732 138078 113147 138080
rect 118326 138078 118372 138138
rect 118436 138136 118483 138140
rect 118478 138080 118483 138136
rect 112732 138076 112738 138078
rect 113081 138075 113147 138078
rect 118366 138076 118372 138078
rect 118436 138076 118483 138080
rect 120574 138076 120580 138140
rect 120644 138138 120650 138140
rect 121361 138138 121427 138141
rect 125409 138140 125475 138141
rect 125358 138138 125364 138140
rect 120644 138136 121427 138138
rect 120644 138080 121366 138136
rect 121422 138080 121427 138136
rect 120644 138078 121427 138080
rect 125318 138078 125364 138138
rect 125428 138136 125475 138140
rect 125470 138080 125475 138136
rect 120644 138076 120650 138078
rect 118417 138075 118483 138076
rect 121361 138075 121427 138078
rect 125358 138076 125364 138078
rect 125428 138076 125475 138080
rect 128118 138076 128124 138140
rect 128188 138138 128194 138140
rect 128261 138138 128327 138141
rect 128188 138136 128327 138138
rect 128188 138080 128266 138136
rect 128322 138080 128327 138136
rect 128188 138078 128327 138080
rect 128188 138076 128194 138078
rect 125409 138075 125475 138076
rect 128261 138075 128327 138078
rect 130510 138076 130516 138140
rect 130580 138138 130586 138140
rect 131021 138138 131087 138141
rect 130580 138136 131087 138138
rect 130580 138080 131026 138136
rect 131082 138080 131087 138136
rect 130580 138078 131087 138080
rect 130580 138076 130586 138078
rect 131021 138075 131087 138078
rect 132718 138076 132724 138140
rect 132788 138138 132794 138140
rect 133781 138138 133847 138141
rect 132788 138136 133847 138138
rect 132788 138080 133786 138136
rect 133842 138080 133847 138136
rect 132788 138078 133847 138080
rect 132788 138076 132794 138078
rect 133781 138075 133847 138078
rect 138238 138076 138244 138140
rect 138308 138138 138314 138140
rect 139301 138138 139367 138141
rect 138308 138136 139367 138138
rect 138308 138080 139306 138136
rect 139362 138080 139367 138136
rect 138308 138078 139367 138080
rect 138308 138076 138314 138078
rect 139301 138075 139367 138078
rect 197353 137322 197419 137325
rect 197353 137320 200032 137322
rect 197353 137264 197358 137320
rect 197414 137264 200032 137320
rect 197353 137262 200032 137264
rect 197353 137259 197419 137262
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 197353 136370 197419 136373
rect 197353 136368 200130 136370
rect 197353 136312 197358 136368
rect 197414 136312 200130 136368
rect 197353 136310 200130 136312
rect 197353 136307 197419 136310
rect 200070 136136 200130 136310
rect 559281 135826 559347 135829
rect 556876 135824 559347 135826
rect 556876 135768 559286 135824
rect 559342 135768 559347 135824
rect 556876 135766 559347 135768
rect 559281 135763 559347 135766
rect 197353 134874 197419 134877
rect 197353 134872 200032 134874
rect 197353 134816 197358 134872
rect 197414 134816 200032 134872
rect 197353 134814 200032 134816
rect 197353 134811 197419 134814
rect 197353 133650 197419 133653
rect 197353 133648 200032 133650
rect 197353 133592 197358 133648
rect 197414 133592 200032 133648
rect 197353 133590 200032 133592
rect 197353 133587 197419 133590
rect 197353 132426 197419 132429
rect 197353 132424 200032 132426
rect 197353 132368 197358 132424
rect 197414 132368 200032 132424
rect 197353 132366 200032 132368
rect 197353 132363 197419 132366
rect 197445 131202 197511 131205
rect 197445 131200 200032 131202
rect 197445 131144 197450 131200
rect 197506 131144 200032 131200
rect 197445 131142 200032 131144
rect 197445 131139 197511 131142
rect 197353 129842 197419 129845
rect 197353 129840 200032 129842
rect 197353 129784 197358 129840
rect 197414 129784 200032 129840
rect 197353 129782 200032 129784
rect 197353 129779 197419 129782
rect 197353 129298 197419 129301
rect 197353 129296 200130 129298
rect 197353 129240 197358 129296
rect 197414 129240 200130 129296
rect 197353 129238 200130 129240
rect 197353 129235 197419 129238
rect 200070 128656 200130 129238
rect 197353 128074 197419 128077
rect 197353 128072 200130 128074
rect 197353 128016 197358 128072
rect 197414 128016 200130 128072
rect 197353 128014 200130 128016
rect 197353 128011 197419 128014
rect 200070 127432 200130 128014
rect 559557 127802 559623 127805
rect 556876 127800 559623 127802
rect 556876 127744 559562 127800
rect 559618 127744 559623 127800
rect 556876 127742 559623 127744
rect 559557 127739 559623 127742
rect 197353 126170 197419 126173
rect 197353 126168 200032 126170
rect 197353 126112 197358 126168
rect 197414 126112 200032 126168
rect 197353 126110 200032 126112
rect 197353 126107 197419 126110
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 197353 124946 197419 124949
rect 197353 124944 200032 124946
rect 197353 124888 197358 124944
rect 197414 124888 200032 124944
rect 197353 124886 200032 124888
rect 197353 124883 197419 124886
rect -960 123572 480 123812
rect 197353 123722 197419 123725
rect 197353 123720 200032 123722
rect 197353 123664 197358 123720
rect 197414 123664 200032 123720
rect 197353 123662 200032 123664
rect 197353 123659 197419 123662
rect 197353 122498 197419 122501
rect 197353 122496 200032 122498
rect 197353 122440 197358 122496
rect 197414 122440 200032 122496
rect 197353 122438 200032 122440
rect 197353 122435 197419 122438
rect 197353 121274 197419 121277
rect 197353 121272 200032 121274
rect 197353 121216 197358 121272
rect 197414 121216 200032 121272
rect 197353 121214 200032 121216
rect 197353 121211 197419 121214
rect 197353 120050 197419 120053
rect 197353 120048 200100 120050
rect 197353 119992 197358 120048
rect 197414 119992 200100 120048
rect 197353 119990 200100 119992
rect 197353 119987 197419 119990
rect 558913 119778 558979 119781
rect 556876 119776 558979 119778
rect 556876 119720 558918 119776
rect 558974 119720 558979 119776
rect 556876 119718 558979 119720
rect 558913 119715 558979 119718
rect 197445 118826 197511 118829
rect 197445 118824 200032 118826
rect 197445 118768 197450 118824
rect 197506 118768 200032 118824
rect 197445 118766 200032 118768
rect 197445 118763 197511 118766
rect 197353 117466 197419 117469
rect 197353 117464 200032 117466
rect 197353 117408 197358 117464
rect 197414 117408 200032 117464
rect 197353 117406 200032 117408
rect 197353 117403 197419 117406
rect 35198 117132 35204 117196
rect 35268 117194 35274 117196
rect 35801 117194 35867 117197
rect 35268 117192 35867 117194
rect 35268 117136 35806 117192
rect 35862 117136 35867 117192
rect 35268 117134 35867 117136
rect 35268 117132 35274 117134
rect 35801 117131 35867 117134
rect 45829 117058 45895 117061
rect 46790 117058 46796 117060
rect 45829 117056 46796 117058
rect 45829 117000 45834 117056
rect 45890 117000 46796 117056
rect 45829 116998 46796 117000
rect 45829 116995 45895 116998
rect 46790 116996 46796 116998
rect 46860 116996 46866 117060
rect 46933 116786 46999 116789
rect 48078 116786 48084 116788
rect 46933 116784 48084 116786
rect 46933 116728 46938 116784
rect 46994 116728 48084 116784
rect 46933 116726 48084 116728
rect 46933 116723 46999 116726
rect 48078 116724 48084 116726
rect 48148 116724 48154 116788
rect 197353 116242 197419 116245
rect 197353 116240 200032 116242
rect 197353 116184 197358 116240
rect 197414 116184 200032 116240
rect 197353 116182 200032 116184
rect 197353 116179 197419 116182
rect 197353 115018 197419 115021
rect 197353 115016 200032 115018
rect 197353 114960 197358 115016
rect 197414 114960 200032 115016
rect 197353 114958 200032 114960
rect 197353 114955 197419 114958
rect 197353 113794 197419 113797
rect 197353 113792 200032 113794
rect 197353 113736 197358 113792
rect 197414 113736 200032 113792
rect 197353 113734 200032 113736
rect 197353 113731 197419 113734
rect 197353 113114 197419 113117
rect 197353 113112 200130 113114
rect 197353 113056 197358 113112
rect 197414 113056 200130 113112
rect 197353 113054 200130 113056
rect 197353 113051 197419 113054
rect 200070 112608 200130 113054
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 559189 111890 559255 111893
rect 556876 111888 559255 111890
rect 556876 111832 559194 111888
rect 559250 111832 559255 111888
rect 556876 111830 559255 111832
rect 559189 111827 559255 111830
rect 197353 111754 197419 111757
rect 197353 111752 200130 111754
rect 197353 111696 197358 111752
rect 197414 111696 200130 111752
rect 197353 111694 200130 111696
rect 197353 111691 197419 111694
rect 200070 111384 200130 111694
rect -960 110666 480 110756
rect 4061 110666 4127 110669
rect -960 110664 4127 110666
rect -960 110608 4066 110664
rect 4122 110608 4127 110664
rect -960 110606 4127 110608
rect -960 110516 480 110606
rect 4061 110603 4127 110606
rect 197353 110122 197419 110125
rect 197353 110120 200032 110122
rect 197353 110064 197358 110120
rect 197414 110064 200032 110120
rect 197353 110062 200032 110064
rect 197353 110059 197419 110062
rect 28901 109306 28967 109309
rect 28901 109304 29378 109306
rect 28901 109248 28906 109304
rect 28962 109248 29378 109304
rect 28901 109246 29378 109248
rect 28901 109243 28967 109246
rect 29318 109220 29378 109246
rect 29318 109160 30032 109220
rect 197353 108898 197419 108901
rect 197353 108896 200032 108898
rect 197353 108840 197358 108896
rect 197414 108840 200032 108896
rect 197353 108838 200032 108840
rect 197353 108835 197419 108838
rect 197537 107674 197603 107677
rect 197537 107672 200032 107674
rect 197537 107616 197542 107672
rect 197598 107616 200032 107672
rect 197537 107614 200032 107616
rect 197537 107611 197603 107614
rect 197445 106314 197511 106317
rect 197445 106312 200032 106314
rect 197445 106256 197450 106312
rect 197506 106256 200032 106312
rect 197445 106254 200032 106256
rect 197445 106251 197511 106254
rect 197353 105090 197419 105093
rect 197353 105088 200032 105090
rect 197353 105032 197358 105088
rect 197414 105032 200032 105088
rect 197353 105030 200032 105032
rect 197353 105027 197419 105030
rect 197353 103866 197419 103869
rect 560201 103866 560267 103869
rect 197353 103864 200032 103866
rect 197353 103808 197358 103864
rect 197414 103808 200032 103864
rect 197353 103806 200032 103808
rect 556876 103864 560267 103866
rect 556876 103808 560206 103864
rect 560262 103808 560267 103864
rect 556876 103806 560267 103808
rect 197353 103803 197419 103806
rect 560201 103803 560267 103806
rect 197353 102642 197419 102645
rect 197353 102640 200032 102642
rect 197353 102584 197358 102640
rect 197414 102584 200032 102640
rect 197353 102582 200032 102584
rect 197353 102579 197419 102582
rect 197353 101418 197419 101421
rect 197353 101416 200032 101418
rect 197353 101360 197358 101416
rect 197414 101360 200032 101416
rect 197353 101358 200032 101360
rect 197353 101355 197419 101358
rect 197353 100194 197419 100197
rect 197353 100192 200032 100194
rect 197353 100136 197358 100192
rect 197414 100136 200032 100192
rect 197353 100134 200032 100136
rect 197353 100131 197419 100134
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 197353 98970 197419 98973
rect 197353 98968 200032 98970
rect 197353 98912 197358 98968
rect 197414 98912 200032 98968
rect 197353 98910 200032 98912
rect 197353 98907 197419 98910
rect 197997 97746 198063 97749
rect 197997 97744 200032 97746
rect -960 97610 480 97700
rect 197997 97688 198002 97744
rect 198058 97688 200032 97744
rect 197997 97686 200032 97688
rect 197997 97683 198063 97686
rect 3877 97610 3943 97613
rect -960 97608 3943 97610
rect -960 97552 3882 97608
rect 3938 97552 3943 97608
rect -960 97550 3943 97552
rect -960 97460 480 97550
rect 3877 97547 3943 97550
rect 198089 95978 198155 95981
rect 200070 95978 200130 96488
rect 198089 95976 200130 95978
rect 198089 95920 198094 95976
rect 198150 95920 200130 95976
rect 198089 95918 200130 95920
rect 198089 95915 198155 95918
rect 559741 95842 559807 95845
rect 556876 95840 559807 95842
rect 556876 95784 559746 95840
rect 559802 95784 559807 95840
rect 556876 95782 559807 95784
rect 559741 95779 559807 95782
rect 197353 94618 197419 94621
rect 200070 94618 200130 95128
rect 197353 94616 200130 94618
rect 197353 94560 197358 94616
rect 197414 94560 200130 94616
rect 197353 94558 200130 94560
rect 197353 94555 197419 94558
rect 198181 93938 198247 93941
rect 198181 93936 200032 93938
rect 198181 93880 198186 93936
rect 198242 93880 200032 93936
rect 198181 93878 200032 93880
rect 198181 93875 198247 93878
rect 197353 92714 197419 92717
rect 197353 92712 200032 92714
rect 197353 92656 197358 92712
rect 197414 92656 200032 92712
rect 197353 92654 200032 92656
rect 197353 92651 197419 92654
rect 197353 91490 197419 91493
rect 197353 91488 200032 91490
rect 197353 91432 197358 91488
rect 197414 91432 200032 91488
rect 197353 91430 200032 91432
rect 197353 91427 197419 91430
rect 197353 90266 197419 90269
rect 197353 90264 200032 90266
rect 197353 90208 197358 90264
rect 197414 90208 200032 90264
rect 197353 90206 200032 90208
rect 197353 90203 197419 90206
rect 197353 89042 197419 89045
rect 197353 89040 200032 89042
rect 197353 88984 197358 89040
rect 197414 88984 200032 89040
rect 197353 88982 200032 88984
rect 197353 88979 197419 88982
rect 560201 87954 560267 87957
rect 556876 87952 560267 87954
rect 556876 87896 560206 87952
rect 560262 87896 560267 87952
rect 556876 87894 560267 87896
rect 560201 87891 560267 87894
rect 197353 87274 197419 87277
rect 200070 87274 200130 87784
rect 197353 87272 200130 87274
rect 197353 87216 197358 87272
rect 197414 87216 200130 87272
rect 197353 87214 200130 87216
rect 197353 87211 197419 87214
rect 197353 86594 197419 86597
rect 197353 86592 200032 86594
rect 197353 86536 197358 86592
rect 197414 86536 200032 86592
rect 197353 86534 200032 86536
rect 197353 86531 197419 86534
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 197353 85370 197419 85373
rect 197353 85368 200032 85370
rect 197353 85312 197358 85368
rect 197414 85312 200032 85368
rect 197353 85310 200032 85312
rect 197353 85307 197419 85310
rect -960 84690 480 84780
rect 3785 84690 3851 84693
rect -960 84688 3851 84690
rect -960 84632 3790 84688
rect 3846 84632 3851 84688
rect -960 84630 3851 84632
rect -960 84540 480 84630
rect 3785 84627 3851 84630
rect 197353 84146 197419 84149
rect 197353 84144 200032 84146
rect 197353 84088 197358 84144
rect 197414 84088 200032 84144
rect 197353 84086 200032 84088
rect 197353 84083 197419 84086
rect 197445 82786 197511 82789
rect 197445 82784 200032 82786
rect 197445 82728 197450 82784
rect 197506 82728 200032 82784
rect 197445 82726 200032 82728
rect 197445 82723 197511 82726
rect 197353 81562 197419 81565
rect 197353 81560 200032 81562
rect 197353 81504 197358 81560
rect 197414 81504 200032 81560
rect 197353 81502 200032 81504
rect 197353 81499 197419 81502
rect 197353 80202 197419 80205
rect 200070 80202 200130 80304
rect 197353 80200 200130 80202
rect 197353 80144 197358 80200
rect 197414 80144 200130 80200
rect 197353 80142 200130 80144
rect 197353 80139 197419 80142
rect 560017 79930 560083 79933
rect 556876 79928 560083 79930
rect 556876 79872 560022 79928
rect 560078 79872 560083 79928
rect 556876 79870 560083 79872
rect 560017 79867 560083 79870
rect 197353 78842 197419 78845
rect 200070 78842 200130 79080
rect 197353 78840 200130 78842
rect 197353 78784 197358 78840
rect 197414 78784 200130 78840
rect 197353 78782 200130 78784
rect 197353 78779 197419 78782
rect 197353 77890 197419 77893
rect 197353 77888 200032 77890
rect 197353 77832 197358 77888
rect 197414 77832 200032 77888
rect 197353 77830 200032 77832
rect 197353 77827 197419 77830
rect 197353 76666 197419 76669
rect 197353 76664 200032 76666
rect 197353 76608 197358 76664
rect 197414 76608 200032 76664
rect 197353 76606 200032 76608
rect 197353 76603 197419 76606
rect 197353 75442 197419 75445
rect 197353 75440 200032 75442
rect 197353 75384 197358 75440
rect 197414 75384 200032 75440
rect 197353 75382 200032 75384
rect 197353 75379 197419 75382
rect 197353 74218 197419 74221
rect 197353 74216 200032 74218
rect 197353 74160 197358 74216
rect 197414 74160 200032 74216
rect 197353 74158 200032 74160
rect 197353 74155 197419 74158
rect 197353 72994 197419 72997
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 197353 72992 200032 72994
rect 197353 72936 197358 72992
rect 197414 72936 200032 72992
rect 197353 72934 200032 72936
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 197353 72931 197419 72934
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 559189 71906 559255 71909
rect 556876 71904 559255 71906
rect 556876 71848 559194 71904
rect 559250 71848 559255 71904
rect 556876 71846 559255 71848
rect 559189 71843 559255 71846
rect -960 71634 480 71724
rect 3693 71634 3759 71637
rect -960 71632 3759 71634
rect -960 71576 3698 71632
rect 3754 71576 3759 71632
rect -960 71574 3759 71576
rect -960 71484 480 71574
rect 3693 71571 3759 71574
rect 198273 71090 198339 71093
rect 200070 71090 200130 71600
rect 198273 71088 200130 71090
rect 198273 71032 198278 71088
rect 198334 71032 200130 71088
rect 198273 71030 200130 71032
rect 198273 71027 198339 71030
rect 197353 70410 197419 70413
rect 197353 70408 200032 70410
rect 197353 70352 197358 70408
rect 197414 70352 200032 70408
rect 197353 70350 200032 70352
rect 197353 70347 197419 70350
rect 198365 69186 198431 69189
rect 198365 69184 200032 69186
rect 198365 69128 198370 69184
rect 198426 69128 200032 69184
rect 198365 69126 200032 69128
rect 198365 69123 198431 69126
rect 198457 67962 198523 67965
rect 198457 67960 200032 67962
rect 198457 67904 198462 67960
rect 198518 67904 200032 67960
rect 198457 67902 200032 67904
rect 198457 67899 198523 67902
rect 168833 67010 168899 67013
rect 167134 67008 168899 67010
rect 167134 66952 168838 67008
rect 168894 66952 168899 67008
rect 167134 66950 168899 66952
rect 167134 66924 167194 66950
rect 168833 66947 168899 66950
rect 166612 66864 167194 66924
rect 198549 66738 198615 66741
rect 198549 66736 200032 66738
rect 198549 66680 198554 66736
rect 198610 66680 200032 66736
rect 198549 66678 200032 66680
rect 198549 66675 198615 66678
rect 168833 66058 168899 66061
rect 167134 66056 168899 66058
rect 167134 66000 168838 66056
rect 168894 66000 168899 66056
rect 167134 65998 168899 66000
rect 167134 65972 167194 65998
rect 168833 65995 168899 65998
rect 166612 65912 167194 65972
rect 198641 65514 198707 65517
rect 198641 65512 200032 65514
rect 198641 65456 198646 65512
rect 198702 65456 200032 65512
rect 198641 65454 200032 65456
rect 198641 65451 198707 65454
rect 168833 63882 168899 63885
rect 167134 63880 168899 63882
rect 167134 63824 168838 63880
rect 168894 63824 168899 63880
rect 167134 63822 168899 63824
rect 167134 63796 167194 63822
rect 168833 63819 168899 63822
rect 197353 63882 197419 63885
rect 200070 63882 200130 64256
rect 560201 64018 560267 64021
rect 556876 64016 560267 64018
rect 556876 63960 560206 64016
rect 560262 63960 560267 64016
rect 556876 63958 560267 63960
rect 560201 63955 560267 63958
rect 197353 63880 200130 63882
rect 197353 63824 197358 63880
rect 197414 63824 200130 63880
rect 197353 63822 200130 63824
rect 197353 63819 197419 63822
rect 166612 63736 167194 63796
rect 197905 63066 197971 63069
rect 197905 63064 200032 63066
rect 197905 63008 197910 63064
rect 197966 63008 200032 63064
rect 197905 63006 200032 63008
rect 197905 63003 197971 63006
rect 169385 62930 169451 62933
rect 167134 62928 169451 62930
rect 167134 62872 169390 62928
rect 169446 62872 169451 62928
rect 167134 62870 169451 62872
rect 167134 62844 167194 62870
rect 169385 62867 169451 62870
rect 166612 62784 167194 62844
rect 197353 61842 197419 61845
rect 197353 61840 200032 61842
rect 197353 61784 197358 61840
rect 197414 61784 200032 61840
rect 197353 61782 200032 61784
rect 197353 61779 197419 61782
rect 168925 61162 168991 61165
rect 167134 61160 168991 61162
rect 167134 61104 168930 61160
rect 168986 61104 168991 61160
rect 167134 61102 168991 61104
rect 167134 61076 167194 61102
rect 168925 61099 168991 61102
rect 166612 61016 167194 61076
rect 197537 60618 197603 60621
rect 197537 60616 200100 60618
rect 197537 60560 197542 60616
rect 197598 60560 200100 60616
rect 197537 60558 200100 60560
rect 197537 60555 197603 60558
rect 168833 60074 168899 60077
rect 167134 60072 168899 60074
rect 167134 60016 168838 60072
rect 168894 60016 168899 60072
rect 167134 60014 168899 60016
rect 167134 59988 167194 60014
rect 168833 60011 168899 60014
rect 166612 59928 167194 59988
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 168833 58306 168899 58309
rect 167134 58304 168899 58306
rect 167134 58248 168838 58304
rect 168894 58248 168899 58304
rect 167134 58246 168899 58248
rect 167134 58220 167194 58246
rect 168833 58243 168899 58246
rect 166612 58160 167194 58220
rect 27429 49466 27495 49469
rect 27429 49464 29378 49466
rect 27429 49408 27434 49464
rect 27490 49408 29378 49464
rect 27429 49406 29378 49408
rect 27429 49403 27495 49406
rect 29318 49380 29378 49406
rect 29318 49320 30032 49380
rect 27337 47834 27403 47837
rect 27337 47832 29378 47834
rect 27337 47776 27342 47832
rect 27398 47776 29378 47832
rect 27337 47774 29378 47776
rect 27337 47771 27403 47774
rect 29318 47748 29378 47774
rect 29318 47688 30032 47748
rect 27245 46474 27311 46477
rect 27245 46472 29378 46474
rect 27245 46416 27250 46472
rect 27306 46416 29378 46472
rect 27245 46414 29378 46416
rect 27245 46411 27311 46414
rect 29318 46388 29378 46414
rect 29318 46328 30032 46388
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3601 45522 3667 45525
rect -960 45520 3667 45522
rect -960 45464 3606 45520
rect 3662 45464 3667 45520
rect -960 45462 3667 45464
rect -960 45372 480 45462
rect 3601 45459 3667 45462
rect 27061 44978 27127 44981
rect 27061 44976 29378 44978
rect 27061 44920 27066 44976
rect 27122 44920 29378 44976
rect 27061 44918 29378 44920
rect 27061 44915 27127 44918
rect 29318 44892 29378 44918
rect 29318 44832 30032 44892
rect 27153 43754 27219 43757
rect 27153 43752 29378 43754
rect 27153 43696 27158 43752
rect 27214 43696 29378 43752
rect 27153 43694 29378 43696
rect 27153 43691 27219 43694
rect 29318 43668 29378 43694
rect 29318 43608 30032 43668
rect 166612 39946 167194 39996
rect 168373 39946 168439 39949
rect 166612 39944 168439 39946
rect 166612 39936 168378 39944
rect 167134 39888 168378 39936
rect 168434 39888 168439 39944
rect 167134 39886 168439 39888
rect 168373 39883 168439 39886
rect 168557 38450 168623 38453
rect 167134 38448 168623 38450
rect 167134 38392 168562 38448
rect 168618 38392 168623 38448
rect 167134 38390 168623 38392
rect 167134 38364 167194 38390
rect 168557 38387 168623 38390
rect 166612 38304 167194 38364
rect 168465 38178 168531 38181
rect 167134 38176 168531 38178
rect 167134 38120 168470 38176
rect 168526 38120 168531 38176
rect 167134 38118 168531 38120
rect 167134 38092 167194 38118
rect 168465 38115 168531 38118
rect 166612 38032 167194 38092
rect 580349 33146 580415 33149
rect 583520 33146 584960 33236
rect 580349 33144 584960 33146
rect 580349 33088 580354 33144
rect 580410 33088 584960 33144
rect 580349 33086 584960 33088
rect 580349 33083 580415 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 125472 29820 125478 29884
rect 125542 29882 125548 29884
rect 128353 29882 128419 29885
rect 125542 29880 128419 29882
rect 125542 29824 128358 29880
rect 128414 29824 128419 29880
rect 125542 29822 128419 29824
rect 125542 29820 125548 29822
rect 128353 29819 128419 29822
rect 75545 29612 75611 29613
rect 88057 29612 88123 29613
rect 90725 29612 90791 29613
rect 75545 29608 75566 29612
rect 75630 29610 75636 29612
rect 75545 29552 75550 29608
rect 75545 29548 75566 29552
rect 75630 29550 75702 29610
rect 88057 29608 88078 29612
rect 88142 29610 88148 29612
rect 90656 29610 90662 29612
rect 88057 29552 88062 29608
rect 75630 29548 75636 29550
rect 88057 29548 88078 29552
rect 88142 29550 88214 29610
rect 90634 29550 90662 29610
rect 88142 29548 88148 29550
rect 90656 29548 90662 29550
rect 90726 29608 90791 29612
rect 90726 29552 90730 29608
rect 90786 29552 90791 29608
rect 90726 29548 90791 29552
rect 75545 29547 75611 29548
rect 88057 29547 88123 29548
rect 90725 29547 90791 29548
rect 122741 29610 122807 29613
rect 130561 29612 130627 29613
rect 123704 29610 123710 29612
rect 122741 29608 123710 29610
rect 122741 29552 122746 29608
rect 122802 29552 123710 29608
rect 122741 29550 123710 29552
rect 122741 29547 122807 29550
rect 123704 29548 123710 29550
rect 123774 29548 123780 29612
rect 130504 29610 130510 29612
rect 130470 29550 130510 29610
rect 130574 29608 130627 29612
rect 130622 29552 130627 29608
rect 130504 29548 130510 29550
rect 130574 29548 130627 29552
rect 130561 29547 130627 29548
rect 138933 29612 138999 29613
rect 138933 29608 138942 29612
rect 139006 29610 139012 29612
rect 138933 29552 138938 29608
rect 138933 29548 138942 29552
rect 139006 29550 139090 29610
rect 139006 29548 139012 29550
rect 138933 29547 138999 29548
rect 60641 28932 60707 28933
rect 68185 28932 68251 28933
rect 78121 28932 78187 28933
rect 80697 28932 80763 28933
rect 83089 28932 83155 28933
rect 103145 28932 103211 28933
rect 128537 28932 128603 28933
rect 134241 28932 134307 28933
rect 135897 28932 135963 28933
rect 138289 28932 138355 28933
rect 60590 28930 60596 28932
rect 60550 28870 60596 28930
rect 60660 28928 60707 28932
rect 68134 28930 68140 28932
rect 60702 28872 60707 28928
rect 60590 28868 60596 28870
rect 60660 28868 60707 28872
rect 68094 28870 68140 28930
rect 68204 28928 68251 28932
rect 78070 28930 78076 28932
rect 68246 28872 68251 28928
rect 68134 28868 68140 28870
rect 68204 28868 68251 28872
rect 78030 28870 78076 28930
rect 78140 28928 78187 28932
rect 80646 28930 80652 28932
rect 78182 28872 78187 28928
rect 78070 28868 78076 28870
rect 78140 28868 78187 28872
rect 80606 28870 80652 28930
rect 80716 28928 80763 28932
rect 83038 28930 83044 28932
rect 80758 28872 80763 28928
rect 80646 28868 80652 28870
rect 80716 28868 80763 28872
rect 82998 28870 83044 28930
rect 83108 28928 83155 28932
rect 103094 28930 103100 28932
rect 83150 28872 83155 28928
rect 83038 28868 83044 28870
rect 83108 28868 83155 28872
rect 103054 28870 103100 28930
rect 103164 28928 103211 28932
rect 128486 28930 128492 28932
rect 103206 28872 103211 28928
rect 103094 28868 103100 28870
rect 103164 28868 103211 28872
rect 128446 28870 128492 28930
rect 128556 28928 128603 28932
rect 134190 28930 134196 28932
rect 128598 28872 128603 28928
rect 128486 28868 128492 28870
rect 128556 28868 128603 28872
rect 134150 28870 134196 28930
rect 134260 28928 134307 28932
rect 135846 28930 135852 28932
rect 134302 28872 134307 28928
rect 134190 28868 134196 28870
rect 134260 28868 134307 28872
rect 135806 28870 135852 28930
rect 135916 28928 135963 28932
rect 138238 28930 138244 28932
rect 135958 28872 135963 28928
rect 135846 28868 135852 28870
rect 135916 28868 135963 28872
rect 138198 28870 138244 28930
rect 138308 28928 138355 28932
rect 188337 28930 188403 28933
rect 138350 28872 138355 28928
rect 138238 28868 138244 28870
rect 138308 28868 138355 28872
rect 60641 28867 60707 28868
rect 68185 28867 68251 28868
rect 78121 28867 78187 28868
rect 80697 28867 80763 28868
rect 83089 28867 83155 28868
rect 103145 28867 103211 28868
rect 128537 28867 128603 28868
rect 134241 28867 134307 28868
rect 135897 28867 135963 28868
rect 138289 28867 138355 28868
rect 142110 28928 188403 28930
rect 142110 28872 188342 28928
rect 188398 28872 188403 28928
rect 142110 28870 188403 28872
rect 133086 28732 133092 28796
rect 133156 28794 133162 28796
rect 142110 28794 142170 28870
rect 188337 28867 188403 28870
rect 170581 28794 170647 28797
rect 133156 28734 142170 28794
rect 151770 28792 170647 28794
rect 151770 28736 170586 28792
rect 170642 28736 170647 28792
rect 151770 28734 170647 28736
rect 133156 28732 133162 28734
rect 135294 28596 135300 28660
rect 135364 28658 135370 28660
rect 151770 28658 151830 28734
rect 170581 28731 170647 28734
rect 135364 28598 151830 28658
rect 135364 28596 135370 28598
rect 149053 28386 149119 28389
rect 178677 28386 178743 28389
rect 149053 28384 178743 28386
rect 149053 28328 149058 28384
rect 149114 28328 178682 28384
rect 178738 28328 178743 28384
rect 149053 28326 178743 28328
rect 149053 28323 149119 28326
rect 178677 28323 178743 28326
rect 63217 28252 63283 28253
rect 112161 28252 112227 28253
rect 115657 28252 115723 28253
rect 129641 28252 129707 28253
rect 132033 28252 132099 28253
rect 143441 28252 143507 28253
rect 63166 28250 63172 28252
rect 63126 28190 63172 28250
rect 63236 28248 63283 28252
rect 112110 28250 112116 28252
rect 63278 28192 63283 28248
rect 63166 28188 63172 28190
rect 63236 28188 63283 28192
rect 112070 28190 112116 28250
rect 112180 28248 112227 28252
rect 115606 28250 115612 28252
rect 112222 28192 112227 28248
rect 112110 28188 112116 28190
rect 112180 28188 112227 28192
rect 115566 28190 115612 28250
rect 115676 28248 115723 28252
rect 129590 28250 129596 28252
rect 115718 28192 115723 28248
rect 115606 28188 115612 28190
rect 115676 28188 115723 28192
rect 129550 28190 129596 28250
rect 129660 28248 129707 28252
rect 131982 28250 131988 28252
rect 129702 28192 129707 28248
rect 129590 28188 129596 28190
rect 129660 28188 129707 28192
rect 131942 28190 131988 28250
rect 132052 28248 132099 28252
rect 143390 28250 143396 28252
rect 132094 28192 132099 28248
rect 131982 28188 131988 28190
rect 132052 28188 132099 28192
rect 143350 28190 143396 28250
rect 143460 28248 143507 28252
rect 181529 28250 181595 28253
rect 143502 28192 143507 28248
rect 143390 28188 143396 28190
rect 143460 28188 143507 28192
rect 63217 28187 63283 28188
rect 112161 28187 112227 28188
rect 115657 28187 115723 28188
rect 129641 28187 129707 28188
rect 132033 28187 132099 28188
rect 143441 28187 143507 28188
rect 151770 28248 181595 28250
rect 151770 28192 181534 28248
rect 181590 28192 181595 28248
rect 151770 28190 181595 28192
rect 143349 28114 143415 28117
rect 151770 28114 151830 28190
rect 181529 28187 181595 28190
rect 143349 28112 151830 28114
rect 143349 28056 143354 28112
rect 143410 28056 151830 28112
rect 143349 28054 151830 28056
rect 143349 28051 143415 28054
rect 122741 27706 122807 27709
rect 122741 27704 122850 27706
rect 122741 27648 122746 27704
rect 122802 27648 122850 27704
rect 122741 27643 122850 27648
rect 42793 27572 42859 27573
rect 42742 27570 42748 27572
rect 42702 27510 42748 27570
rect 42812 27568 42859 27572
rect 42854 27512 42859 27568
rect 42742 27508 42748 27510
rect 42812 27508 42859 27512
rect 42793 27507 42859 27508
rect 43621 27572 43687 27573
rect 64873 27572 64939 27573
rect 43621 27568 43668 27572
rect 43732 27570 43738 27572
rect 43621 27512 43626 27568
rect 43621 27508 43668 27512
rect 43732 27510 43778 27570
rect 43732 27508 43738 27510
rect 64822 27508 64828 27572
rect 64892 27570 64939 27572
rect 64892 27568 64984 27570
rect 64934 27512 64984 27568
rect 64892 27510 64984 27512
rect 64892 27508 64939 27510
rect 70710 27508 70716 27572
rect 70780 27570 70786 27572
rect 71589 27570 71655 27573
rect 70780 27568 71655 27570
rect 70780 27512 71594 27568
rect 71650 27512 71655 27568
rect 70780 27510 71655 27512
rect 70780 27508 70786 27510
rect 43621 27507 43687 27508
rect 64873 27507 64939 27508
rect 71589 27507 71655 27510
rect 73654 27508 73660 27572
rect 73724 27570 73730 27572
rect 73981 27570 74047 27573
rect 73724 27568 74047 27570
rect 73724 27512 73986 27568
rect 74042 27512 74047 27568
rect 73724 27510 74047 27512
rect 73724 27508 73730 27510
rect 73981 27507 74047 27510
rect 86350 27508 86356 27572
rect 86420 27570 86426 27572
rect 86585 27570 86651 27573
rect 86420 27568 86651 27570
rect 86420 27512 86590 27568
rect 86646 27512 86651 27568
rect 86420 27510 86651 27512
rect 86420 27508 86426 27510
rect 86585 27507 86651 27510
rect 92749 27572 92815 27573
rect 95233 27572 95299 27573
rect 92749 27568 92796 27572
rect 92860 27570 92866 27572
rect 95182 27570 95188 27572
rect 92749 27512 92754 27568
rect 92749 27508 92796 27512
rect 92860 27510 92906 27570
rect 95142 27510 95188 27570
rect 95252 27568 95299 27572
rect 95294 27512 95299 27568
rect 92860 27508 92866 27510
rect 95182 27508 95188 27510
rect 95252 27508 95299 27512
rect 92749 27507 92815 27508
rect 95233 27507 95299 27508
rect 98269 27572 98335 27573
rect 98269 27568 98316 27572
rect 98380 27570 98386 27572
rect 100201 27570 100267 27573
rect 100518 27570 100524 27572
rect 98269 27512 98274 27568
rect 98269 27508 98316 27512
rect 98380 27510 98426 27570
rect 100201 27568 100524 27570
rect 100201 27512 100206 27568
rect 100262 27512 100524 27568
rect 100201 27510 100524 27512
rect 98380 27508 98386 27510
rect 98269 27507 98335 27508
rect 100201 27507 100267 27510
rect 100518 27508 100524 27510
rect 100588 27508 100594 27572
rect 105302 27508 105308 27572
rect 105372 27570 105378 27572
rect 105537 27570 105603 27573
rect 105372 27568 105603 27570
rect 105372 27512 105542 27568
rect 105598 27512 105603 27568
rect 105372 27510 105603 27512
rect 105372 27508 105378 27510
rect 105537 27507 105603 27510
rect 106273 27570 106339 27573
rect 108021 27572 108087 27573
rect 107326 27570 107332 27572
rect 106273 27568 107332 27570
rect 106273 27512 106278 27568
rect 106334 27512 107332 27568
rect 106273 27510 107332 27512
rect 106273 27507 106339 27510
rect 107326 27508 107332 27510
rect 107396 27508 107402 27572
rect 108021 27568 108068 27572
rect 108132 27570 108138 27572
rect 108021 27512 108026 27568
rect 108021 27508 108068 27512
rect 108132 27510 108178 27570
rect 108132 27508 108138 27510
rect 108430 27508 108436 27572
rect 108500 27570 108506 27572
rect 108757 27570 108823 27573
rect 108500 27568 108823 27570
rect 108500 27512 108762 27568
rect 108818 27512 108823 27568
rect 108500 27510 108823 27512
rect 108500 27508 108506 27510
rect 108021 27507 108087 27508
rect 108757 27507 108823 27510
rect 110086 27508 110092 27572
rect 110156 27570 110162 27572
rect 110321 27570 110387 27573
rect 110156 27568 110387 27570
rect 110156 27512 110326 27568
rect 110382 27512 110387 27568
rect 110156 27510 110387 27512
rect 110156 27508 110162 27510
rect 110321 27507 110387 27510
rect 110822 27508 110828 27572
rect 110892 27570 110898 27572
rect 110965 27570 111031 27573
rect 110892 27568 111031 27570
rect 110892 27512 110970 27568
rect 111026 27512 111031 27568
rect 110892 27510 111031 27512
rect 110892 27508 110898 27510
rect 110965 27507 111031 27510
rect 112662 27508 112668 27572
rect 112732 27570 112738 27572
rect 112897 27570 112963 27573
rect 112732 27568 112963 27570
rect 112732 27512 112902 27568
rect 112958 27512 112963 27568
rect 112732 27510 112963 27512
rect 112732 27508 112738 27510
rect 112897 27507 112963 27510
rect 116710 27508 116716 27572
rect 116780 27570 116786 27572
rect 117129 27570 117195 27573
rect 116780 27568 117195 27570
rect 116780 27512 117134 27568
rect 117190 27512 117195 27568
rect 116780 27510 117195 27512
rect 116780 27508 116786 27510
rect 117129 27507 117195 27510
rect 117814 27508 117820 27572
rect 117884 27570 117890 27572
rect 118233 27570 118299 27573
rect 118417 27572 118483 27573
rect 117884 27568 118299 27570
rect 117884 27512 118238 27568
rect 118294 27512 118299 27568
rect 117884 27510 118299 27512
rect 117884 27508 117890 27510
rect 118233 27507 118299 27510
rect 118366 27508 118372 27572
rect 118436 27570 118483 27572
rect 118436 27568 118528 27570
rect 118478 27512 118528 27568
rect 118436 27510 118528 27512
rect 118436 27508 118483 27510
rect 120206 27508 120212 27572
rect 120276 27570 120282 27572
rect 120809 27570 120875 27573
rect 120276 27568 120875 27570
rect 120276 27512 120814 27568
rect 120870 27512 120875 27568
rect 120276 27510 120875 27512
rect 122790 27570 122850 27643
rect 124121 27570 124187 27573
rect 126329 27572 126395 27573
rect 128169 27572 128235 27573
rect 132769 27572 132835 27573
rect 126278 27570 126284 27572
rect 122790 27568 124187 27570
rect 122790 27512 124126 27568
rect 124182 27512 124187 27568
rect 122790 27510 124187 27512
rect 126238 27510 126284 27570
rect 126348 27568 126395 27572
rect 128118 27570 128124 27572
rect 126390 27512 126395 27568
rect 120276 27508 120282 27510
rect 118417 27507 118483 27508
rect 120809 27507 120875 27510
rect 124121 27507 124187 27510
rect 126278 27508 126284 27510
rect 126348 27508 126395 27512
rect 128078 27510 128124 27570
rect 128188 27568 128235 27572
rect 132718 27570 132724 27572
rect 128230 27512 128235 27568
rect 128118 27508 128124 27510
rect 128188 27508 128235 27512
rect 132678 27510 132724 27570
rect 132788 27568 132835 27572
rect 132830 27512 132835 27568
rect 132718 27508 132724 27510
rect 132788 27508 132835 27512
rect 126329 27507 126395 27508
rect 128169 27507 128235 27508
rect 132769 27507 132835 27508
rect 135345 27570 135411 27573
rect 136398 27570 136404 27572
rect 135345 27568 136404 27570
rect 135345 27512 135350 27568
rect 135406 27512 136404 27568
rect 135345 27510 136404 27512
rect 135345 27507 135411 27510
rect 136398 27508 136404 27510
rect 136468 27508 136474 27572
rect 137185 27570 137251 27573
rect 140129 27572 140195 27573
rect 141233 27572 141299 27573
rect 137870 27570 137876 27572
rect 137185 27568 137876 27570
rect 137185 27512 137190 27568
rect 137246 27512 137876 27568
rect 137185 27510 137876 27512
rect 137185 27507 137251 27510
rect 137870 27508 137876 27510
rect 137940 27508 137946 27572
rect 140078 27570 140084 27572
rect 140038 27510 140084 27570
rect 140148 27568 140195 27572
rect 141182 27570 141188 27572
rect 140190 27512 140195 27568
rect 140078 27508 140084 27510
rect 140148 27508 140195 27512
rect 141142 27510 141188 27570
rect 141252 27568 141299 27572
rect 141294 27512 141299 27568
rect 141182 27508 141188 27510
rect 141252 27508 141299 27512
rect 147070 27508 147076 27572
rect 147140 27570 147146 27572
rect 147673 27570 147739 27573
rect 150065 27572 150131 27573
rect 150617 27572 150683 27573
rect 148358 27570 148364 27572
rect 147140 27568 148364 27570
rect 147140 27512 147678 27568
rect 147734 27512 148364 27568
rect 147140 27510 148364 27512
rect 147140 27508 147146 27510
rect 140129 27507 140195 27508
rect 141233 27507 141299 27508
rect 147673 27507 147739 27510
rect 148358 27508 148364 27510
rect 148428 27508 148434 27572
rect 150014 27570 150020 27572
rect 149974 27510 150020 27570
rect 150084 27568 150131 27572
rect 150566 27570 150572 27572
rect 150126 27512 150131 27568
rect 150014 27508 150020 27510
rect 150084 27508 150131 27512
rect 150526 27510 150572 27570
rect 150636 27568 150683 27572
rect 150678 27512 150683 27568
rect 150566 27508 150572 27510
rect 150636 27508 150683 27512
rect 150065 27507 150131 27508
rect 150617 27507 150683 27508
rect 110454 27372 110460 27436
rect 110524 27434 110530 27436
rect 111517 27434 111583 27437
rect 110524 27432 111583 27434
rect 110524 27376 111522 27432
rect 111578 27376 111583 27432
rect 110524 27374 111583 27376
rect 110524 27372 110530 27374
rect 111517 27371 111583 27374
rect 120073 27434 120139 27437
rect 121310 27434 121316 27436
rect 120073 27432 121316 27434
rect 120073 27376 120078 27432
rect 120134 27376 121316 27432
rect 120073 27374 121316 27376
rect 120073 27371 120139 27374
rect 121310 27372 121316 27374
rect 121380 27372 121386 27436
rect 177297 27434 177363 27437
rect 121502 27432 177363 27434
rect 121502 27376 177302 27432
rect 177358 27376 177363 27432
rect 121502 27374 177363 27376
rect 120625 27300 120691 27301
rect 120574 27298 120580 27300
rect 120534 27238 120580 27298
rect 120644 27296 120691 27300
rect 120686 27240 120691 27296
rect 120574 27236 120580 27238
rect 120644 27236 120691 27240
rect 120625 27235 120691 27236
rect 113766 27100 113772 27164
rect 113836 27162 113842 27164
rect 121502 27162 121562 27374
rect 177297 27371 177363 27374
rect 170489 27298 170555 27301
rect 113836 27102 121562 27162
rect 122790 27296 170555 27298
rect 122790 27240 170494 27296
rect 170550 27240 170555 27296
rect 122790 27238 170555 27240
rect 113836 27100 113842 27102
rect 114318 26964 114324 27028
rect 114388 27026 114394 27028
rect 122790 27026 122850 27238
rect 170489 27235 170555 27238
rect 123753 27164 123819 27165
rect 123702 27162 123708 27164
rect 123662 27102 123708 27162
rect 123772 27160 123819 27164
rect 123814 27104 123819 27160
rect 123702 27100 123708 27102
rect 123772 27100 123819 27104
rect 127198 27100 127204 27164
rect 127268 27162 127274 27164
rect 178769 27162 178835 27165
rect 127268 27160 178835 27162
rect 127268 27104 178774 27160
rect 178830 27104 178835 27160
rect 127268 27102 178835 27104
rect 127268 27100 127274 27102
rect 123753 27099 123819 27100
rect 178769 27099 178835 27102
rect 114388 26966 122850 27026
rect 114388 26964 114394 26966
rect 124806 26964 124812 27028
rect 124876 27026 124882 27028
rect 174629 27026 174695 27029
rect 124876 27024 174695 27026
rect 124876 26968 174634 27024
rect 174690 26968 174695 27024
rect 124876 26966 174695 26968
rect 124876 26964 124882 26966
rect 174629 26963 174695 26966
rect 122598 26828 122604 26892
rect 122668 26890 122674 26892
rect 170673 26890 170739 26893
rect 122668 26888 170739 26890
rect 122668 26832 170678 26888
rect 170734 26832 170739 26888
rect 122668 26830 170739 26832
rect 122668 26828 122674 26830
rect 170673 26827 170739 26830
rect 130694 26692 130700 26756
rect 130764 26754 130770 26756
rect 177481 26754 177547 26757
rect 130764 26752 177547 26754
rect 130764 26696 177486 26752
rect 177542 26696 177547 26752
rect 130764 26694 177547 26696
rect 130764 26692 130770 26694
rect 177481 26691 177547 26694
rect 142654 26556 142660 26620
rect 142724 26618 142730 26620
rect 143441 26618 143507 26621
rect 142724 26616 143507 26618
rect 142724 26560 143446 26616
rect 143502 26560 143507 26616
rect 142724 26558 143507 26560
rect 142724 26556 142730 26558
rect 143441 26555 143507 26558
rect 115238 26346 115244 26348
rect 114510 26286 115244 26346
rect 114510 26210 114570 26286
rect 115238 26284 115244 26286
rect 115308 26284 115314 26348
rect 118918 26284 118924 26348
rect 118988 26346 118994 26348
rect 196801 26346 196867 26349
rect 118988 26344 196867 26346
rect 118988 26288 196806 26344
rect 196862 26288 196867 26344
rect 118988 26286 196867 26288
rect 118988 26284 118994 26286
rect 196801 26283 196867 26286
rect 170397 26210 170463 26213
rect 114510 26208 170463 26210
rect 114510 26152 170402 26208
rect 170458 26152 170463 26208
rect 114510 26150 170463 26152
rect 170397 26147 170463 26150
rect 137185 24850 137251 24853
rect 193949 24850 194015 24853
rect 137185 24848 194015 24850
rect 137185 24792 137190 24848
rect 137246 24792 193954 24848
rect 194010 24792 194015 24848
rect 137185 24790 194015 24792
rect 137185 24787 137251 24790
rect 193949 24787 194015 24790
rect 579613 19818 579679 19821
rect 583520 19818 584960 19908
rect 579613 19816 584960 19818
rect 579613 19760 579618 19816
rect 579674 19760 584960 19816
rect 579613 19758 584960 19760
rect 579613 19755 579679 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect -960 6430 674 6490
rect 583520 6476 584960 6566
rect -960 6354 480 6430
rect 614 6354 674 6430
rect -960 6340 674 6354
rect 246 6294 674 6340
rect 246 5810 306 6294
rect 246 5750 6930 5810
rect 6870 5674 6930 5750
rect 174486 5674 174492 5676
rect 6870 5614 174492 5674
rect 174486 5612 174492 5614
rect 174556 5612 174562 5676
<< via3 >>
rect 196572 700572 196636 700636
rect 174676 700436 174740 700500
rect 174492 700300 174556 700364
rect 35756 674868 35820 674932
rect 46796 674868 46860 674932
rect 48084 674868 48148 674932
rect 246252 659696 246316 659700
rect 246252 659640 246302 659696
rect 246302 659640 246316 659696
rect 246252 659636 246316 659640
rect 256556 659636 256620 659700
rect 340092 659696 340156 659700
rect 340092 659640 340142 659696
rect 340142 659640 340156 659696
rect 340092 659636 340156 659640
rect 488948 659696 489012 659700
rect 488948 659640 488962 659696
rect 488962 659640 489012 659696
rect 488948 659636 489012 659640
rect 499988 659636 500052 659700
rect 338252 612172 338316 612236
rect 338068 610948 338132 611012
rect 144790 589732 144854 589796
rect 146014 589732 146078 589796
rect 43116 588100 43180 588164
rect 63172 588100 63236 588164
rect 73108 588100 73172 588164
rect 83044 588100 83108 588164
rect 85620 588100 85684 588164
rect 95556 588100 95620 588164
rect 103100 588100 103164 588164
rect 109540 588100 109604 588164
rect 112116 588100 112180 588164
rect 113036 588100 113100 588164
rect 115612 588100 115676 588164
rect 122972 588100 123036 588164
rect 129596 588100 129660 588164
rect 133092 588100 133156 588164
rect 143396 588100 143460 588164
rect 149468 588100 149532 588164
rect 43668 587828 43732 587892
rect 60596 587888 60660 587892
rect 60596 587832 60646 587888
rect 60646 587832 60660 587888
rect 60596 587828 60660 587832
rect 68140 587828 68204 587892
rect 88196 587888 88260 587892
rect 88196 587832 88246 587888
rect 88246 587832 88260 587888
rect 88196 587828 88260 587832
rect 98316 587828 98380 587892
rect 100524 587888 100588 587892
rect 100524 587832 100574 587888
rect 100574 587832 100588 587888
rect 100524 587828 100588 587832
rect 105308 587828 105372 587892
rect 107332 587828 107396 587892
rect 108436 587828 108500 587892
rect 110460 587888 110524 587892
rect 110460 587832 110510 587888
rect 110510 587832 110524 587888
rect 110460 587828 110524 587832
rect 110828 587828 110892 587892
rect 114324 587828 114388 587892
rect 115244 587828 115308 587892
rect 113772 587692 113836 587756
rect 116716 587828 116780 587892
rect 118924 587828 118988 587892
rect 120212 587888 120276 587892
rect 120212 587832 120262 587888
rect 120262 587832 120276 587888
rect 120212 587828 120276 587832
rect 121316 587828 121380 587892
rect 122604 587888 122668 587892
rect 122604 587832 122654 587888
rect 122654 587832 122668 587888
rect 122604 587828 122668 587832
rect 124812 587828 124876 587892
rect 126284 587828 126348 587892
rect 128492 587828 128556 587892
rect 130700 587828 130764 587892
rect 131620 587828 131684 587892
rect 132724 587828 132788 587892
rect 136220 587828 136284 587892
rect 137876 587888 137940 587892
rect 137876 587832 137926 587888
rect 137926 587832 137940 587888
rect 137876 587828 137940 587832
rect 138244 587828 138308 587892
rect 140084 587888 140148 587892
rect 140084 587832 140134 587888
rect 140134 587832 140148 587888
rect 140084 587828 140148 587832
rect 142660 587888 142724 587892
rect 142660 587832 142710 587888
rect 142710 587832 142724 587888
rect 142660 587828 142724 587832
rect 147076 587828 147140 587892
rect 148364 587828 148428 587892
rect 150572 587828 150636 587892
rect 120580 587692 120644 587756
rect 130516 587692 130580 587756
rect 134196 587692 134260 587756
rect 166948 587692 167012 587756
rect 135300 587556 135364 587620
rect 170076 587556 170140 587620
rect 127204 587420 127268 587484
rect 123708 587284 123772 587348
rect 170260 587284 170324 587348
rect 117820 587012 117884 587076
rect 136588 587072 136652 587076
rect 136588 587016 136602 587072
rect 136602 587016 136652 587072
rect 136588 587012 136652 587016
rect 138980 587072 139044 587076
rect 138980 587016 139030 587072
rect 139030 587016 139044 587072
rect 138980 587012 139044 587016
rect 64828 586528 64892 586532
rect 64828 586472 64878 586528
rect 64878 586472 64892 586528
rect 64828 586468 64892 586472
rect 70716 586604 70780 586668
rect 75316 586604 75380 586668
rect 78076 586604 78140 586668
rect 80652 586604 80716 586668
rect 90588 586604 90652 586668
rect 92796 586604 92860 586668
rect 108068 586604 108132 586668
rect 118188 586604 118252 586668
rect 125364 586604 125428 586668
rect 128124 586604 128188 586668
rect 141004 586604 141068 586668
rect 168420 584836 168484 584900
rect 167132 584700 167196 584764
rect 172652 584428 172716 584492
rect 168604 581708 168668 581772
rect 167684 581572 167748 581636
rect 252508 577764 252572 577828
rect 252926 577764 252990 577828
rect 284892 577764 284956 577828
rect 285294 577764 285358 577828
rect 445156 577764 445220 577828
rect 445502 577764 445566 577828
rect 492694 577824 492758 577828
rect 492694 577768 492734 577824
rect 492734 577768 492758 577824
rect 492694 577764 492758 577768
rect 493102 577764 493166 577828
rect 492628 577628 492692 577692
rect 280108 577492 280172 577556
rect 281486 577492 281550 577556
rect 441844 577008 441908 577012
rect 441844 576952 441858 577008
rect 441858 576952 441908 577008
rect 441844 576948 441908 576952
rect 462820 577008 462884 577012
rect 462820 576952 462870 577008
rect 462870 576952 462884 577008
rect 462820 576948 462884 576952
rect 492996 576872 493060 576876
rect 492996 576816 493010 576872
rect 493010 576816 493060 576872
rect 492996 576812 493060 576816
rect 253060 576192 253124 576196
rect 253060 576136 253110 576192
rect 253110 576136 253124 576192
rect 253060 576132 253124 576136
rect 292436 576192 292500 576196
rect 292436 576136 292486 576192
rect 292486 576136 292500 576192
rect 292436 576132 292500 576136
rect 455460 576192 455524 576196
rect 455460 576136 455510 576192
rect 455510 576136 455524 576192
rect 455460 576132 455524 576136
rect 459324 576192 459388 576196
rect 459324 576136 459338 576192
rect 459338 576136 459388 576192
rect 459324 576132 459388 576136
rect 469260 576132 469324 576196
rect 341564 575996 341628 576060
rect 284156 575376 284220 575380
rect 284156 575320 284206 575376
rect 284206 575320 284220 575376
rect 284156 575316 284220 575320
rect 285260 575376 285324 575380
rect 285260 575320 285310 575376
rect 285310 575320 285324 575376
rect 285260 575316 285324 575320
rect 286548 575376 286612 575380
rect 286548 575320 286598 575376
rect 286598 575320 286612 575376
rect 286548 575316 286612 575320
rect 287652 575316 287716 575380
rect 297036 575316 297100 575380
rect 300532 575316 300596 575380
rect 301636 575316 301700 575380
rect 302740 575316 302804 575380
rect 304212 575316 304276 575380
rect 305132 575316 305196 575380
rect 306236 575376 306300 575380
rect 306236 575320 306286 575376
rect 306286 575320 306300 575376
rect 306236 575316 306300 575320
rect 307524 575376 307588 575380
rect 307524 575320 307574 575376
rect 307574 575320 307588 575376
rect 307524 575316 307588 575320
rect 320404 575376 320468 575380
rect 320404 575320 320454 575376
rect 320454 575320 320468 575376
rect 320404 575316 320468 575320
rect 330156 575376 330220 575380
rect 330156 575320 330206 575376
rect 330206 575320 330220 575376
rect 330156 575316 330220 575320
rect 336964 575316 337028 575380
rect 415348 575376 415412 575380
rect 415348 575320 415398 575376
rect 415398 575320 415412 575376
rect 415348 575316 415412 575320
rect 425284 575316 425348 575380
rect 284892 575180 284956 575244
rect 290228 575180 290292 575244
rect 293908 575240 293972 575244
rect 293908 575184 293958 575240
rect 293958 575184 293972 575240
rect 293908 575180 293972 575184
rect 314516 575180 314580 575244
rect 426756 575180 426820 575244
rect 438348 575180 438412 575244
rect 467604 575180 467668 575244
rect 280108 575104 280172 575108
rect 280108 575048 280158 575104
rect 280158 575048 280172 575104
rect 280108 575044 280172 575048
rect 291516 575044 291580 575108
rect 295196 575044 295260 575108
rect 312676 575044 312740 575108
rect 442764 575044 442828 575108
rect 448836 575044 448900 575108
rect 280292 574968 280356 574972
rect 280292 574912 280306 574968
rect 280306 574912 280356 574968
rect 280292 574908 280356 574912
rect 282684 574908 282748 574972
rect 288020 574908 288084 574972
rect 290044 574908 290108 574972
rect 310836 574908 310900 574972
rect 431356 574908 431420 574972
rect 284524 574772 284588 574836
rect 288940 574772 289004 574836
rect 290964 574832 291028 574836
rect 290964 574776 291014 574832
rect 291014 574776 291028 574832
rect 290964 574772 291028 574776
rect 292804 574772 292868 574836
rect 310100 574772 310164 574836
rect 432644 574772 432708 574836
rect 440004 574772 440068 574836
rect 445156 574772 445220 574836
rect 307892 574636 307956 574700
rect 308628 574636 308692 574700
rect 452516 574636 452580 574700
rect 288756 574500 288820 574564
rect 296300 574500 296364 574564
rect 298324 574500 298388 574564
rect 299060 574500 299124 574564
rect 300164 574500 300228 574564
rect 451412 574500 451476 574564
rect 456380 574500 456444 574564
rect 463924 574500 463988 574564
rect 253796 574424 253860 574428
rect 253796 574368 253810 574424
rect 253810 574368 253860 574424
rect 253796 574364 253860 574368
rect 274036 574364 274100 574428
rect 276612 574364 276676 574428
rect 293724 574424 293788 574428
rect 293724 574368 293774 574424
rect 293774 574368 293788 574424
rect 293724 574364 293788 574368
rect 294644 574424 294708 574428
rect 294644 574368 294694 574424
rect 294694 574368 294708 574424
rect 294644 574364 294708 574368
rect 433748 574364 433812 574428
rect 458220 574424 458284 574428
rect 458220 574368 458234 574424
rect 458234 574368 458284 574424
rect 458220 574364 458284 574368
rect 460796 574364 460860 574428
rect 465028 574424 465092 574428
rect 465028 574368 465078 574424
rect 465078 574368 465092 574424
rect 465028 574364 465092 574368
rect 492628 574424 492692 574428
rect 492628 574368 492678 574424
rect 492678 574368 492692 574424
rect 492628 574364 492692 574368
rect 252692 574228 252756 574292
rect 270356 574228 270420 574292
rect 275324 574228 275388 574292
rect 278820 574288 278884 574292
rect 278820 574232 278834 574288
rect 278834 574232 278884 574288
rect 278820 574228 278884 574232
rect 286732 574228 286796 574292
rect 298876 574228 298940 574292
rect 303844 574228 303908 574292
rect 313780 574228 313844 574292
rect 436324 574228 436388 574292
rect 440740 574228 440804 574292
rect 444052 574228 444116 574292
rect 445340 574228 445404 574292
rect 446628 574228 446692 574292
rect 447548 574228 447612 574292
rect 450308 574228 450372 574292
rect 452700 574288 452764 574292
rect 452700 574232 452750 574288
rect 452750 574232 452764 574288
rect 452700 574228 452764 574232
rect 454908 574228 454972 574292
rect 457116 574228 457180 574292
rect 461348 574228 461412 574292
rect 465212 574228 465276 574292
rect 471468 574228 471532 574292
rect 492628 574228 492692 574292
rect 252508 574092 252572 574156
rect 269068 574152 269132 574156
rect 269068 574096 269118 574152
rect 269118 574096 269132 574152
rect 269068 574092 269132 574096
rect 271460 574092 271524 574156
rect 272748 574092 272812 574156
rect 278084 574092 278148 574156
rect 278268 574092 278332 574156
rect 279004 574092 279068 574156
rect 280660 574092 280724 574156
rect 282500 574092 282564 574156
rect 283788 574092 283852 574156
rect 296484 574092 296548 574156
rect 298140 574152 298204 574156
rect 298140 574096 298154 574152
rect 298154 574096 298204 574152
rect 298140 574092 298204 574096
rect 301452 574092 301516 574156
rect 302556 574092 302620 574156
rect 305316 574092 305380 574156
rect 306604 574092 306668 574156
rect 318932 574092 318996 574156
rect 336780 574092 336844 574156
rect 434852 574092 434916 574156
rect 437244 574092 437308 574156
rect 437796 574092 437860 574156
rect 439084 574092 439148 574156
rect 440372 574092 440436 574156
rect 442580 574092 442644 574156
rect 443684 574092 443748 574156
rect 444420 574152 444484 574156
rect 444420 574096 444470 574152
rect 444470 574096 444484 574152
rect 444420 574092 444484 574096
rect 446812 574092 446876 574156
rect 447916 574092 447980 574156
rect 449020 574092 449084 574156
rect 450676 574092 450740 574156
rect 451596 574092 451660 574156
rect 453804 574092 453868 574156
rect 454356 574092 454420 574156
rect 456564 574092 456628 574156
rect 457852 574092 457916 574156
rect 458956 574092 459020 574156
rect 460612 574092 460676 574156
rect 461532 574092 461596 574156
rect 462636 574092 462700 574156
rect 464292 574092 464356 574156
rect 466500 574152 466564 574156
rect 466500 574096 466514 574152
rect 466514 574096 466564 574152
rect 466500 574092 466564 574096
rect 466868 574092 466932 574156
rect 467788 574152 467852 574156
rect 467788 574096 467838 574152
rect 467838 574096 467852 574152
rect 467788 574092 467852 574096
rect 470548 574152 470612 574156
rect 470548 574096 470598 574152
rect 470598 574096 470612 574152
rect 470548 574092 470612 574096
rect 472756 574092 472820 574156
rect 474228 574092 474292 574156
rect 475332 574092 475396 574156
rect 476804 574092 476868 574156
rect 35756 563136 35820 563140
rect 35756 563080 35770 563136
rect 35770 563080 35820 563136
rect 35756 563076 35820 563080
rect 46796 563136 46860 563140
rect 46796 563080 46810 563136
rect 46810 563080 46860 563136
rect 46796 563076 46860 563080
rect 48094 561776 48158 561780
rect 48094 561720 48098 561776
rect 48098 561720 48158 561776
rect 48094 561716 48158 561720
rect 341564 543144 341628 543148
rect 341564 543088 341614 543144
rect 341614 543088 341628 543144
rect 341564 543084 341628 543088
rect 337148 542948 337212 543012
rect 338988 542948 339052 543012
rect 528324 540228 528388 540292
rect 198596 539684 198660 539748
rect 216812 539684 216876 539748
rect 529060 539684 529124 539748
rect 218100 539608 218164 539612
rect 218100 539552 218114 539608
rect 218114 539552 218164 539608
rect 218100 539548 218164 539552
rect 205772 539200 205836 539204
rect 205772 539144 205786 539200
rect 205786 539144 205836 539200
rect 205772 539140 205836 539144
rect 540836 538792 540900 538796
rect 540836 538736 540850 538792
rect 540850 538736 540900 538792
rect 540836 538732 540900 538736
rect 115414 477804 115478 477868
rect 122622 477864 122686 477868
rect 122622 477808 122654 477864
rect 122654 477808 122686 477864
rect 122622 477804 122686 477808
rect 63172 476172 63236 476236
rect 65748 476172 65812 476236
rect 83044 476172 83108 476236
rect 85620 476172 85684 476236
rect 105676 476172 105740 476236
rect 113036 476172 113100 476236
rect 129596 476172 129660 476236
rect 131988 476172 132052 476236
rect 133092 476172 133156 476236
rect 143396 476172 143460 476236
rect 95372 476036 95436 476100
rect 167132 476172 167196 476236
rect 147076 476036 147140 476100
rect 148364 476096 148428 476100
rect 148364 476040 148378 476096
rect 148378 476040 148428 476096
rect 148364 476036 148428 476040
rect 122604 475764 122668 475828
rect 141188 475764 141252 475828
rect 42748 475552 42812 475556
rect 42748 475496 42798 475552
rect 42798 475496 42812 475552
rect 42748 475492 42812 475496
rect 120212 475492 120276 475556
rect 124812 475492 124876 475556
rect 43668 475356 43732 475420
rect 128492 475356 128556 475420
rect 150572 475492 150636 475556
rect 196388 475356 196452 475420
rect 126284 475220 126348 475284
rect 130700 475220 130764 475284
rect 138244 475220 138308 475284
rect 199516 475220 199580 475284
rect 127204 475084 127268 475148
rect 132724 475084 132788 475148
rect 198044 475084 198108 475148
rect 108068 474948 108132 475012
rect 110092 474948 110156 475012
rect 110460 474948 110524 475012
rect 113772 474948 113836 475012
rect 117820 474948 117884 475012
rect 121316 475008 121380 475012
rect 121316 474952 121366 475008
rect 121366 474952 121380 475008
rect 121316 474948 121380 474952
rect 135300 474948 135364 475012
rect 199332 474948 199396 475012
rect 60596 474872 60660 474876
rect 60596 474816 60646 474872
rect 60646 474816 60660 474872
rect 60596 474812 60660 474816
rect 68140 474812 68204 474876
rect 70716 474812 70780 474876
rect 73660 474812 73724 474876
rect 75316 474812 75380 474876
rect 78076 474812 78140 474876
rect 80652 474812 80716 474876
rect 88196 474872 88260 474876
rect 88196 474816 88246 474872
rect 88246 474816 88260 474872
rect 88196 474812 88260 474816
rect 90772 474812 90836 474876
rect 93716 474872 93780 474876
rect 93716 474816 93766 474872
rect 93766 474816 93780 474872
rect 93716 474812 93780 474816
rect 98316 474812 98380 474876
rect 100524 474812 100588 474876
rect 102732 474812 102796 474876
rect 107332 474812 107396 474876
rect 108436 474812 108500 474876
rect 110828 474812 110892 474876
rect 112668 474812 112732 474876
rect 114324 474812 114388 474876
rect 115244 474812 115308 474876
rect 116716 474812 116780 474876
rect 118372 474812 118436 474876
rect 118924 474812 118988 474876
rect 120580 474812 120644 474876
rect 123708 474812 123772 474876
rect 125364 474812 125428 474876
rect 128124 474812 128188 474876
rect 130516 474812 130580 474876
rect 134196 474812 134260 474876
rect 136220 474812 136284 474876
rect 136588 474872 136652 474876
rect 136588 474816 136602 474872
rect 136602 474816 136652 474872
rect 136588 474812 136652 474816
rect 137876 474872 137940 474876
rect 137876 474816 137926 474872
rect 137926 474816 137940 474872
rect 137876 474812 137940 474816
rect 138980 474812 139044 474876
rect 140084 474812 140148 474876
rect 142660 474812 142724 474876
rect 150020 474812 150084 474876
rect 197860 474812 197924 474876
rect 338436 462028 338500 462092
rect 338436 461484 338500 461548
rect 168972 455772 169036 455836
rect 198964 455636 199028 455700
rect 197308 455500 197372 455564
rect 198780 454004 198844 454068
rect 288950 453792 289014 453796
rect 288950 453736 288954 453792
rect 288954 453736 289014 453792
rect 288950 453732 289014 453736
rect 294798 453792 294862 453796
rect 294798 453736 294842 453792
rect 294842 453736 294862 453792
rect 294798 453732 294862 453736
rect 429590 453732 429654 453796
rect 430542 453732 430606 453796
rect 431766 453732 431830 453796
rect 213334 453596 213398 453660
rect 284326 453656 284390 453660
rect 284326 453600 284354 453656
rect 284354 453600 284390 453656
rect 284326 453596 284390 453600
rect 286774 453656 286838 453660
rect 286774 453600 286782 453656
rect 286782 453600 286838 453656
rect 286774 453596 286838 453600
rect 290174 453656 290238 453660
rect 290174 453600 290186 453656
rect 290186 453600 290238 453656
rect 290174 453596 290238 453600
rect 291262 453596 291326 453660
rect 293710 453656 293774 453660
rect 293710 453600 293738 453656
rect 293738 453600 293774 453656
rect 293710 453596 293774 453600
rect 297110 453656 297174 453660
rect 297110 453600 297142 453656
rect 297142 453600 297174 453656
rect 297110 453596 297174 453600
rect 298470 453656 298534 453660
rect 298470 453600 298522 453656
rect 298522 453600 298534 453656
rect 298470 453596 298534 453600
rect 299558 453656 299622 453660
rect 299558 453600 299570 453656
rect 299570 453600 299622 453656
rect 299558 453596 299622 453600
rect 311118 453656 311182 453660
rect 311118 453600 311126 453656
rect 311126 453600 311182 453656
rect 311118 453596 311182 453600
rect 312342 453656 312406 453660
rect 312342 453600 312358 453656
rect 312358 453600 312406 453656
rect 312342 453596 312406 453600
rect 443598 453656 443662 453660
rect 443598 453600 443642 453656
rect 443642 453600 443662 453656
rect 443598 453596 443662 453600
rect 532740 453596 532804 453660
rect 533222 453596 533286 453660
rect 196388 453188 196452 453252
rect 199516 453052 199580 453116
rect 279556 453052 279620 453116
rect 199332 452916 199396 452980
rect 285260 452916 285324 452980
rect 198044 452780 198108 452844
rect 295932 452780 295996 452844
rect 197860 452644 197924 452708
rect 35204 452508 35268 452572
rect 230612 452508 230676 452572
rect 233188 452508 233252 452572
rect 235580 452508 235644 452572
rect 238156 452508 238220 452572
rect 240732 452508 240796 452572
rect 243124 452568 243188 452572
rect 243124 452512 243174 452568
rect 243174 452512 243188 452568
rect 243124 452508 243188 452512
rect 245516 452568 245580 452572
rect 245516 452512 245566 452568
rect 245566 452512 245580 452568
rect 245516 452508 245580 452512
rect 253060 452508 253124 452572
rect 255636 452568 255700 452572
rect 255636 452512 255686 452568
rect 255686 452512 255700 452568
rect 255636 452508 255700 452512
rect 260604 452508 260668 452572
rect 263180 452508 263244 452572
rect 265572 452568 265636 452572
rect 265572 452512 265622 452568
rect 265622 452512 265636 452568
rect 265572 452508 265636 452512
rect 268332 452508 268396 452572
rect 270540 452508 270604 452572
rect 273116 452568 273180 452572
rect 273116 452512 273166 452568
rect 273166 452512 273180 452568
rect 273116 452508 273180 452512
rect 275692 452508 275756 452572
rect 278084 452508 278148 452572
rect 280476 452508 280540 452572
rect 282132 452568 282196 452572
rect 282132 452512 282146 452568
rect 282146 452512 282196 452568
rect 282132 452508 282196 452512
rect 283052 452508 283116 452572
rect 285628 452568 285692 452572
rect 285628 452512 285642 452568
rect 285642 452512 285692 452568
rect 285628 452508 285692 452512
rect 288204 452508 288268 452572
rect 290596 452508 290660 452572
rect 292620 452568 292684 452572
rect 292620 452512 292634 452568
rect 292634 452512 292684 452568
rect 292620 452508 292684 452512
rect 292988 452568 293052 452572
rect 292988 452512 293038 452568
rect 293038 452512 293052 452568
rect 292988 452508 293052 452512
rect 295564 452508 295628 452572
rect 298140 452508 298204 452572
rect 300348 452508 300412 452572
rect 302004 452568 302068 452572
rect 302004 452512 302018 452568
rect 302018 452512 302068 452568
rect 302004 452508 302068 452512
rect 303108 452568 303172 452572
rect 303108 452512 303122 452568
rect 303122 452512 303172 452568
rect 303108 452508 303172 452512
rect 304212 452568 304276 452572
rect 304212 452512 304226 452568
rect 304226 452512 304276 452568
rect 304212 452508 304276 452512
rect 305316 452568 305380 452572
rect 305316 452512 305330 452568
rect 305330 452512 305380 452568
rect 305316 452508 305380 452512
rect 306420 452568 306484 452572
rect 306420 452512 306434 452568
rect 306434 452512 306484 452568
rect 306420 452508 306484 452512
rect 307892 452568 307956 452572
rect 307892 452512 307906 452568
rect 307906 452512 307956 452568
rect 307892 452508 307956 452512
rect 308996 452568 309060 452572
rect 308996 452512 309010 452568
rect 309010 452512 309060 452568
rect 308996 452508 309060 452512
rect 309916 452568 309980 452572
rect 309916 452512 309930 452568
rect 309930 452512 309980 452568
rect 309916 452508 309980 452512
rect 313412 452568 313476 452572
rect 313412 452512 313426 452568
rect 313426 452512 313476 452568
rect 313412 452508 313476 452512
rect 314700 452568 314764 452572
rect 314700 452512 314714 452568
rect 314714 452512 314764 452568
rect 314700 452508 314764 452512
rect 315988 452508 316052 452572
rect 316908 452508 316972 452572
rect 318380 452508 318444 452572
rect 320404 452508 320468 452572
rect 426020 452508 426084 452572
rect 427124 452508 427188 452572
rect 428228 452508 428292 452572
rect 429516 452508 429580 452572
rect 433012 452508 433076 452572
rect 434116 452508 434180 452572
rect 435404 452508 435468 452572
rect 436508 452508 436572 452572
rect 450676 452508 450740 452572
rect 452884 452568 452948 452572
rect 452884 452512 452898 452568
rect 452898 452512 452948 452568
rect 452884 452508 452948 452512
rect 466132 452568 466196 452572
rect 466132 452512 466182 452568
rect 466182 452512 466196 452568
rect 466132 452508 466196 452512
rect 467052 452508 467116 452572
rect 467972 452568 468036 452572
rect 467972 452512 467986 452568
rect 467986 452512 468036 452568
rect 467972 452508 468036 452512
rect 468524 452508 468588 452572
rect 470916 452508 470980 452572
rect 473492 452568 473556 452572
rect 473492 452512 473542 452568
rect 473542 452512 473556 452568
rect 473492 452508 473556 452512
rect 476068 452568 476132 452572
rect 476068 452512 476082 452568
rect 476082 452512 476132 452568
rect 476068 452508 476132 452512
rect 478276 452508 478340 452572
rect 481036 452568 481100 452572
rect 481036 452512 481086 452568
rect 481086 452512 481100 452568
rect 481036 452508 481100 452512
rect 483428 452568 483492 452572
rect 483428 452512 483478 452568
rect 483478 452512 483492 452568
rect 483428 452508 483492 452512
rect 486004 452508 486068 452572
rect 488396 452568 488460 452572
rect 488396 452512 488446 452568
rect 488446 452512 488460 452568
rect 488396 452508 488460 452512
rect 490972 452568 491036 452572
rect 490972 452512 491022 452568
rect 491022 452512 491036 452568
rect 490972 452508 491036 452512
rect 493548 452568 493612 452572
rect 493548 452512 493598 452568
rect 493598 452512 493612 452568
rect 493548 452508 493612 452512
rect 495940 452568 496004 452572
rect 495940 452512 495990 452568
rect 495990 452512 496004 452568
rect 495940 452508 496004 452512
rect 498516 452508 498580 452572
rect 501092 452508 501156 452572
rect 503484 452568 503548 452572
rect 503484 452512 503534 452568
rect 503534 452512 503548 452568
rect 503484 452508 503548 452512
rect 505876 452568 505940 452572
rect 505876 452512 505926 452568
rect 505926 452512 505940 452568
rect 505876 452508 505940 452512
rect 508452 452508 508516 452572
rect 511028 452508 511092 452572
rect 513420 452508 513484 452572
rect 515996 452568 516060 452572
rect 515996 452512 516046 452568
rect 516046 452512 516060 452568
rect 515996 452508 516060 452512
rect 213316 452432 213380 452436
rect 213316 452376 213366 452432
rect 213366 452376 213380 452432
rect 213316 452372 213380 452376
rect 533292 452372 533356 452436
rect 198964 452236 199028 452300
rect 280844 452236 280908 452300
rect 283236 452296 283300 452300
rect 283236 452240 283250 452296
rect 283250 452240 283300 452296
rect 283236 452236 283300 452240
rect 197308 452100 197372 452164
rect 277164 452100 277228 452164
rect 287836 452236 287900 452300
rect 300716 452236 300780 452300
rect 302924 452236 302988 452300
rect 305868 452236 305932 452300
rect 319484 452296 319548 452300
rect 319484 452240 319498 452296
rect 319498 452240 319548 452296
rect 319484 452236 319548 452240
rect 438348 452236 438412 452300
rect 455276 452236 455340 452300
rect 463372 452236 463436 452300
rect 469076 452236 469140 452300
rect 442396 452100 442460 452164
rect 443500 452100 443564 452164
rect 445892 452100 445956 452164
rect 446076 452100 446140 452164
rect 449388 452100 449452 452164
rect 451780 452100 451844 452164
rect 453620 452160 453684 452164
rect 453620 452104 453670 452160
rect 453670 452104 453684 452160
rect 453620 452100 453684 452104
rect 456012 452100 456076 452164
rect 459692 452160 459756 452164
rect 459692 452104 459742 452160
rect 459742 452104 459756 452160
rect 459692 452100 459756 452104
rect 462268 452100 462332 452164
rect 463556 452160 463620 452164
rect 463556 452104 463606 452160
rect 463606 452104 463620 452160
rect 463556 452100 463620 452104
rect 465764 452100 465828 452164
rect 198780 451964 198844 452028
rect 46796 451828 46860 451892
rect 167500 451828 167564 451892
rect 278452 451828 278516 451892
rect 438716 451556 438780 451620
rect 441292 451556 441356 451620
rect 458404 451556 458468 451620
rect 532740 451420 532804 451484
rect 48084 451344 48148 451348
rect 48084 451288 48098 451344
rect 48098 451288 48148 451344
rect 48084 451284 48148 451288
rect 248092 451284 248156 451348
rect 250668 451284 250732 451348
rect 258028 451284 258092 451348
rect 308260 451284 308324 451348
rect 437612 451344 437676 451348
rect 437612 451288 437626 451344
rect 437626 451288 437676 451344
rect 437612 451284 437676 451288
rect 440004 451284 440068 451348
rect 440740 451284 440804 451348
rect 444604 451284 444668 451348
rect 446996 451284 447060 451348
rect 448100 451284 448164 451348
rect 448468 451344 448532 451348
rect 448468 451288 448518 451344
rect 448518 451288 448532 451344
rect 448468 451284 448532 451288
rect 451044 451284 451108 451348
rect 453988 451284 454052 451348
rect 456380 451284 456444 451348
rect 457668 451284 457732 451348
rect 458588 451284 458652 451348
rect 464292 451284 464356 451348
rect 170444 451148 170508 451212
rect 167132 449924 167196 449988
rect 461164 449244 461228 449308
rect 460980 449108 461044 449172
rect 168604 448564 168668 448628
rect 174676 447884 174740 447948
rect 338252 447884 338316 447948
rect 336964 447748 337028 447812
rect 336780 447612 336844 447676
rect 338068 439452 338132 439516
rect 174492 438092 174556 438156
rect 196572 432516 196636 432580
rect 341564 428088 341628 428092
rect 341564 428032 341614 428088
rect 341614 428032 341628 428088
rect 341564 428028 341628 428032
rect 170628 427620 170692 427684
rect 338436 425716 338500 425780
rect 166948 425580 167012 425644
rect 170076 423600 170140 423604
rect 170076 423544 170126 423600
rect 170126 423544 170140 423600
rect 170076 423540 170140 423544
rect 198780 422860 198844 422924
rect 337148 421772 337212 421836
rect 338988 421772 339052 421836
rect 340092 421832 340156 421836
rect 340092 421776 340106 421832
rect 340106 421776 340156 421832
rect 340092 421772 340156 421776
rect 171548 421228 171612 421292
rect 170260 421092 170324 421156
rect 167684 420956 167748 421020
rect 168604 420956 168668 421020
rect 174676 420956 174740 421020
rect 174492 419596 174556 419660
rect 168420 382332 168484 382396
rect 168236 379476 168300 379540
rect 43116 364244 43180 364308
rect 112116 364244 112180 364308
rect 115428 364244 115492 364308
rect 132908 364304 132972 364308
rect 132908 364248 132958 364304
rect 132958 364248 132972 364304
rect 132908 364244 132972 364248
rect 135300 364244 135364 364308
rect 143396 364304 143460 364308
rect 143396 364248 143410 364304
rect 143410 364248 143460 364304
rect 143396 364244 143460 364248
rect 144684 364244 144748 364308
rect 145972 364244 146036 364308
rect 43484 364108 43548 364172
rect 63172 364108 63236 364172
rect 65748 364108 65812 364172
rect 73108 364168 73172 364172
rect 73108 364112 73158 364168
rect 73158 364112 73172 364168
rect 73108 364108 73172 364112
rect 75684 364108 75748 364172
rect 83044 364108 83108 364172
rect 85620 364168 85684 364172
rect 85620 364112 85670 364168
rect 85670 364112 85684 364168
rect 85620 364108 85684 364112
rect 93164 364108 93228 364172
rect 95556 364168 95620 364172
rect 95556 364112 95606 364168
rect 95606 364112 95620 364168
rect 95556 364108 95620 364112
rect 103100 364168 103164 364172
rect 103100 364112 103150 364168
rect 103150 364112 103164 364168
rect 103100 364108 103164 364112
rect 105676 364108 105740 364172
rect 109540 364168 109604 364172
rect 109540 364112 109590 364168
rect 109590 364112 109604 364168
rect 109540 364108 109604 364112
rect 113036 364168 113100 364172
rect 113036 364112 113086 364168
rect 113086 364112 113100 364168
rect 113036 364108 113100 364112
rect 113220 364108 113284 364172
rect 115612 364108 115676 364172
rect 122972 364108 123036 364172
rect 125916 364168 125980 364172
rect 125916 364112 125966 364168
rect 125966 364112 125980 364168
rect 125916 364108 125980 364112
rect 129596 364168 129660 364172
rect 129596 364112 129610 364168
rect 129610 364112 129660 364168
rect 129596 364108 129660 364112
rect 131988 364168 132052 364172
rect 131988 364112 132038 364168
rect 132038 364112 132052 364168
rect 131988 364108 132052 364112
rect 133092 364168 133156 364172
rect 133092 364112 133142 364168
rect 133142 364112 133156 364168
rect 133092 364108 133156 364112
rect 135852 364168 135916 364172
rect 135852 364112 135902 364168
rect 135902 364112 135916 364168
rect 135852 364108 135916 364112
rect 142292 364108 142356 364172
rect 149468 364108 149532 364172
rect 167132 364168 167196 364172
rect 167132 364112 167182 364168
rect 167182 364112 167196 364168
rect 167132 364108 167196 364112
rect 120212 363972 120276 364036
rect 170628 363972 170692 364036
rect 122604 363836 122668 363900
rect 136588 363896 136652 363900
rect 136588 363840 136602 363896
rect 136602 363840 136652 363896
rect 136588 363836 136652 363840
rect 127204 363700 127268 363764
rect 166948 363836 167012 363900
rect 150572 363564 150636 363628
rect 123708 363428 123772 363492
rect 138244 363488 138308 363492
rect 138244 363432 138294 363488
rect 138294 363432 138308 363488
rect 138244 363428 138308 363432
rect 108068 363292 108132 363356
rect 118924 363292 118988 363356
rect 167132 363292 167196 363356
rect 110460 363156 110524 363220
rect 117820 363156 117884 363220
rect 120580 363156 120644 363220
rect 124812 363156 124876 363220
rect 130700 363156 130764 363220
rect 60596 363080 60660 363084
rect 60596 363024 60646 363080
rect 60646 363024 60660 363080
rect 60596 363020 60660 363024
rect 68140 363020 68204 363084
rect 70716 363020 70780 363084
rect 78076 363020 78140 363084
rect 80652 363020 80716 363084
rect 88196 363080 88260 363084
rect 88196 363024 88246 363080
rect 88246 363024 88260 363080
rect 88196 363020 88260 363024
rect 90772 363020 90836 363084
rect 98316 363020 98380 363084
rect 100524 363020 100588 363084
rect 107332 363020 107396 363084
rect 108436 363020 108500 363084
rect 110828 363020 110892 363084
rect 114324 363080 114388 363084
rect 114324 363024 114374 363080
rect 114374 363024 114388 363080
rect 114324 363020 114388 363024
rect 116716 363020 116780 363084
rect 118372 363020 118436 363084
rect 121316 363020 121380 363084
rect 125364 363080 125428 363084
rect 125364 363024 125414 363080
rect 125414 363024 125428 363080
rect 125364 363020 125428 363024
rect 128124 363080 128188 363084
rect 128124 363024 128174 363080
rect 128174 363024 128188 363080
rect 128124 363020 128188 363024
rect 128492 363020 128556 363084
rect 130516 363020 130580 363084
rect 134196 363020 134260 363084
rect 137876 363080 137940 363084
rect 137876 363024 137926 363080
rect 137926 363024 137940 363080
rect 137876 363020 137940 363024
rect 138980 363020 139044 363084
rect 140084 363020 140148 363084
rect 141188 363020 141252 363084
rect 148364 363020 148428 363084
rect 170444 361660 170508 361724
rect 168604 353228 168668 353292
rect 168604 352548 168668 352612
rect 172652 342892 172716 342956
rect 48084 340716 48148 340780
rect 46796 340172 46860 340236
rect 174676 340036 174740 340100
rect 35204 339552 35268 339556
rect 35204 339496 35218 339552
rect 35218 339496 35268 339552
rect 35204 339492 35268 339496
rect 168052 259524 168116 259588
rect 60606 253736 60670 253740
rect 60606 253680 60646 253736
rect 60646 253680 60670 253736
rect 60606 253676 60670 253680
rect 65638 253676 65702 253740
rect 70670 253736 70734 253740
rect 70670 253680 70674 253736
rect 70674 253680 70730 253736
rect 70730 253680 70734 253736
rect 70670 253676 70734 253680
rect 75566 253736 75630 253740
rect 75566 253680 75606 253736
rect 75606 253680 75630 253736
rect 75566 253676 75630 253680
rect 98278 253736 98342 253740
rect 98278 253680 98330 253736
rect 98330 253680 98342 253736
rect 98278 253676 98342 253680
rect 115612 253736 115676 253740
rect 115612 253680 115662 253736
rect 115662 253680 115676 253736
rect 115612 253676 115676 253680
rect 118270 253736 118334 253740
rect 118270 253680 118330 253736
rect 118330 253680 118334 253736
rect 118270 253676 118334 253680
rect 123030 253736 123094 253740
rect 123030 253680 123078 253736
rect 123078 253680 123094 253736
rect 123030 253676 123094 253680
rect 125478 253736 125542 253740
rect 125478 253680 125506 253736
rect 125506 253680 125542 253736
rect 125478 253676 125542 253680
rect 128062 253736 128126 253740
rect 128062 253680 128082 253736
rect 128082 253680 128126 253736
rect 128062 253676 128126 253680
rect 43334 253600 43398 253604
rect 43334 253544 43350 253600
rect 43350 253544 43398 253600
rect 43334 253540 43398 253544
rect 130516 253600 130580 253604
rect 130516 253544 130566 253600
rect 130566 253544 130580 253600
rect 130516 253540 130580 253544
rect 136494 253600 136558 253604
rect 136494 253544 136510 253600
rect 136510 253544 136558 253600
rect 136494 253540 136558 253544
rect 132908 253464 132972 253468
rect 132908 253408 132958 253464
rect 132958 253408 132972 253464
rect 132908 253404 132972 253408
rect 63172 252452 63236 252516
rect 68140 252512 68204 252516
rect 68140 252456 68190 252512
rect 68190 252456 68204 252512
rect 68140 252452 68204 252456
rect 73108 252512 73172 252516
rect 73108 252456 73158 252512
rect 73158 252456 73172 252512
rect 73108 252452 73172 252456
rect 78076 252512 78140 252516
rect 78076 252456 78126 252512
rect 78126 252456 78140 252512
rect 78076 252452 78140 252456
rect 80652 252452 80716 252516
rect 83044 252452 83108 252516
rect 85620 252512 85684 252516
rect 85620 252456 85670 252512
rect 85670 252456 85684 252512
rect 85620 252452 85684 252456
rect 88196 252512 88260 252516
rect 88196 252456 88246 252512
rect 88246 252456 88260 252512
rect 88196 252452 88260 252456
rect 90772 252512 90836 252516
rect 90772 252456 90822 252512
rect 90822 252456 90836 252512
rect 90772 252452 90836 252456
rect 93164 252512 93228 252516
rect 93164 252456 93214 252512
rect 93214 252456 93228 252512
rect 93164 252452 93228 252456
rect 95556 252512 95620 252516
rect 95556 252456 95606 252512
rect 95606 252456 95620 252512
rect 95556 252452 95620 252456
rect 100524 252512 100588 252516
rect 100524 252456 100574 252512
rect 100574 252456 100588 252512
rect 100524 252452 100588 252456
rect 103100 252512 103164 252516
rect 103100 252456 103150 252512
rect 103150 252456 103164 252512
rect 103100 252452 103164 252456
rect 105676 252452 105740 252516
rect 108068 252452 108132 252516
rect 110460 252512 110524 252516
rect 110460 252456 110510 252512
rect 110510 252456 110524 252512
rect 110460 252452 110524 252456
rect 113036 252512 113100 252516
rect 113036 252456 113086 252512
rect 113086 252456 113100 252512
rect 113036 252452 113100 252456
rect 115428 252452 115492 252516
rect 120580 252452 120644 252516
rect 135852 252452 135916 252516
rect 143396 252512 143460 252516
rect 143396 252456 143410 252512
rect 143410 252456 143460 252512
rect 143396 252452 143460 252456
rect 144868 252452 144932 252516
rect 145972 252452 146036 252516
rect 147076 252452 147140 252516
rect 148364 252512 148428 252516
rect 148364 252456 148378 252512
rect 148378 252456 148428 252512
rect 148364 252452 148428 252456
rect 150572 252452 150636 252516
rect 43116 252316 43180 252380
rect 109540 252316 109604 252380
rect 110828 252316 110892 252380
rect 112116 252316 112180 252380
rect 113220 252316 113284 252380
rect 125916 252316 125980 252380
rect 129596 252376 129660 252380
rect 129596 252320 129610 252376
rect 129610 252320 129660 252376
rect 129596 252316 129660 252320
rect 131988 252376 132052 252380
rect 131988 252320 132038 252376
rect 132038 252320 132052 252376
rect 131988 252316 132052 252320
rect 133092 252316 133156 252380
rect 138244 252376 138308 252380
rect 138244 252320 138294 252376
rect 138294 252320 138308 252376
rect 138244 252316 138308 252320
rect 142292 252316 142356 252380
rect 168052 252180 168116 252244
rect 150020 252044 150084 252108
rect 114324 251968 114388 251972
rect 114324 251912 114374 251968
rect 114374 251912 114388 251968
rect 114324 251908 114388 251912
rect 141188 251908 141252 251972
rect 120212 251636 120276 251700
rect 135300 251636 135364 251700
rect 107332 251228 107396 251292
rect 108436 251228 108500 251292
rect 116716 251228 116780 251292
rect 117820 251228 117884 251292
rect 118924 251228 118988 251292
rect 121316 251288 121380 251292
rect 121316 251232 121330 251288
rect 121330 251232 121380 251288
rect 121316 251228 121380 251232
rect 122604 251228 122668 251292
rect 123708 251228 123772 251292
rect 124812 251228 124876 251292
rect 127204 251228 127268 251292
rect 128492 251228 128556 251292
rect 130700 251228 130764 251292
rect 134196 251228 134260 251292
rect 137876 251288 137940 251292
rect 137876 251232 137926 251288
rect 137926 251232 137940 251288
rect 137876 251228 137940 251232
rect 138980 251228 139044 251292
rect 140084 251228 140148 251292
rect 198596 250412 198660 250476
rect 198780 247964 198844 248028
rect 167500 245652 167564 245716
rect 168236 238640 168300 238644
rect 168236 238584 168250 238640
rect 168250 238584 168300 238640
rect 168236 238580 168300 238584
rect 168972 228924 169036 228988
rect 35204 227760 35268 227764
rect 35204 227704 35218 227760
rect 35218 227704 35268 227760
rect 35204 227700 35268 227704
rect 46796 227760 46860 227764
rect 46796 227704 46810 227760
rect 46810 227704 46860 227760
rect 46796 227700 46860 227704
rect 48084 227700 48148 227764
rect 170260 227020 170324 227084
rect 171548 226884 171612 226948
rect 123030 141748 123094 141812
rect 133094 141808 133158 141812
rect 133094 141752 133142 141808
rect 133142 141752 133158 141808
rect 133094 141748 133158 141752
rect 108478 141672 108542 141676
rect 108478 141616 108486 141672
rect 108486 141616 108542 141672
rect 108478 141612 108542 141616
rect 112150 141672 112214 141676
rect 112150 141616 112166 141672
rect 112166 141616 112214 141672
rect 112150 141612 112214 141616
rect 123710 141672 123774 141676
rect 123710 141616 123758 141672
rect 123758 141616 123774 141672
rect 123710 141612 123774 141616
rect 128470 141612 128534 141676
rect 134182 141612 134246 141676
rect 136494 141672 136558 141676
rect 136494 141616 136546 141672
rect 136546 141616 136558 141672
rect 136494 141612 136558 141616
rect 140030 141672 140094 141676
rect 140030 141616 140042 141672
rect 140042 141616 140094 141672
rect 140030 141612 140094 141616
rect 142342 141672 142406 141676
rect 142342 141616 142398 141672
rect 142398 141616 142406 141672
rect 142342 141612 142406 141616
rect 109540 140720 109604 140724
rect 109540 140664 109590 140720
rect 109590 140664 109604 140720
rect 109540 140660 109604 140664
rect 113220 140720 113284 140724
rect 113220 140664 113270 140720
rect 113270 140664 113284 140720
rect 113220 140660 113284 140664
rect 116716 140720 116780 140724
rect 116716 140664 116766 140720
rect 116766 140664 116780 140720
rect 116716 140660 116780 140664
rect 118924 140720 118988 140724
rect 118924 140664 118974 140720
rect 118974 140664 118988 140720
rect 118924 140660 118988 140664
rect 125916 140720 125980 140724
rect 125916 140664 125966 140720
rect 125966 140664 125980 140720
rect 125916 140660 125980 140664
rect 131988 140720 132052 140724
rect 131988 140664 132038 140720
rect 132038 140664 132052 140720
rect 131988 140660 132052 140664
rect 135300 140720 135364 140724
rect 135300 140664 135350 140720
rect 135350 140664 135364 140720
rect 135300 140660 135364 140664
rect 137876 140720 137940 140724
rect 137876 140664 137926 140720
rect 137926 140664 137940 140720
rect 137876 140660 137940 140664
rect 138980 140720 139044 140724
rect 138980 140664 139030 140720
rect 139030 140664 139044 140720
rect 138980 140660 139044 140664
rect 141188 140720 141252 140724
rect 141188 140664 141238 140720
rect 141238 140664 141252 140720
rect 141188 140660 141252 140664
rect 143396 140720 143460 140724
rect 143396 140664 143446 140720
rect 143446 140664 143460 140720
rect 143396 140660 143460 140664
rect 149468 140720 149532 140724
rect 149468 140664 149518 140720
rect 149518 140664 149532 140720
rect 149468 140660 149532 140664
rect 43116 140176 43180 140180
rect 43116 140120 43130 140176
rect 43130 140120 43180 140176
rect 43116 140116 43180 140120
rect 63172 140176 63236 140180
rect 63172 140120 63222 140176
rect 63222 140120 63236 140176
rect 63172 140116 63236 140120
rect 65748 140176 65812 140180
rect 65748 140120 65798 140176
rect 65798 140120 65812 140176
rect 65748 140116 65812 140120
rect 115428 140176 115492 140180
rect 115428 140120 115478 140176
rect 115478 140120 115492 140176
rect 115428 140116 115492 140120
rect 115612 140116 115676 140180
rect 129596 140176 129660 140180
rect 129596 140120 129646 140176
rect 129646 140120 129660 140176
rect 129596 140116 129660 140120
rect 43668 139300 43732 139364
rect 60596 139360 60660 139364
rect 60596 139304 60646 139360
rect 60646 139304 60660 139360
rect 60596 139300 60660 139304
rect 107332 139360 107396 139364
rect 107332 139304 107382 139360
rect 107382 139304 107396 139360
rect 107332 139300 107396 139304
rect 110828 139360 110892 139364
rect 110828 139304 110878 139360
rect 110878 139304 110892 139360
rect 110828 139300 110892 139304
rect 114324 139360 114388 139364
rect 114324 139304 114374 139360
rect 114374 139304 114388 139360
rect 114324 139300 114388 139304
rect 117820 139360 117884 139364
rect 117820 139304 117870 139360
rect 117870 139304 117884 139360
rect 117820 139300 117884 139304
rect 120212 139300 120276 139364
rect 121316 139360 121380 139364
rect 121316 139304 121366 139360
rect 121366 139304 121380 139360
rect 121316 139300 121380 139304
rect 122604 139360 122668 139364
rect 122604 139304 122654 139360
rect 122654 139304 122668 139360
rect 122604 139300 122668 139304
rect 124812 139300 124876 139364
rect 127204 139300 127268 139364
rect 130700 139360 130764 139364
rect 130700 139304 130750 139360
rect 130750 139304 130764 139360
rect 130700 139300 130764 139304
rect 148364 139360 148428 139364
rect 148364 139304 148414 139360
rect 148414 139304 148428 139360
rect 148364 139300 148428 139304
rect 150572 139300 150636 139364
rect 136220 139028 136284 139092
rect 68140 138620 68204 138684
rect 70716 138076 70780 138140
rect 73660 138076 73724 138140
rect 75316 138076 75380 138140
rect 78076 138076 78140 138140
rect 80652 138076 80716 138140
rect 83780 138076 83844 138140
rect 86356 138076 86420 138140
rect 88196 138136 88260 138140
rect 88196 138080 88246 138136
rect 88246 138080 88260 138136
rect 88196 138076 88260 138080
rect 90772 138076 90836 138140
rect 93716 138136 93780 138140
rect 93716 138080 93766 138136
rect 93766 138080 93780 138136
rect 93716 138076 93780 138080
rect 96292 138076 96356 138140
rect 98316 138076 98380 138140
rect 100524 138076 100588 138140
rect 102732 138076 102796 138140
rect 105308 138076 105372 138140
rect 108068 138076 108132 138140
rect 110460 138076 110524 138140
rect 112668 138076 112732 138140
rect 118372 138136 118436 138140
rect 118372 138080 118422 138136
rect 118422 138080 118436 138136
rect 118372 138076 118436 138080
rect 120580 138076 120644 138140
rect 125364 138136 125428 138140
rect 125364 138080 125414 138136
rect 125414 138080 125428 138136
rect 125364 138076 125428 138080
rect 128124 138076 128188 138140
rect 130516 138076 130580 138140
rect 132724 138076 132788 138140
rect 138244 138076 138308 138140
rect 35204 117132 35268 117196
rect 46796 116996 46860 117060
rect 48084 116724 48148 116788
rect 125478 29820 125542 29884
rect 75566 29608 75630 29612
rect 75566 29552 75606 29608
rect 75606 29552 75630 29608
rect 75566 29548 75630 29552
rect 88078 29608 88142 29612
rect 88078 29552 88118 29608
rect 88118 29552 88142 29608
rect 88078 29548 88142 29552
rect 90662 29548 90726 29612
rect 123710 29548 123774 29612
rect 130510 29608 130574 29612
rect 130510 29552 130566 29608
rect 130566 29552 130574 29608
rect 130510 29548 130574 29552
rect 138942 29608 139006 29612
rect 138942 29552 138994 29608
rect 138994 29552 139006 29608
rect 138942 29548 139006 29552
rect 60596 28928 60660 28932
rect 60596 28872 60646 28928
rect 60646 28872 60660 28928
rect 60596 28868 60660 28872
rect 68140 28928 68204 28932
rect 68140 28872 68190 28928
rect 68190 28872 68204 28928
rect 68140 28868 68204 28872
rect 78076 28928 78140 28932
rect 78076 28872 78126 28928
rect 78126 28872 78140 28928
rect 78076 28868 78140 28872
rect 80652 28928 80716 28932
rect 80652 28872 80702 28928
rect 80702 28872 80716 28928
rect 80652 28868 80716 28872
rect 83044 28928 83108 28932
rect 83044 28872 83094 28928
rect 83094 28872 83108 28928
rect 83044 28868 83108 28872
rect 103100 28928 103164 28932
rect 103100 28872 103150 28928
rect 103150 28872 103164 28928
rect 103100 28868 103164 28872
rect 128492 28928 128556 28932
rect 128492 28872 128542 28928
rect 128542 28872 128556 28928
rect 128492 28868 128556 28872
rect 134196 28928 134260 28932
rect 134196 28872 134246 28928
rect 134246 28872 134260 28928
rect 134196 28868 134260 28872
rect 135852 28928 135916 28932
rect 135852 28872 135902 28928
rect 135902 28872 135916 28928
rect 135852 28868 135916 28872
rect 138244 28928 138308 28932
rect 138244 28872 138294 28928
rect 138294 28872 138308 28928
rect 138244 28868 138308 28872
rect 133092 28732 133156 28796
rect 135300 28596 135364 28660
rect 63172 28248 63236 28252
rect 63172 28192 63222 28248
rect 63222 28192 63236 28248
rect 63172 28188 63236 28192
rect 112116 28248 112180 28252
rect 112116 28192 112166 28248
rect 112166 28192 112180 28248
rect 112116 28188 112180 28192
rect 115612 28248 115676 28252
rect 115612 28192 115662 28248
rect 115662 28192 115676 28248
rect 115612 28188 115676 28192
rect 129596 28248 129660 28252
rect 129596 28192 129646 28248
rect 129646 28192 129660 28248
rect 129596 28188 129660 28192
rect 131988 28248 132052 28252
rect 131988 28192 132038 28248
rect 132038 28192 132052 28248
rect 131988 28188 132052 28192
rect 143396 28248 143460 28252
rect 143396 28192 143446 28248
rect 143446 28192 143460 28248
rect 143396 28188 143460 28192
rect 42748 27568 42812 27572
rect 42748 27512 42798 27568
rect 42798 27512 42812 27568
rect 42748 27508 42812 27512
rect 43668 27568 43732 27572
rect 43668 27512 43682 27568
rect 43682 27512 43732 27568
rect 43668 27508 43732 27512
rect 64828 27568 64892 27572
rect 64828 27512 64878 27568
rect 64878 27512 64892 27568
rect 64828 27508 64892 27512
rect 70716 27508 70780 27572
rect 73660 27508 73724 27572
rect 86356 27508 86420 27572
rect 92796 27568 92860 27572
rect 92796 27512 92810 27568
rect 92810 27512 92860 27568
rect 92796 27508 92860 27512
rect 95188 27568 95252 27572
rect 95188 27512 95238 27568
rect 95238 27512 95252 27568
rect 95188 27508 95252 27512
rect 98316 27568 98380 27572
rect 98316 27512 98330 27568
rect 98330 27512 98380 27568
rect 98316 27508 98380 27512
rect 100524 27508 100588 27572
rect 105308 27508 105372 27572
rect 107332 27508 107396 27572
rect 108068 27568 108132 27572
rect 108068 27512 108082 27568
rect 108082 27512 108132 27568
rect 108068 27508 108132 27512
rect 108436 27508 108500 27572
rect 110092 27508 110156 27572
rect 110828 27508 110892 27572
rect 112668 27508 112732 27572
rect 116716 27508 116780 27572
rect 117820 27508 117884 27572
rect 118372 27568 118436 27572
rect 118372 27512 118422 27568
rect 118422 27512 118436 27568
rect 118372 27508 118436 27512
rect 120212 27508 120276 27572
rect 126284 27568 126348 27572
rect 126284 27512 126334 27568
rect 126334 27512 126348 27568
rect 126284 27508 126348 27512
rect 128124 27568 128188 27572
rect 128124 27512 128174 27568
rect 128174 27512 128188 27568
rect 128124 27508 128188 27512
rect 132724 27568 132788 27572
rect 132724 27512 132774 27568
rect 132774 27512 132788 27568
rect 132724 27508 132788 27512
rect 136404 27508 136468 27572
rect 137876 27508 137940 27572
rect 140084 27568 140148 27572
rect 140084 27512 140134 27568
rect 140134 27512 140148 27568
rect 140084 27508 140148 27512
rect 141188 27568 141252 27572
rect 141188 27512 141238 27568
rect 141238 27512 141252 27568
rect 141188 27508 141252 27512
rect 147076 27508 147140 27572
rect 148364 27508 148428 27572
rect 150020 27568 150084 27572
rect 150020 27512 150070 27568
rect 150070 27512 150084 27568
rect 150020 27508 150084 27512
rect 150572 27568 150636 27572
rect 150572 27512 150622 27568
rect 150622 27512 150636 27568
rect 150572 27508 150636 27512
rect 110460 27372 110524 27436
rect 121316 27372 121380 27436
rect 120580 27296 120644 27300
rect 120580 27240 120630 27296
rect 120630 27240 120644 27296
rect 120580 27236 120644 27240
rect 113772 27100 113836 27164
rect 114324 26964 114388 27028
rect 123708 27160 123772 27164
rect 123708 27104 123758 27160
rect 123758 27104 123772 27160
rect 123708 27100 123772 27104
rect 127204 27100 127268 27164
rect 124812 26964 124876 27028
rect 122604 26828 122668 26892
rect 130700 26692 130764 26756
rect 142660 26556 142724 26620
rect 115244 26284 115308 26348
rect 118924 26284 118988 26348
rect 174492 5612 174556 5676
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 684274 -8106 711002
rect -8726 684038 -8694 684274
rect -8458 684038 -8374 684274
rect -8138 684038 -8106 684274
rect -8726 664274 -8106 684038
rect -8726 664038 -8694 664274
rect -8458 664038 -8374 664274
rect -8138 664038 -8106 664274
rect -8726 644274 -8106 664038
rect -8726 644038 -8694 644274
rect -8458 644038 -8374 644274
rect -8138 644038 -8106 644274
rect -8726 624274 -8106 644038
rect -8726 624038 -8694 624274
rect -8458 624038 -8374 624274
rect -8138 624038 -8106 624274
rect -8726 604274 -8106 624038
rect -8726 604038 -8694 604274
rect -8458 604038 -8374 604274
rect -8138 604038 -8106 604274
rect -8726 584274 -8106 604038
rect -8726 584038 -8694 584274
rect -8458 584038 -8374 584274
rect -8138 584038 -8106 584274
rect -8726 564274 -8106 584038
rect -8726 564038 -8694 564274
rect -8458 564038 -8374 564274
rect -8138 564038 -8106 564274
rect -8726 544274 -8106 564038
rect -8726 544038 -8694 544274
rect -8458 544038 -8374 544274
rect -8138 544038 -8106 544274
rect -8726 524274 -8106 544038
rect -8726 524038 -8694 524274
rect -8458 524038 -8374 524274
rect -8138 524038 -8106 524274
rect -8726 504274 -8106 524038
rect -8726 504038 -8694 504274
rect -8458 504038 -8374 504274
rect -8138 504038 -8106 504274
rect -8726 484274 -8106 504038
rect -8726 484038 -8694 484274
rect -8458 484038 -8374 484274
rect -8138 484038 -8106 484274
rect -8726 464274 -8106 484038
rect -8726 464038 -8694 464274
rect -8458 464038 -8374 464274
rect -8138 464038 -8106 464274
rect -8726 444274 -8106 464038
rect -8726 444038 -8694 444274
rect -8458 444038 -8374 444274
rect -8138 444038 -8106 444274
rect -8726 424274 -8106 444038
rect -8726 424038 -8694 424274
rect -8458 424038 -8374 424274
rect -8138 424038 -8106 424274
rect -8726 404274 -8106 424038
rect -8726 404038 -8694 404274
rect -8458 404038 -8374 404274
rect -8138 404038 -8106 404274
rect -8726 384274 -8106 404038
rect -8726 384038 -8694 384274
rect -8458 384038 -8374 384274
rect -8138 384038 -8106 384274
rect -8726 364274 -8106 384038
rect -8726 364038 -8694 364274
rect -8458 364038 -8374 364274
rect -8138 364038 -8106 364274
rect -8726 344274 -8106 364038
rect -8726 344038 -8694 344274
rect -8458 344038 -8374 344274
rect -8138 344038 -8106 344274
rect -8726 324274 -8106 344038
rect -8726 324038 -8694 324274
rect -8458 324038 -8374 324274
rect -8138 324038 -8106 324274
rect -8726 304274 -8106 324038
rect -8726 304038 -8694 304274
rect -8458 304038 -8374 304274
rect -8138 304038 -8106 304274
rect -8726 284274 -8106 304038
rect -8726 284038 -8694 284274
rect -8458 284038 -8374 284274
rect -8138 284038 -8106 284274
rect -8726 264274 -8106 284038
rect -8726 264038 -8694 264274
rect -8458 264038 -8374 264274
rect -8138 264038 -8106 264274
rect -8726 244274 -8106 264038
rect -8726 244038 -8694 244274
rect -8458 244038 -8374 244274
rect -8138 244038 -8106 244274
rect -8726 224274 -8106 244038
rect -8726 224038 -8694 224274
rect -8458 224038 -8374 224274
rect -8138 224038 -8106 224274
rect -8726 204274 -8106 224038
rect -8726 204038 -8694 204274
rect -8458 204038 -8374 204274
rect -8138 204038 -8106 204274
rect -8726 184274 -8106 204038
rect -8726 184038 -8694 184274
rect -8458 184038 -8374 184274
rect -8138 184038 -8106 184274
rect -8726 164274 -8106 184038
rect -8726 164038 -8694 164274
rect -8458 164038 -8374 164274
rect -8138 164038 -8106 164274
rect -8726 144274 -8106 164038
rect -8726 144038 -8694 144274
rect -8458 144038 -8374 144274
rect -8138 144038 -8106 144274
rect -8726 124274 -8106 144038
rect -8726 124038 -8694 124274
rect -8458 124038 -8374 124274
rect -8138 124038 -8106 124274
rect -8726 104274 -8106 124038
rect -8726 104038 -8694 104274
rect -8458 104038 -8374 104274
rect -8138 104038 -8106 104274
rect -8726 84274 -8106 104038
rect -8726 84038 -8694 84274
rect -8458 84038 -8374 84274
rect -8138 84038 -8106 84274
rect -8726 64274 -8106 84038
rect -8726 64038 -8694 64274
rect -8458 64038 -8374 64274
rect -8138 64038 -8106 64274
rect -8726 44274 -8106 64038
rect -8726 44038 -8694 44274
rect -8458 44038 -8374 44274
rect -8138 44038 -8106 44274
rect -8726 24274 -8106 44038
rect -8726 24038 -8694 24274
rect -8458 24038 -8374 24274
rect -8138 24038 -8106 24274
rect -8726 -7066 -8106 24038
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 694274 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 694038 -7734 694274
rect -7498 694038 -7414 694274
rect -7178 694038 -7146 694274
rect -7766 674274 -7146 694038
rect -7766 674038 -7734 674274
rect -7498 674038 -7414 674274
rect -7178 674038 -7146 674274
rect -7766 654274 -7146 674038
rect -7766 654038 -7734 654274
rect -7498 654038 -7414 654274
rect -7178 654038 -7146 654274
rect -7766 634274 -7146 654038
rect -7766 634038 -7734 634274
rect -7498 634038 -7414 634274
rect -7178 634038 -7146 634274
rect -7766 614274 -7146 634038
rect -7766 614038 -7734 614274
rect -7498 614038 -7414 614274
rect -7178 614038 -7146 614274
rect -7766 594274 -7146 614038
rect -7766 594038 -7734 594274
rect -7498 594038 -7414 594274
rect -7178 594038 -7146 594274
rect -7766 574274 -7146 594038
rect -7766 574038 -7734 574274
rect -7498 574038 -7414 574274
rect -7178 574038 -7146 574274
rect -7766 554274 -7146 574038
rect -7766 554038 -7734 554274
rect -7498 554038 -7414 554274
rect -7178 554038 -7146 554274
rect -7766 534274 -7146 554038
rect -7766 534038 -7734 534274
rect -7498 534038 -7414 534274
rect -7178 534038 -7146 534274
rect -7766 514274 -7146 534038
rect -7766 514038 -7734 514274
rect -7498 514038 -7414 514274
rect -7178 514038 -7146 514274
rect -7766 494274 -7146 514038
rect -7766 494038 -7734 494274
rect -7498 494038 -7414 494274
rect -7178 494038 -7146 494274
rect -7766 474274 -7146 494038
rect -7766 474038 -7734 474274
rect -7498 474038 -7414 474274
rect -7178 474038 -7146 474274
rect -7766 454274 -7146 474038
rect -7766 454038 -7734 454274
rect -7498 454038 -7414 454274
rect -7178 454038 -7146 454274
rect -7766 434274 -7146 454038
rect -7766 434038 -7734 434274
rect -7498 434038 -7414 434274
rect -7178 434038 -7146 434274
rect -7766 414274 -7146 434038
rect -7766 414038 -7734 414274
rect -7498 414038 -7414 414274
rect -7178 414038 -7146 414274
rect -7766 394274 -7146 414038
rect -7766 394038 -7734 394274
rect -7498 394038 -7414 394274
rect -7178 394038 -7146 394274
rect -7766 374274 -7146 394038
rect -7766 374038 -7734 374274
rect -7498 374038 -7414 374274
rect -7178 374038 -7146 374274
rect -7766 354274 -7146 374038
rect -7766 354038 -7734 354274
rect -7498 354038 -7414 354274
rect -7178 354038 -7146 354274
rect -7766 334274 -7146 354038
rect -7766 334038 -7734 334274
rect -7498 334038 -7414 334274
rect -7178 334038 -7146 334274
rect -7766 314274 -7146 334038
rect -7766 314038 -7734 314274
rect -7498 314038 -7414 314274
rect -7178 314038 -7146 314274
rect -7766 294274 -7146 314038
rect -7766 294038 -7734 294274
rect -7498 294038 -7414 294274
rect -7178 294038 -7146 294274
rect -7766 274274 -7146 294038
rect -7766 274038 -7734 274274
rect -7498 274038 -7414 274274
rect -7178 274038 -7146 274274
rect -7766 254274 -7146 274038
rect -7766 254038 -7734 254274
rect -7498 254038 -7414 254274
rect -7178 254038 -7146 254274
rect -7766 234274 -7146 254038
rect -7766 234038 -7734 234274
rect -7498 234038 -7414 234274
rect -7178 234038 -7146 234274
rect -7766 214274 -7146 234038
rect -7766 214038 -7734 214274
rect -7498 214038 -7414 214274
rect -7178 214038 -7146 214274
rect -7766 194274 -7146 214038
rect -7766 194038 -7734 194274
rect -7498 194038 -7414 194274
rect -7178 194038 -7146 194274
rect -7766 174274 -7146 194038
rect -7766 174038 -7734 174274
rect -7498 174038 -7414 174274
rect -7178 174038 -7146 174274
rect -7766 154274 -7146 174038
rect -7766 154038 -7734 154274
rect -7498 154038 -7414 154274
rect -7178 154038 -7146 154274
rect -7766 134274 -7146 154038
rect -7766 134038 -7734 134274
rect -7498 134038 -7414 134274
rect -7178 134038 -7146 134274
rect -7766 114274 -7146 134038
rect -7766 114038 -7734 114274
rect -7498 114038 -7414 114274
rect -7178 114038 -7146 114274
rect -7766 94274 -7146 114038
rect -7766 94038 -7734 94274
rect -7498 94038 -7414 94274
rect -7178 94038 -7146 94274
rect -7766 74274 -7146 94038
rect -7766 74038 -7734 74274
rect -7498 74038 -7414 74274
rect -7178 74038 -7146 74274
rect -7766 54274 -7146 74038
rect -7766 54038 -7734 54274
rect -7498 54038 -7414 54274
rect -7178 54038 -7146 54274
rect -7766 34274 -7146 54038
rect -7766 34038 -7734 34274
rect -7498 34038 -7414 34274
rect -7178 34038 -7146 34274
rect -7766 14274 -7146 34038
rect -7766 14038 -7734 14274
rect -7498 14038 -7414 14274
rect -7178 14038 -7146 14274
rect -7766 -6106 -7146 14038
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 700614 -6186 709082
rect -6806 700378 -6774 700614
rect -6538 700378 -6454 700614
rect -6218 700378 -6186 700614
rect -6806 680614 -6186 700378
rect -6806 680378 -6774 680614
rect -6538 680378 -6454 680614
rect -6218 680378 -6186 680614
rect -6806 660614 -6186 680378
rect -6806 660378 -6774 660614
rect -6538 660378 -6454 660614
rect -6218 660378 -6186 660614
rect -6806 640614 -6186 660378
rect -6806 640378 -6774 640614
rect -6538 640378 -6454 640614
rect -6218 640378 -6186 640614
rect -6806 620614 -6186 640378
rect -6806 620378 -6774 620614
rect -6538 620378 -6454 620614
rect -6218 620378 -6186 620614
rect -6806 600614 -6186 620378
rect -6806 600378 -6774 600614
rect -6538 600378 -6454 600614
rect -6218 600378 -6186 600614
rect -6806 580614 -6186 600378
rect -6806 580378 -6774 580614
rect -6538 580378 -6454 580614
rect -6218 580378 -6186 580614
rect -6806 560614 -6186 580378
rect -6806 560378 -6774 560614
rect -6538 560378 -6454 560614
rect -6218 560378 -6186 560614
rect -6806 540614 -6186 560378
rect -6806 540378 -6774 540614
rect -6538 540378 -6454 540614
rect -6218 540378 -6186 540614
rect -6806 520614 -6186 540378
rect -6806 520378 -6774 520614
rect -6538 520378 -6454 520614
rect -6218 520378 -6186 520614
rect -6806 500614 -6186 520378
rect -6806 500378 -6774 500614
rect -6538 500378 -6454 500614
rect -6218 500378 -6186 500614
rect -6806 480614 -6186 500378
rect -6806 480378 -6774 480614
rect -6538 480378 -6454 480614
rect -6218 480378 -6186 480614
rect -6806 460614 -6186 480378
rect -6806 460378 -6774 460614
rect -6538 460378 -6454 460614
rect -6218 460378 -6186 460614
rect -6806 440614 -6186 460378
rect -6806 440378 -6774 440614
rect -6538 440378 -6454 440614
rect -6218 440378 -6186 440614
rect -6806 420614 -6186 440378
rect -6806 420378 -6774 420614
rect -6538 420378 -6454 420614
rect -6218 420378 -6186 420614
rect -6806 400614 -6186 420378
rect -6806 400378 -6774 400614
rect -6538 400378 -6454 400614
rect -6218 400378 -6186 400614
rect -6806 380614 -6186 400378
rect -6806 380378 -6774 380614
rect -6538 380378 -6454 380614
rect -6218 380378 -6186 380614
rect -6806 360614 -6186 380378
rect -6806 360378 -6774 360614
rect -6538 360378 -6454 360614
rect -6218 360378 -6186 360614
rect -6806 340614 -6186 360378
rect -6806 340378 -6774 340614
rect -6538 340378 -6454 340614
rect -6218 340378 -6186 340614
rect -6806 320614 -6186 340378
rect -6806 320378 -6774 320614
rect -6538 320378 -6454 320614
rect -6218 320378 -6186 320614
rect -6806 300614 -6186 320378
rect -6806 300378 -6774 300614
rect -6538 300378 -6454 300614
rect -6218 300378 -6186 300614
rect -6806 280614 -6186 300378
rect -6806 280378 -6774 280614
rect -6538 280378 -6454 280614
rect -6218 280378 -6186 280614
rect -6806 260614 -6186 280378
rect -6806 260378 -6774 260614
rect -6538 260378 -6454 260614
rect -6218 260378 -6186 260614
rect -6806 240614 -6186 260378
rect -6806 240378 -6774 240614
rect -6538 240378 -6454 240614
rect -6218 240378 -6186 240614
rect -6806 220614 -6186 240378
rect -6806 220378 -6774 220614
rect -6538 220378 -6454 220614
rect -6218 220378 -6186 220614
rect -6806 200614 -6186 220378
rect -6806 200378 -6774 200614
rect -6538 200378 -6454 200614
rect -6218 200378 -6186 200614
rect -6806 180614 -6186 200378
rect -6806 180378 -6774 180614
rect -6538 180378 -6454 180614
rect -6218 180378 -6186 180614
rect -6806 160614 -6186 180378
rect -6806 160378 -6774 160614
rect -6538 160378 -6454 160614
rect -6218 160378 -6186 160614
rect -6806 140614 -6186 160378
rect -6806 140378 -6774 140614
rect -6538 140378 -6454 140614
rect -6218 140378 -6186 140614
rect -6806 120614 -6186 140378
rect -6806 120378 -6774 120614
rect -6538 120378 -6454 120614
rect -6218 120378 -6186 120614
rect -6806 100614 -6186 120378
rect -6806 100378 -6774 100614
rect -6538 100378 -6454 100614
rect -6218 100378 -6186 100614
rect -6806 80614 -6186 100378
rect -6806 80378 -6774 80614
rect -6538 80378 -6454 80614
rect -6218 80378 -6186 80614
rect -6806 60614 -6186 80378
rect -6806 60378 -6774 60614
rect -6538 60378 -6454 60614
rect -6218 60378 -6186 60614
rect -6806 40614 -6186 60378
rect -6806 40378 -6774 40614
rect -6538 40378 -6454 40614
rect -6218 40378 -6186 40614
rect -6806 20614 -6186 40378
rect -6806 20378 -6774 20614
rect -6538 20378 -6454 20614
rect -6218 20378 -6186 20614
rect -6806 -5146 -6186 20378
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 690614 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 690378 -5814 690614
rect -5578 690378 -5494 690614
rect -5258 690378 -5226 690614
rect -5846 670614 -5226 690378
rect -5846 670378 -5814 670614
rect -5578 670378 -5494 670614
rect -5258 670378 -5226 670614
rect -5846 650614 -5226 670378
rect -5846 650378 -5814 650614
rect -5578 650378 -5494 650614
rect -5258 650378 -5226 650614
rect -5846 630614 -5226 650378
rect -5846 630378 -5814 630614
rect -5578 630378 -5494 630614
rect -5258 630378 -5226 630614
rect -5846 610614 -5226 630378
rect -5846 610378 -5814 610614
rect -5578 610378 -5494 610614
rect -5258 610378 -5226 610614
rect -5846 590614 -5226 610378
rect -5846 590378 -5814 590614
rect -5578 590378 -5494 590614
rect -5258 590378 -5226 590614
rect -5846 570614 -5226 590378
rect -5846 570378 -5814 570614
rect -5578 570378 -5494 570614
rect -5258 570378 -5226 570614
rect -5846 550614 -5226 570378
rect -5846 550378 -5814 550614
rect -5578 550378 -5494 550614
rect -5258 550378 -5226 550614
rect -5846 530614 -5226 550378
rect -5846 530378 -5814 530614
rect -5578 530378 -5494 530614
rect -5258 530378 -5226 530614
rect -5846 510614 -5226 530378
rect -5846 510378 -5814 510614
rect -5578 510378 -5494 510614
rect -5258 510378 -5226 510614
rect -5846 490614 -5226 510378
rect -5846 490378 -5814 490614
rect -5578 490378 -5494 490614
rect -5258 490378 -5226 490614
rect -5846 470614 -5226 490378
rect -5846 470378 -5814 470614
rect -5578 470378 -5494 470614
rect -5258 470378 -5226 470614
rect -5846 450614 -5226 470378
rect -5846 450378 -5814 450614
rect -5578 450378 -5494 450614
rect -5258 450378 -5226 450614
rect -5846 430614 -5226 450378
rect -5846 430378 -5814 430614
rect -5578 430378 -5494 430614
rect -5258 430378 -5226 430614
rect -5846 410614 -5226 430378
rect -5846 410378 -5814 410614
rect -5578 410378 -5494 410614
rect -5258 410378 -5226 410614
rect -5846 390614 -5226 410378
rect -5846 390378 -5814 390614
rect -5578 390378 -5494 390614
rect -5258 390378 -5226 390614
rect -5846 370614 -5226 390378
rect -5846 370378 -5814 370614
rect -5578 370378 -5494 370614
rect -5258 370378 -5226 370614
rect -5846 350614 -5226 370378
rect -5846 350378 -5814 350614
rect -5578 350378 -5494 350614
rect -5258 350378 -5226 350614
rect -5846 330614 -5226 350378
rect -5846 330378 -5814 330614
rect -5578 330378 -5494 330614
rect -5258 330378 -5226 330614
rect -5846 310614 -5226 330378
rect -5846 310378 -5814 310614
rect -5578 310378 -5494 310614
rect -5258 310378 -5226 310614
rect -5846 290614 -5226 310378
rect -5846 290378 -5814 290614
rect -5578 290378 -5494 290614
rect -5258 290378 -5226 290614
rect -5846 270614 -5226 290378
rect -5846 270378 -5814 270614
rect -5578 270378 -5494 270614
rect -5258 270378 -5226 270614
rect -5846 250614 -5226 270378
rect -5846 250378 -5814 250614
rect -5578 250378 -5494 250614
rect -5258 250378 -5226 250614
rect -5846 230614 -5226 250378
rect -5846 230378 -5814 230614
rect -5578 230378 -5494 230614
rect -5258 230378 -5226 230614
rect -5846 210614 -5226 230378
rect -5846 210378 -5814 210614
rect -5578 210378 -5494 210614
rect -5258 210378 -5226 210614
rect -5846 190614 -5226 210378
rect -5846 190378 -5814 190614
rect -5578 190378 -5494 190614
rect -5258 190378 -5226 190614
rect -5846 170614 -5226 190378
rect -5846 170378 -5814 170614
rect -5578 170378 -5494 170614
rect -5258 170378 -5226 170614
rect -5846 150614 -5226 170378
rect -5846 150378 -5814 150614
rect -5578 150378 -5494 150614
rect -5258 150378 -5226 150614
rect -5846 130614 -5226 150378
rect -5846 130378 -5814 130614
rect -5578 130378 -5494 130614
rect -5258 130378 -5226 130614
rect -5846 110614 -5226 130378
rect -5846 110378 -5814 110614
rect -5578 110378 -5494 110614
rect -5258 110378 -5226 110614
rect -5846 90614 -5226 110378
rect -5846 90378 -5814 90614
rect -5578 90378 -5494 90614
rect -5258 90378 -5226 90614
rect -5846 70614 -5226 90378
rect -5846 70378 -5814 70614
rect -5578 70378 -5494 70614
rect -5258 70378 -5226 70614
rect -5846 50614 -5226 70378
rect -5846 50378 -5814 50614
rect -5578 50378 -5494 50614
rect -5258 50378 -5226 50614
rect -5846 30614 -5226 50378
rect -5846 30378 -5814 30614
rect -5578 30378 -5494 30614
rect -5258 30378 -5226 30614
rect -5846 10614 -5226 30378
rect -5846 10378 -5814 10614
rect -5578 10378 -5494 10614
rect -5258 10378 -5226 10614
rect -5846 -4186 -5226 10378
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 696954 -4266 707162
rect -4886 696718 -4854 696954
rect -4618 696718 -4534 696954
rect -4298 696718 -4266 696954
rect -4886 676954 -4266 696718
rect -4886 676718 -4854 676954
rect -4618 676718 -4534 676954
rect -4298 676718 -4266 676954
rect -4886 656954 -4266 676718
rect -4886 656718 -4854 656954
rect -4618 656718 -4534 656954
rect -4298 656718 -4266 656954
rect -4886 636954 -4266 656718
rect -4886 636718 -4854 636954
rect -4618 636718 -4534 636954
rect -4298 636718 -4266 636954
rect -4886 616954 -4266 636718
rect -4886 616718 -4854 616954
rect -4618 616718 -4534 616954
rect -4298 616718 -4266 616954
rect -4886 596954 -4266 616718
rect -4886 596718 -4854 596954
rect -4618 596718 -4534 596954
rect -4298 596718 -4266 596954
rect -4886 576954 -4266 596718
rect -4886 576718 -4854 576954
rect -4618 576718 -4534 576954
rect -4298 576718 -4266 576954
rect -4886 556954 -4266 576718
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 536954 -4266 556718
rect -4886 536718 -4854 536954
rect -4618 536718 -4534 536954
rect -4298 536718 -4266 536954
rect -4886 516954 -4266 536718
rect -4886 516718 -4854 516954
rect -4618 516718 -4534 516954
rect -4298 516718 -4266 516954
rect -4886 496954 -4266 516718
rect -4886 496718 -4854 496954
rect -4618 496718 -4534 496954
rect -4298 496718 -4266 496954
rect -4886 476954 -4266 496718
rect -4886 476718 -4854 476954
rect -4618 476718 -4534 476954
rect -4298 476718 -4266 476954
rect -4886 456954 -4266 476718
rect -4886 456718 -4854 456954
rect -4618 456718 -4534 456954
rect -4298 456718 -4266 456954
rect -4886 436954 -4266 456718
rect -4886 436718 -4854 436954
rect -4618 436718 -4534 436954
rect -4298 436718 -4266 436954
rect -4886 416954 -4266 436718
rect -4886 416718 -4854 416954
rect -4618 416718 -4534 416954
rect -4298 416718 -4266 416954
rect -4886 396954 -4266 416718
rect -4886 396718 -4854 396954
rect -4618 396718 -4534 396954
rect -4298 396718 -4266 396954
rect -4886 376954 -4266 396718
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 356954 -4266 376718
rect -4886 356718 -4854 356954
rect -4618 356718 -4534 356954
rect -4298 356718 -4266 356954
rect -4886 336954 -4266 356718
rect -4886 336718 -4854 336954
rect -4618 336718 -4534 336954
rect -4298 336718 -4266 336954
rect -4886 316954 -4266 336718
rect -4886 316718 -4854 316954
rect -4618 316718 -4534 316954
rect -4298 316718 -4266 316954
rect -4886 296954 -4266 316718
rect -4886 296718 -4854 296954
rect -4618 296718 -4534 296954
rect -4298 296718 -4266 296954
rect -4886 276954 -4266 296718
rect -4886 276718 -4854 276954
rect -4618 276718 -4534 276954
rect -4298 276718 -4266 276954
rect -4886 256954 -4266 276718
rect -4886 256718 -4854 256954
rect -4618 256718 -4534 256954
rect -4298 256718 -4266 256954
rect -4886 236954 -4266 256718
rect -4886 236718 -4854 236954
rect -4618 236718 -4534 236954
rect -4298 236718 -4266 236954
rect -4886 216954 -4266 236718
rect -4886 216718 -4854 216954
rect -4618 216718 -4534 216954
rect -4298 216718 -4266 216954
rect -4886 196954 -4266 216718
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 176954 -4266 196718
rect -4886 176718 -4854 176954
rect -4618 176718 -4534 176954
rect -4298 176718 -4266 176954
rect -4886 156954 -4266 176718
rect -4886 156718 -4854 156954
rect -4618 156718 -4534 156954
rect -4298 156718 -4266 156954
rect -4886 136954 -4266 156718
rect -4886 136718 -4854 136954
rect -4618 136718 -4534 136954
rect -4298 136718 -4266 136954
rect -4886 116954 -4266 136718
rect -4886 116718 -4854 116954
rect -4618 116718 -4534 116954
rect -4298 116718 -4266 116954
rect -4886 96954 -4266 116718
rect -4886 96718 -4854 96954
rect -4618 96718 -4534 96954
rect -4298 96718 -4266 96954
rect -4886 76954 -4266 96718
rect -4886 76718 -4854 76954
rect -4618 76718 -4534 76954
rect -4298 76718 -4266 76954
rect -4886 56954 -4266 76718
rect -4886 56718 -4854 56954
rect -4618 56718 -4534 56954
rect -4298 56718 -4266 56954
rect -4886 36954 -4266 56718
rect -4886 36718 -4854 36954
rect -4618 36718 -4534 36954
rect -4298 36718 -4266 36954
rect -4886 16954 -4266 36718
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 -3226 -4266 16718
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 686954 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 686718 -3894 686954
rect -3658 686718 -3574 686954
rect -3338 686718 -3306 686954
rect -3926 666954 -3306 686718
rect -3926 666718 -3894 666954
rect -3658 666718 -3574 666954
rect -3338 666718 -3306 666954
rect -3926 646954 -3306 666718
rect -3926 646718 -3894 646954
rect -3658 646718 -3574 646954
rect -3338 646718 -3306 646954
rect -3926 626954 -3306 646718
rect -3926 626718 -3894 626954
rect -3658 626718 -3574 626954
rect -3338 626718 -3306 626954
rect -3926 606954 -3306 626718
rect -3926 606718 -3894 606954
rect -3658 606718 -3574 606954
rect -3338 606718 -3306 606954
rect -3926 586954 -3306 606718
rect -3926 586718 -3894 586954
rect -3658 586718 -3574 586954
rect -3338 586718 -3306 586954
rect -3926 566954 -3306 586718
rect -3926 566718 -3894 566954
rect -3658 566718 -3574 566954
rect -3338 566718 -3306 566954
rect -3926 546954 -3306 566718
rect -3926 546718 -3894 546954
rect -3658 546718 -3574 546954
rect -3338 546718 -3306 546954
rect -3926 526954 -3306 546718
rect -3926 526718 -3894 526954
rect -3658 526718 -3574 526954
rect -3338 526718 -3306 526954
rect -3926 506954 -3306 526718
rect -3926 506718 -3894 506954
rect -3658 506718 -3574 506954
rect -3338 506718 -3306 506954
rect -3926 486954 -3306 506718
rect -3926 486718 -3894 486954
rect -3658 486718 -3574 486954
rect -3338 486718 -3306 486954
rect -3926 466954 -3306 486718
rect -3926 466718 -3894 466954
rect -3658 466718 -3574 466954
rect -3338 466718 -3306 466954
rect -3926 446954 -3306 466718
rect -3926 446718 -3894 446954
rect -3658 446718 -3574 446954
rect -3338 446718 -3306 446954
rect -3926 426954 -3306 446718
rect -3926 426718 -3894 426954
rect -3658 426718 -3574 426954
rect -3338 426718 -3306 426954
rect -3926 406954 -3306 426718
rect -3926 406718 -3894 406954
rect -3658 406718 -3574 406954
rect -3338 406718 -3306 406954
rect -3926 386954 -3306 406718
rect -3926 386718 -3894 386954
rect -3658 386718 -3574 386954
rect -3338 386718 -3306 386954
rect -3926 366954 -3306 386718
rect -3926 366718 -3894 366954
rect -3658 366718 -3574 366954
rect -3338 366718 -3306 366954
rect -3926 346954 -3306 366718
rect -3926 346718 -3894 346954
rect -3658 346718 -3574 346954
rect -3338 346718 -3306 346954
rect -3926 326954 -3306 346718
rect -3926 326718 -3894 326954
rect -3658 326718 -3574 326954
rect -3338 326718 -3306 326954
rect -3926 306954 -3306 326718
rect -3926 306718 -3894 306954
rect -3658 306718 -3574 306954
rect -3338 306718 -3306 306954
rect -3926 286954 -3306 306718
rect -3926 286718 -3894 286954
rect -3658 286718 -3574 286954
rect -3338 286718 -3306 286954
rect -3926 266954 -3306 286718
rect -3926 266718 -3894 266954
rect -3658 266718 -3574 266954
rect -3338 266718 -3306 266954
rect -3926 246954 -3306 266718
rect -3926 246718 -3894 246954
rect -3658 246718 -3574 246954
rect -3338 246718 -3306 246954
rect -3926 226954 -3306 246718
rect -3926 226718 -3894 226954
rect -3658 226718 -3574 226954
rect -3338 226718 -3306 226954
rect -3926 206954 -3306 226718
rect -3926 206718 -3894 206954
rect -3658 206718 -3574 206954
rect -3338 206718 -3306 206954
rect -3926 186954 -3306 206718
rect -3926 186718 -3894 186954
rect -3658 186718 -3574 186954
rect -3338 186718 -3306 186954
rect -3926 166954 -3306 186718
rect -3926 166718 -3894 166954
rect -3658 166718 -3574 166954
rect -3338 166718 -3306 166954
rect -3926 146954 -3306 166718
rect -3926 146718 -3894 146954
rect -3658 146718 -3574 146954
rect -3338 146718 -3306 146954
rect -3926 126954 -3306 146718
rect -3926 126718 -3894 126954
rect -3658 126718 -3574 126954
rect -3338 126718 -3306 126954
rect -3926 106954 -3306 126718
rect -3926 106718 -3894 106954
rect -3658 106718 -3574 106954
rect -3338 106718 -3306 106954
rect -3926 86954 -3306 106718
rect -3926 86718 -3894 86954
rect -3658 86718 -3574 86954
rect -3338 86718 -3306 86954
rect -3926 66954 -3306 86718
rect -3926 66718 -3894 66954
rect -3658 66718 -3574 66954
rect -3338 66718 -3306 66954
rect -3926 46954 -3306 66718
rect -3926 46718 -3894 46954
rect -3658 46718 -3574 46954
rect -3338 46718 -3306 46954
rect -3926 26954 -3306 46718
rect -3926 26718 -3894 26954
rect -3658 26718 -3574 26954
rect -3338 26718 -3306 26954
rect -3926 6954 -3306 26718
rect -3926 6718 -3894 6954
rect -3658 6718 -3574 6954
rect -3338 6718 -3306 6954
rect -3926 -2266 -3306 6718
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 693294 -2346 705242
rect -2966 693058 -2934 693294
rect -2698 693058 -2614 693294
rect -2378 693058 -2346 693294
rect -2966 673294 -2346 693058
rect -2966 673058 -2934 673294
rect -2698 673058 -2614 673294
rect -2378 673058 -2346 673294
rect -2966 653294 -2346 673058
rect -2966 653058 -2934 653294
rect -2698 653058 -2614 653294
rect -2378 653058 -2346 653294
rect -2966 633294 -2346 653058
rect -2966 633058 -2934 633294
rect -2698 633058 -2614 633294
rect -2378 633058 -2346 633294
rect -2966 613294 -2346 633058
rect -2966 613058 -2934 613294
rect -2698 613058 -2614 613294
rect -2378 613058 -2346 613294
rect -2966 593294 -2346 613058
rect -2966 593058 -2934 593294
rect -2698 593058 -2614 593294
rect -2378 593058 -2346 593294
rect -2966 573294 -2346 593058
rect -2966 573058 -2934 573294
rect -2698 573058 -2614 573294
rect -2378 573058 -2346 573294
rect -2966 553294 -2346 573058
rect -2966 553058 -2934 553294
rect -2698 553058 -2614 553294
rect -2378 553058 -2346 553294
rect -2966 533294 -2346 553058
rect -2966 533058 -2934 533294
rect -2698 533058 -2614 533294
rect -2378 533058 -2346 533294
rect -2966 513294 -2346 533058
rect -2966 513058 -2934 513294
rect -2698 513058 -2614 513294
rect -2378 513058 -2346 513294
rect -2966 493294 -2346 513058
rect -2966 493058 -2934 493294
rect -2698 493058 -2614 493294
rect -2378 493058 -2346 493294
rect -2966 473294 -2346 493058
rect -2966 473058 -2934 473294
rect -2698 473058 -2614 473294
rect -2378 473058 -2346 473294
rect -2966 453294 -2346 473058
rect -2966 453058 -2934 453294
rect -2698 453058 -2614 453294
rect -2378 453058 -2346 453294
rect -2966 433294 -2346 453058
rect -2966 433058 -2934 433294
rect -2698 433058 -2614 433294
rect -2378 433058 -2346 433294
rect -2966 413294 -2346 433058
rect -2966 413058 -2934 413294
rect -2698 413058 -2614 413294
rect -2378 413058 -2346 413294
rect -2966 393294 -2346 413058
rect -2966 393058 -2934 393294
rect -2698 393058 -2614 393294
rect -2378 393058 -2346 393294
rect -2966 373294 -2346 393058
rect -2966 373058 -2934 373294
rect -2698 373058 -2614 373294
rect -2378 373058 -2346 373294
rect -2966 353294 -2346 373058
rect -2966 353058 -2934 353294
rect -2698 353058 -2614 353294
rect -2378 353058 -2346 353294
rect -2966 333294 -2346 353058
rect -2966 333058 -2934 333294
rect -2698 333058 -2614 333294
rect -2378 333058 -2346 333294
rect -2966 313294 -2346 333058
rect -2966 313058 -2934 313294
rect -2698 313058 -2614 313294
rect -2378 313058 -2346 313294
rect -2966 293294 -2346 313058
rect -2966 293058 -2934 293294
rect -2698 293058 -2614 293294
rect -2378 293058 -2346 293294
rect -2966 273294 -2346 293058
rect -2966 273058 -2934 273294
rect -2698 273058 -2614 273294
rect -2378 273058 -2346 273294
rect -2966 253294 -2346 273058
rect -2966 253058 -2934 253294
rect -2698 253058 -2614 253294
rect -2378 253058 -2346 253294
rect -2966 233294 -2346 253058
rect -2966 233058 -2934 233294
rect -2698 233058 -2614 233294
rect -2378 233058 -2346 233294
rect -2966 213294 -2346 233058
rect -2966 213058 -2934 213294
rect -2698 213058 -2614 213294
rect -2378 213058 -2346 213294
rect -2966 193294 -2346 213058
rect -2966 193058 -2934 193294
rect -2698 193058 -2614 193294
rect -2378 193058 -2346 193294
rect -2966 173294 -2346 193058
rect -2966 173058 -2934 173294
rect -2698 173058 -2614 173294
rect -2378 173058 -2346 173294
rect -2966 153294 -2346 173058
rect -2966 153058 -2934 153294
rect -2698 153058 -2614 153294
rect -2378 153058 -2346 153294
rect -2966 133294 -2346 153058
rect -2966 133058 -2934 133294
rect -2698 133058 -2614 133294
rect -2378 133058 -2346 133294
rect -2966 113294 -2346 133058
rect -2966 113058 -2934 113294
rect -2698 113058 -2614 113294
rect -2378 113058 -2346 113294
rect -2966 93294 -2346 113058
rect -2966 93058 -2934 93294
rect -2698 93058 -2614 93294
rect -2378 93058 -2346 93294
rect -2966 73294 -2346 93058
rect -2966 73058 -2934 73294
rect -2698 73058 -2614 73294
rect -2378 73058 -2346 73294
rect -2966 53294 -2346 73058
rect -2966 53058 -2934 53294
rect -2698 53058 -2614 53294
rect -2378 53058 -2346 53294
rect -2966 33294 -2346 53058
rect -2966 33058 -2934 33294
rect -2698 33058 -2614 33294
rect -2378 33058 -2346 33294
rect -2966 13294 -2346 33058
rect -2966 13058 -2934 13294
rect -2698 13058 -2614 13294
rect -2378 13058 -2346 13294
rect -2966 -1306 -2346 13058
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 683294 -1386 704282
rect -2006 683058 -1974 683294
rect -1738 683058 -1654 683294
rect -1418 683058 -1386 683294
rect -2006 663294 -1386 683058
rect -2006 663058 -1974 663294
rect -1738 663058 -1654 663294
rect -1418 663058 -1386 663294
rect -2006 643294 -1386 663058
rect -2006 643058 -1974 643294
rect -1738 643058 -1654 643294
rect -1418 643058 -1386 643294
rect -2006 623294 -1386 643058
rect -2006 623058 -1974 623294
rect -1738 623058 -1654 623294
rect -1418 623058 -1386 623294
rect -2006 603294 -1386 623058
rect -2006 603058 -1974 603294
rect -1738 603058 -1654 603294
rect -1418 603058 -1386 603294
rect -2006 583294 -1386 603058
rect -2006 583058 -1974 583294
rect -1738 583058 -1654 583294
rect -1418 583058 -1386 583294
rect -2006 563294 -1386 583058
rect -2006 563058 -1974 563294
rect -1738 563058 -1654 563294
rect -1418 563058 -1386 563294
rect -2006 543294 -1386 563058
rect -2006 543058 -1974 543294
rect -1738 543058 -1654 543294
rect -1418 543058 -1386 543294
rect -2006 523294 -1386 543058
rect -2006 523058 -1974 523294
rect -1738 523058 -1654 523294
rect -1418 523058 -1386 523294
rect -2006 503294 -1386 523058
rect -2006 503058 -1974 503294
rect -1738 503058 -1654 503294
rect -1418 503058 -1386 503294
rect -2006 483294 -1386 503058
rect -2006 483058 -1974 483294
rect -1738 483058 -1654 483294
rect -1418 483058 -1386 483294
rect -2006 463294 -1386 483058
rect -2006 463058 -1974 463294
rect -1738 463058 -1654 463294
rect -1418 463058 -1386 463294
rect -2006 443294 -1386 463058
rect -2006 443058 -1974 443294
rect -1738 443058 -1654 443294
rect -1418 443058 -1386 443294
rect -2006 423294 -1386 443058
rect -2006 423058 -1974 423294
rect -1738 423058 -1654 423294
rect -1418 423058 -1386 423294
rect -2006 403294 -1386 423058
rect -2006 403058 -1974 403294
rect -1738 403058 -1654 403294
rect -1418 403058 -1386 403294
rect -2006 383294 -1386 403058
rect -2006 383058 -1974 383294
rect -1738 383058 -1654 383294
rect -1418 383058 -1386 383294
rect -2006 363294 -1386 383058
rect -2006 363058 -1974 363294
rect -1738 363058 -1654 363294
rect -1418 363058 -1386 363294
rect -2006 343294 -1386 363058
rect -2006 343058 -1974 343294
rect -1738 343058 -1654 343294
rect -1418 343058 -1386 343294
rect -2006 323294 -1386 343058
rect -2006 323058 -1974 323294
rect -1738 323058 -1654 323294
rect -1418 323058 -1386 323294
rect -2006 303294 -1386 323058
rect -2006 303058 -1974 303294
rect -1738 303058 -1654 303294
rect -1418 303058 -1386 303294
rect -2006 283294 -1386 303058
rect -2006 283058 -1974 283294
rect -1738 283058 -1654 283294
rect -1418 283058 -1386 283294
rect -2006 263294 -1386 283058
rect -2006 263058 -1974 263294
rect -1738 263058 -1654 263294
rect -1418 263058 -1386 263294
rect -2006 243294 -1386 263058
rect -2006 243058 -1974 243294
rect -1738 243058 -1654 243294
rect -1418 243058 -1386 243294
rect -2006 223294 -1386 243058
rect -2006 223058 -1974 223294
rect -1738 223058 -1654 223294
rect -1418 223058 -1386 223294
rect -2006 203294 -1386 223058
rect -2006 203058 -1974 203294
rect -1738 203058 -1654 203294
rect -1418 203058 -1386 203294
rect -2006 183294 -1386 203058
rect -2006 183058 -1974 183294
rect -1738 183058 -1654 183294
rect -1418 183058 -1386 183294
rect -2006 163294 -1386 183058
rect -2006 163058 -1974 163294
rect -1738 163058 -1654 163294
rect -1418 163058 -1386 163294
rect -2006 143294 -1386 163058
rect -2006 143058 -1974 143294
rect -1738 143058 -1654 143294
rect -1418 143058 -1386 143294
rect -2006 123294 -1386 143058
rect -2006 123058 -1974 123294
rect -1738 123058 -1654 123294
rect -1418 123058 -1386 123294
rect -2006 103294 -1386 123058
rect -2006 103058 -1974 103294
rect -1738 103058 -1654 103294
rect -1418 103058 -1386 103294
rect -2006 83294 -1386 103058
rect -2006 83058 -1974 83294
rect -1738 83058 -1654 83294
rect -1418 83058 -1386 83294
rect -2006 63294 -1386 83058
rect -2006 63058 -1974 63294
rect -1738 63058 -1654 63294
rect -1418 63058 -1386 63294
rect -2006 43294 -1386 63058
rect -2006 43058 -1974 43294
rect -1738 43058 -1654 43294
rect -1418 43058 -1386 43294
rect -2006 23294 -1386 43058
rect -2006 23058 -1974 23294
rect -1738 23058 -1654 23294
rect -1418 23058 -1386 23294
rect -2006 3294 -1386 23058
rect -2006 3058 -1974 3294
rect -1738 3058 -1654 3294
rect -1418 3058 -1386 3294
rect -2006 -346 -1386 3058
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 683294 2414 704282
rect 1794 683058 1826 683294
rect 2062 683058 2146 683294
rect 2382 683058 2414 683294
rect 1794 663294 2414 683058
rect 1794 663058 1826 663294
rect 2062 663058 2146 663294
rect 2382 663058 2414 663294
rect 1794 643294 2414 663058
rect 1794 643058 1826 643294
rect 2062 643058 2146 643294
rect 2382 643058 2414 643294
rect 1794 623294 2414 643058
rect 1794 623058 1826 623294
rect 2062 623058 2146 623294
rect 2382 623058 2414 623294
rect 1794 603294 2414 623058
rect 1794 603058 1826 603294
rect 2062 603058 2146 603294
rect 2382 603058 2414 603294
rect 1794 583294 2414 603058
rect 1794 583058 1826 583294
rect 2062 583058 2146 583294
rect 2382 583058 2414 583294
rect 1794 563294 2414 583058
rect 1794 563058 1826 563294
rect 2062 563058 2146 563294
rect 2382 563058 2414 563294
rect 1794 543294 2414 563058
rect 1794 543058 1826 543294
rect 2062 543058 2146 543294
rect 2382 543058 2414 543294
rect 1794 523294 2414 543058
rect 1794 523058 1826 523294
rect 2062 523058 2146 523294
rect 2382 523058 2414 523294
rect 1794 503294 2414 523058
rect 1794 503058 1826 503294
rect 2062 503058 2146 503294
rect 2382 503058 2414 503294
rect 1794 483294 2414 503058
rect 1794 483058 1826 483294
rect 2062 483058 2146 483294
rect 2382 483058 2414 483294
rect 1794 463294 2414 483058
rect 1794 463058 1826 463294
rect 2062 463058 2146 463294
rect 2382 463058 2414 463294
rect 1794 443294 2414 463058
rect 1794 443058 1826 443294
rect 2062 443058 2146 443294
rect 2382 443058 2414 443294
rect 1794 423294 2414 443058
rect 1794 423058 1826 423294
rect 2062 423058 2146 423294
rect 2382 423058 2414 423294
rect 1794 403294 2414 423058
rect 1794 403058 1826 403294
rect 2062 403058 2146 403294
rect 2382 403058 2414 403294
rect 1794 383294 2414 403058
rect 1794 383058 1826 383294
rect 2062 383058 2146 383294
rect 2382 383058 2414 383294
rect 1794 363294 2414 383058
rect 1794 363058 1826 363294
rect 2062 363058 2146 363294
rect 2382 363058 2414 363294
rect 1794 343294 2414 363058
rect 1794 343058 1826 343294
rect 2062 343058 2146 343294
rect 2382 343058 2414 343294
rect 1794 323294 2414 343058
rect 1794 323058 1826 323294
rect 2062 323058 2146 323294
rect 2382 323058 2414 323294
rect 1794 303294 2414 323058
rect 1794 303058 1826 303294
rect 2062 303058 2146 303294
rect 2382 303058 2414 303294
rect 1794 283294 2414 303058
rect 1794 283058 1826 283294
rect 2062 283058 2146 283294
rect 2382 283058 2414 283294
rect 1794 263294 2414 283058
rect 1794 263058 1826 263294
rect 2062 263058 2146 263294
rect 2382 263058 2414 263294
rect 1794 243294 2414 263058
rect 1794 243058 1826 243294
rect 2062 243058 2146 243294
rect 2382 243058 2414 243294
rect 1794 223294 2414 243058
rect 1794 223058 1826 223294
rect 2062 223058 2146 223294
rect 2382 223058 2414 223294
rect 1794 203294 2414 223058
rect 1794 203058 1826 203294
rect 2062 203058 2146 203294
rect 2382 203058 2414 203294
rect 1794 183294 2414 203058
rect 1794 183058 1826 183294
rect 2062 183058 2146 183294
rect 2382 183058 2414 183294
rect 1794 163294 2414 183058
rect 1794 163058 1826 163294
rect 2062 163058 2146 163294
rect 2382 163058 2414 163294
rect 1794 143294 2414 163058
rect 1794 143058 1826 143294
rect 2062 143058 2146 143294
rect 2382 143058 2414 143294
rect 1794 123294 2414 143058
rect 1794 123058 1826 123294
rect 2062 123058 2146 123294
rect 2382 123058 2414 123294
rect 1794 103294 2414 123058
rect 1794 103058 1826 103294
rect 2062 103058 2146 103294
rect 2382 103058 2414 103294
rect 1794 83294 2414 103058
rect 1794 83058 1826 83294
rect 2062 83058 2146 83294
rect 2382 83058 2414 83294
rect 1794 63294 2414 83058
rect 1794 63058 1826 63294
rect 2062 63058 2146 63294
rect 2382 63058 2414 63294
rect 1794 43294 2414 63058
rect 1794 43058 1826 43294
rect 2062 43058 2146 43294
rect 2382 43058 2414 43294
rect 1794 23294 2414 43058
rect 1794 23058 1826 23294
rect 2062 23058 2146 23294
rect 2382 23058 2414 23294
rect 1794 3294 2414 23058
rect 1794 3058 1826 3294
rect 2062 3058 2146 3294
rect 2382 3058 2414 3294
rect 1794 -346 2414 3058
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 686954 6134 706202
rect 5514 686718 5546 686954
rect 5782 686718 5866 686954
rect 6102 686718 6134 686954
rect 5514 666954 6134 686718
rect 5514 666718 5546 666954
rect 5782 666718 5866 666954
rect 6102 666718 6134 666954
rect 5514 646954 6134 666718
rect 5514 646718 5546 646954
rect 5782 646718 5866 646954
rect 6102 646718 6134 646954
rect 5514 626954 6134 646718
rect 5514 626718 5546 626954
rect 5782 626718 5866 626954
rect 6102 626718 6134 626954
rect 5514 606954 6134 626718
rect 5514 606718 5546 606954
rect 5782 606718 5866 606954
rect 6102 606718 6134 606954
rect 5514 586954 6134 606718
rect 5514 586718 5546 586954
rect 5782 586718 5866 586954
rect 6102 586718 6134 586954
rect 5514 566954 6134 586718
rect 5514 566718 5546 566954
rect 5782 566718 5866 566954
rect 6102 566718 6134 566954
rect 5514 546954 6134 566718
rect 5514 546718 5546 546954
rect 5782 546718 5866 546954
rect 6102 546718 6134 546954
rect 5514 526954 6134 546718
rect 5514 526718 5546 526954
rect 5782 526718 5866 526954
rect 6102 526718 6134 526954
rect 5514 506954 6134 526718
rect 5514 506718 5546 506954
rect 5782 506718 5866 506954
rect 6102 506718 6134 506954
rect 5514 486954 6134 506718
rect 5514 486718 5546 486954
rect 5782 486718 5866 486954
rect 6102 486718 6134 486954
rect 5514 466954 6134 486718
rect 5514 466718 5546 466954
rect 5782 466718 5866 466954
rect 6102 466718 6134 466954
rect 5514 446954 6134 466718
rect 5514 446718 5546 446954
rect 5782 446718 5866 446954
rect 6102 446718 6134 446954
rect 5514 426954 6134 446718
rect 5514 426718 5546 426954
rect 5782 426718 5866 426954
rect 6102 426718 6134 426954
rect 5514 406954 6134 426718
rect 5514 406718 5546 406954
rect 5782 406718 5866 406954
rect 6102 406718 6134 406954
rect 5514 386954 6134 406718
rect 5514 386718 5546 386954
rect 5782 386718 5866 386954
rect 6102 386718 6134 386954
rect 5514 366954 6134 386718
rect 5514 366718 5546 366954
rect 5782 366718 5866 366954
rect 6102 366718 6134 366954
rect 5514 346954 6134 366718
rect 5514 346718 5546 346954
rect 5782 346718 5866 346954
rect 6102 346718 6134 346954
rect 5514 326954 6134 346718
rect 5514 326718 5546 326954
rect 5782 326718 5866 326954
rect 6102 326718 6134 326954
rect 5514 306954 6134 326718
rect 5514 306718 5546 306954
rect 5782 306718 5866 306954
rect 6102 306718 6134 306954
rect 5514 286954 6134 306718
rect 5514 286718 5546 286954
rect 5782 286718 5866 286954
rect 6102 286718 6134 286954
rect 5514 266954 6134 286718
rect 5514 266718 5546 266954
rect 5782 266718 5866 266954
rect 6102 266718 6134 266954
rect 5514 246954 6134 266718
rect 5514 246718 5546 246954
rect 5782 246718 5866 246954
rect 6102 246718 6134 246954
rect 5514 226954 6134 246718
rect 5514 226718 5546 226954
rect 5782 226718 5866 226954
rect 6102 226718 6134 226954
rect 5514 206954 6134 226718
rect 5514 206718 5546 206954
rect 5782 206718 5866 206954
rect 6102 206718 6134 206954
rect 5514 186954 6134 206718
rect 5514 186718 5546 186954
rect 5782 186718 5866 186954
rect 6102 186718 6134 186954
rect 5514 166954 6134 186718
rect 5514 166718 5546 166954
rect 5782 166718 5866 166954
rect 6102 166718 6134 166954
rect 5514 146954 6134 166718
rect 5514 146718 5546 146954
rect 5782 146718 5866 146954
rect 6102 146718 6134 146954
rect 5514 126954 6134 146718
rect 5514 126718 5546 126954
rect 5782 126718 5866 126954
rect 6102 126718 6134 126954
rect 5514 106954 6134 126718
rect 5514 106718 5546 106954
rect 5782 106718 5866 106954
rect 6102 106718 6134 106954
rect 5514 86954 6134 106718
rect 5514 86718 5546 86954
rect 5782 86718 5866 86954
rect 6102 86718 6134 86954
rect 5514 66954 6134 86718
rect 5514 66718 5546 66954
rect 5782 66718 5866 66954
rect 6102 66718 6134 66954
rect 5514 46954 6134 66718
rect 5514 46718 5546 46954
rect 5782 46718 5866 46954
rect 6102 46718 6134 46954
rect 5514 26954 6134 46718
rect 5514 26718 5546 26954
rect 5782 26718 5866 26954
rect 6102 26718 6134 26954
rect 5514 6954 6134 26718
rect 5514 6718 5546 6954
rect 5782 6718 5866 6954
rect 6102 6718 6134 6954
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6718
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 690614 9854 708122
rect 9234 690378 9266 690614
rect 9502 690378 9586 690614
rect 9822 690378 9854 690614
rect 9234 670614 9854 690378
rect 9234 670378 9266 670614
rect 9502 670378 9586 670614
rect 9822 670378 9854 670614
rect 9234 650614 9854 670378
rect 9234 650378 9266 650614
rect 9502 650378 9586 650614
rect 9822 650378 9854 650614
rect 9234 630614 9854 650378
rect 9234 630378 9266 630614
rect 9502 630378 9586 630614
rect 9822 630378 9854 630614
rect 9234 610614 9854 630378
rect 9234 610378 9266 610614
rect 9502 610378 9586 610614
rect 9822 610378 9854 610614
rect 9234 590614 9854 610378
rect 9234 590378 9266 590614
rect 9502 590378 9586 590614
rect 9822 590378 9854 590614
rect 9234 570614 9854 590378
rect 9234 570378 9266 570614
rect 9502 570378 9586 570614
rect 9822 570378 9854 570614
rect 9234 550614 9854 570378
rect 9234 550378 9266 550614
rect 9502 550378 9586 550614
rect 9822 550378 9854 550614
rect 9234 530614 9854 550378
rect 9234 530378 9266 530614
rect 9502 530378 9586 530614
rect 9822 530378 9854 530614
rect 9234 510614 9854 530378
rect 9234 510378 9266 510614
rect 9502 510378 9586 510614
rect 9822 510378 9854 510614
rect 9234 490614 9854 510378
rect 9234 490378 9266 490614
rect 9502 490378 9586 490614
rect 9822 490378 9854 490614
rect 9234 470614 9854 490378
rect 9234 470378 9266 470614
rect 9502 470378 9586 470614
rect 9822 470378 9854 470614
rect 9234 450614 9854 470378
rect 9234 450378 9266 450614
rect 9502 450378 9586 450614
rect 9822 450378 9854 450614
rect 9234 430614 9854 450378
rect 9234 430378 9266 430614
rect 9502 430378 9586 430614
rect 9822 430378 9854 430614
rect 9234 410614 9854 430378
rect 9234 410378 9266 410614
rect 9502 410378 9586 410614
rect 9822 410378 9854 410614
rect 9234 390614 9854 410378
rect 9234 390378 9266 390614
rect 9502 390378 9586 390614
rect 9822 390378 9854 390614
rect 9234 370614 9854 390378
rect 9234 370378 9266 370614
rect 9502 370378 9586 370614
rect 9822 370378 9854 370614
rect 9234 350614 9854 370378
rect 9234 350378 9266 350614
rect 9502 350378 9586 350614
rect 9822 350378 9854 350614
rect 9234 330614 9854 350378
rect 9234 330378 9266 330614
rect 9502 330378 9586 330614
rect 9822 330378 9854 330614
rect 9234 310614 9854 330378
rect 9234 310378 9266 310614
rect 9502 310378 9586 310614
rect 9822 310378 9854 310614
rect 9234 290614 9854 310378
rect 9234 290378 9266 290614
rect 9502 290378 9586 290614
rect 9822 290378 9854 290614
rect 9234 270614 9854 290378
rect 9234 270378 9266 270614
rect 9502 270378 9586 270614
rect 9822 270378 9854 270614
rect 9234 250614 9854 270378
rect 9234 250378 9266 250614
rect 9502 250378 9586 250614
rect 9822 250378 9854 250614
rect 9234 230614 9854 250378
rect 9234 230378 9266 230614
rect 9502 230378 9586 230614
rect 9822 230378 9854 230614
rect 9234 210614 9854 230378
rect 9234 210378 9266 210614
rect 9502 210378 9586 210614
rect 9822 210378 9854 210614
rect 9234 190614 9854 210378
rect 9234 190378 9266 190614
rect 9502 190378 9586 190614
rect 9822 190378 9854 190614
rect 9234 170614 9854 190378
rect 9234 170378 9266 170614
rect 9502 170378 9586 170614
rect 9822 170378 9854 170614
rect 9234 150614 9854 170378
rect 9234 150378 9266 150614
rect 9502 150378 9586 150614
rect 9822 150378 9854 150614
rect 9234 130614 9854 150378
rect 9234 130378 9266 130614
rect 9502 130378 9586 130614
rect 9822 130378 9854 130614
rect 9234 110614 9854 130378
rect 9234 110378 9266 110614
rect 9502 110378 9586 110614
rect 9822 110378 9854 110614
rect 9234 90614 9854 110378
rect 9234 90378 9266 90614
rect 9502 90378 9586 90614
rect 9822 90378 9854 90614
rect 9234 70614 9854 90378
rect 9234 70378 9266 70614
rect 9502 70378 9586 70614
rect 9822 70378 9854 70614
rect 9234 50614 9854 70378
rect 9234 50378 9266 50614
rect 9502 50378 9586 50614
rect 9822 50378 9854 50614
rect 9234 30614 9854 50378
rect 9234 30378 9266 30614
rect 9502 30378 9586 30614
rect 9822 30378 9854 30614
rect 9234 10614 9854 30378
rect 9234 10378 9266 10614
rect 9502 10378 9586 10614
rect 9822 10378 9854 10614
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10378
rect 11794 705798 12414 705830
rect 11794 705562 11826 705798
rect 12062 705562 12146 705798
rect 12382 705562 12414 705798
rect 11794 705478 12414 705562
rect 11794 705242 11826 705478
rect 12062 705242 12146 705478
rect 12382 705242 12414 705478
rect 11794 693294 12414 705242
rect 11794 693058 11826 693294
rect 12062 693058 12146 693294
rect 12382 693058 12414 693294
rect 11794 673294 12414 693058
rect 11794 673058 11826 673294
rect 12062 673058 12146 673294
rect 12382 673058 12414 673294
rect 11794 653294 12414 673058
rect 11794 653058 11826 653294
rect 12062 653058 12146 653294
rect 12382 653058 12414 653294
rect 11794 633294 12414 653058
rect 11794 633058 11826 633294
rect 12062 633058 12146 633294
rect 12382 633058 12414 633294
rect 11794 613294 12414 633058
rect 11794 613058 11826 613294
rect 12062 613058 12146 613294
rect 12382 613058 12414 613294
rect 11794 593294 12414 613058
rect 11794 593058 11826 593294
rect 12062 593058 12146 593294
rect 12382 593058 12414 593294
rect 11794 573294 12414 593058
rect 11794 573058 11826 573294
rect 12062 573058 12146 573294
rect 12382 573058 12414 573294
rect 11794 553294 12414 573058
rect 11794 553058 11826 553294
rect 12062 553058 12146 553294
rect 12382 553058 12414 553294
rect 11794 533294 12414 553058
rect 11794 533058 11826 533294
rect 12062 533058 12146 533294
rect 12382 533058 12414 533294
rect 11794 513294 12414 533058
rect 11794 513058 11826 513294
rect 12062 513058 12146 513294
rect 12382 513058 12414 513294
rect 11794 493294 12414 513058
rect 11794 493058 11826 493294
rect 12062 493058 12146 493294
rect 12382 493058 12414 493294
rect 11794 473294 12414 493058
rect 11794 473058 11826 473294
rect 12062 473058 12146 473294
rect 12382 473058 12414 473294
rect 11794 453294 12414 473058
rect 11794 453058 11826 453294
rect 12062 453058 12146 453294
rect 12382 453058 12414 453294
rect 11794 433294 12414 453058
rect 11794 433058 11826 433294
rect 12062 433058 12146 433294
rect 12382 433058 12414 433294
rect 11794 413294 12414 433058
rect 11794 413058 11826 413294
rect 12062 413058 12146 413294
rect 12382 413058 12414 413294
rect 11794 393294 12414 413058
rect 11794 393058 11826 393294
rect 12062 393058 12146 393294
rect 12382 393058 12414 393294
rect 11794 373294 12414 393058
rect 11794 373058 11826 373294
rect 12062 373058 12146 373294
rect 12382 373058 12414 373294
rect 11794 353294 12414 373058
rect 11794 353058 11826 353294
rect 12062 353058 12146 353294
rect 12382 353058 12414 353294
rect 11794 333294 12414 353058
rect 11794 333058 11826 333294
rect 12062 333058 12146 333294
rect 12382 333058 12414 333294
rect 11794 313294 12414 333058
rect 11794 313058 11826 313294
rect 12062 313058 12146 313294
rect 12382 313058 12414 313294
rect 11794 293294 12414 313058
rect 11794 293058 11826 293294
rect 12062 293058 12146 293294
rect 12382 293058 12414 293294
rect 11794 273294 12414 293058
rect 11794 273058 11826 273294
rect 12062 273058 12146 273294
rect 12382 273058 12414 273294
rect 11794 253294 12414 273058
rect 11794 253058 11826 253294
rect 12062 253058 12146 253294
rect 12382 253058 12414 253294
rect 11794 233294 12414 253058
rect 11794 233058 11826 233294
rect 12062 233058 12146 233294
rect 12382 233058 12414 233294
rect 11794 213294 12414 233058
rect 11794 213058 11826 213294
rect 12062 213058 12146 213294
rect 12382 213058 12414 213294
rect 11794 193294 12414 213058
rect 11794 193058 11826 193294
rect 12062 193058 12146 193294
rect 12382 193058 12414 193294
rect 11794 173294 12414 193058
rect 11794 173058 11826 173294
rect 12062 173058 12146 173294
rect 12382 173058 12414 173294
rect 11794 153294 12414 173058
rect 11794 153058 11826 153294
rect 12062 153058 12146 153294
rect 12382 153058 12414 153294
rect 11794 133294 12414 153058
rect 11794 133058 11826 133294
rect 12062 133058 12146 133294
rect 12382 133058 12414 133294
rect 11794 113294 12414 133058
rect 11794 113058 11826 113294
rect 12062 113058 12146 113294
rect 12382 113058 12414 113294
rect 11794 93294 12414 113058
rect 11794 93058 11826 93294
rect 12062 93058 12146 93294
rect 12382 93058 12414 93294
rect 11794 73294 12414 93058
rect 11794 73058 11826 73294
rect 12062 73058 12146 73294
rect 12382 73058 12414 73294
rect 11794 53294 12414 73058
rect 11794 53058 11826 53294
rect 12062 53058 12146 53294
rect 12382 53058 12414 53294
rect 11794 33294 12414 53058
rect 11794 33058 11826 33294
rect 12062 33058 12146 33294
rect 12382 33058 12414 33294
rect 11794 13294 12414 33058
rect 11794 13058 11826 13294
rect 12062 13058 12146 13294
rect 12382 13058 12414 13294
rect 11794 -1306 12414 13058
rect 11794 -1542 11826 -1306
rect 12062 -1542 12146 -1306
rect 12382 -1542 12414 -1306
rect 11794 -1626 12414 -1542
rect 11794 -1862 11826 -1626
rect 12062 -1862 12146 -1626
rect 12382 -1862 12414 -1626
rect 11794 -1894 12414 -1862
rect 12954 694274 13574 710042
rect 22954 711558 23574 711590
rect 22954 711322 22986 711558
rect 23222 711322 23306 711558
rect 23542 711322 23574 711558
rect 22954 711238 23574 711322
rect 22954 711002 22986 711238
rect 23222 711002 23306 711238
rect 23542 711002 23574 711238
rect 19234 709638 19854 709670
rect 19234 709402 19266 709638
rect 19502 709402 19586 709638
rect 19822 709402 19854 709638
rect 19234 709318 19854 709402
rect 19234 709082 19266 709318
rect 19502 709082 19586 709318
rect 19822 709082 19854 709318
rect 12954 694038 12986 694274
rect 13222 694038 13306 694274
rect 13542 694038 13574 694274
rect 12954 674274 13574 694038
rect 12954 674038 12986 674274
rect 13222 674038 13306 674274
rect 13542 674038 13574 674274
rect 12954 654274 13574 674038
rect 12954 654038 12986 654274
rect 13222 654038 13306 654274
rect 13542 654038 13574 654274
rect 12954 634274 13574 654038
rect 12954 634038 12986 634274
rect 13222 634038 13306 634274
rect 13542 634038 13574 634274
rect 12954 614274 13574 634038
rect 12954 614038 12986 614274
rect 13222 614038 13306 614274
rect 13542 614038 13574 614274
rect 12954 594274 13574 614038
rect 12954 594038 12986 594274
rect 13222 594038 13306 594274
rect 13542 594038 13574 594274
rect 12954 574274 13574 594038
rect 12954 574038 12986 574274
rect 13222 574038 13306 574274
rect 13542 574038 13574 574274
rect 12954 554274 13574 574038
rect 12954 554038 12986 554274
rect 13222 554038 13306 554274
rect 13542 554038 13574 554274
rect 12954 534274 13574 554038
rect 12954 534038 12986 534274
rect 13222 534038 13306 534274
rect 13542 534038 13574 534274
rect 12954 514274 13574 534038
rect 12954 514038 12986 514274
rect 13222 514038 13306 514274
rect 13542 514038 13574 514274
rect 12954 494274 13574 514038
rect 12954 494038 12986 494274
rect 13222 494038 13306 494274
rect 13542 494038 13574 494274
rect 12954 474274 13574 494038
rect 12954 474038 12986 474274
rect 13222 474038 13306 474274
rect 13542 474038 13574 474274
rect 12954 454274 13574 474038
rect 12954 454038 12986 454274
rect 13222 454038 13306 454274
rect 13542 454038 13574 454274
rect 12954 434274 13574 454038
rect 12954 434038 12986 434274
rect 13222 434038 13306 434274
rect 13542 434038 13574 434274
rect 12954 414274 13574 434038
rect 12954 414038 12986 414274
rect 13222 414038 13306 414274
rect 13542 414038 13574 414274
rect 12954 394274 13574 414038
rect 12954 394038 12986 394274
rect 13222 394038 13306 394274
rect 13542 394038 13574 394274
rect 12954 374274 13574 394038
rect 12954 374038 12986 374274
rect 13222 374038 13306 374274
rect 13542 374038 13574 374274
rect 12954 354274 13574 374038
rect 12954 354038 12986 354274
rect 13222 354038 13306 354274
rect 13542 354038 13574 354274
rect 12954 334274 13574 354038
rect 12954 334038 12986 334274
rect 13222 334038 13306 334274
rect 13542 334038 13574 334274
rect 12954 314274 13574 334038
rect 12954 314038 12986 314274
rect 13222 314038 13306 314274
rect 13542 314038 13574 314274
rect 12954 294274 13574 314038
rect 12954 294038 12986 294274
rect 13222 294038 13306 294274
rect 13542 294038 13574 294274
rect 12954 274274 13574 294038
rect 12954 274038 12986 274274
rect 13222 274038 13306 274274
rect 13542 274038 13574 274274
rect 12954 254274 13574 274038
rect 12954 254038 12986 254274
rect 13222 254038 13306 254274
rect 13542 254038 13574 254274
rect 12954 234274 13574 254038
rect 12954 234038 12986 234274
rect 13222 234038 13306 234274
rect 13542 234038 13574 234274
rect 12954 214274 13574 234038
rect 12954 214038 12986 214274
rect 13222 214038 13306 214274
rect 13542 214038 13574 214274
rect 12954 194274 13574 214038
rect 12954 194038 12986 194274
rect 13222 194038 13306 194274
rect 13542 194038 13574 194274
rect 12954 174274 13574 194038
rect 12954 174038 12986 174274
rect 13222 174038 13306 174274
rect 13542 174038 13574 174274
rect 12954 154274 13574 174038
rect 12954 154038 12986 154274
rect 13222 154038 13306 154274
rect 13542 154038 13574 154274
rect 12954 134274 13574 154038
rect 12954 134038 12986 134274
rect 13222 134038 13306 134274
rect 13542 134038 13574 134274
rect 12954 114274 13574 134038
rect 12954 114038 12986 114274
rect 13222 114038 13306 114274
rect 13542 114038 13574 114274
rect 12954 94274 13574 114038
rect 12954 94038 12986 94274
rect 13222 94038 13306 94274
rect 13542 94038 13574 94274
rect 12954 74274 13574 94038
rect 12954 74038 12986 74274
rect 13222 74038 13306 74274
rect 13542 74038 13574 74274
rect 12954 54274 13574 74038
rect 12954 54038 12986 54274
rect 13222 54038 13306 54274
rect 13542 54038 13574 54274
rect 12954 34274 13574 54038
rect 12954 34038 12986 34274
rect 13222 34038 13306 34274
rect 13542 34038 13574 34274
rect 12954 14274 13574 34038
rect 12954 14038 12986 14274
rect 13222 14038 13306 14274
rect 13542 14038 13574 14274
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14038
rect 15514 707718 16134 707750
rect 15514 707482 15546 707718
rect 15782 707482 15866 707718
rect 16102 707482 16134 707718
rect 15514 707398 16134 707482
rect 15514 707162 15546 707398
rect 15782 707162 15866 707398
rect 16102 707162 16134 707398
rect 15514 696954 16134 707162
rect 15514 696718 15546 696954
rect 15782 696718 15866 696954
rect 16102 696718 16134 696954
rect 15514 676954 16134 696718
rect 15514 676718 15546 676954
rect 15782 676718 15866 676954
rect 16102 676718 16134 676954
rect 15514 656954 16134 676718
rect 15514 656718 15546 656954
rect 15782 656718 15866 656954
rect 16102 656718 16134 656954
rect 15514 636954 16134 656718
rect 15514 636718 15546 636954
rect 15782 636718 15866 636954
rect 16102 636718 16134 636954
rect 15514 616954 16134 636718
rect 15514 616718 15546 616954
rect 15782 616718 15866 616954
rect 16102 616718 16134 616954
rect 15514 596954 16134 616718
rect 15514 596718 15546 596954
rect 15782 596718 15866 596954
rect 16102 596718 16134 596954
rect 15514 576954 16134 596718
rect 15514 576718 15546 576954
rect 15782 576718 15866 576954
rect 16102 576718 16134 576954
rect 15514 556954 16134 576718
rect 15514 556718 15546 556954
rect 15782 556718 15866 556954
rect 16102 556718 16134 556954
rect 15514 536954 16134 556718
rect 15514 536718 15546 536954
rect 15782 536718 15866 536954
rect 16102 536718 16134 536954
rect 15514 516954 16134 536718
rect 15514 516718 15546 516954
rect 15782 516718 15866 516954
rect 16102 516718 16134 516954
rect 15514 496954 16134 516718
rect 15514 496718 15546 496954
rect 15782 496718 15866 496954
rect 16102 496718 16134 496954
rect 15514 476954 16134 496718
rect 15514 476718 15546 476954
rect 15782 476718 15866 476954
rect 16102 476718 16134 476954
rect 15514 456954 16134 476718
rect 15514 456718 15546 456954
rect 15782 456718 15866 456954
rect 16102 456718 16134 456954
rect 15514 436954 16134 456718
rect 15514 436718 15546 436954
rect 15782 436718 15866 436954
rect 16102 436718 16134 436954
rect 15514 416954 16134 436718
rect 15514 416718 15546 416954
rect 15782 416718 15866 416954
rect 16102 416718 16134 416954
rect 15514 396954 16134 416718
rect 15514 396718 15546 396954
rect 15782 396718 15866 396954
rect 16102 396718 16134 396954
rect 15514 376954 16134 396718
rect 15514 376718 15546 376954
rect 15782 376718 15866 376954
rect 16102 376718 16134 376954
rect 15514 356954 16134 376718
rect 15514 356718 15546 356954
rect 15782 356718 15866 356954
rect 16102 356718 16134 356954
rect 15514 336954 16134 356718
rect 15514 336718 15546 336954
rect 15782 336718 15866 336954
rect 16102 336718 16134 336954
rect 15514 316954 16134 336718
rect 15514 316718 15546 316954
rect 15782 316718 15866 316954
rect 16102 316718 16134 316954
rect 15514 296954 16134 316718
rect 15514 296718 15546 296954
rect 15782 296718 15866 296954
rect 16102 296718 16134 296954
rect 15514 276954 16134 296718
rect 15514 276718 15546 276954
rect 15782 276718 15866 276954
rect 16102 276718 16134 276954
rect 15514 256954 16134 276718
rect 15514 256718 15546 256954
rect 15782 256718 15866 256954
rect 16102 256718 16134 256954
rect 15514 236954 16134 256718
rect 15514 236718 15546 236954
rect 15782 236718 15866 236954
rect 16102 236718 16134 236954
rect 15514 216954 16134 236718
rect 15514 216718 15546 216954
rect 15782 216718 15866 216954
rect 16102 216718 16134 216954
rect 15514 196954 16134 216718
rect 15514 196718 15546 196954
rect 15782 196718 15866 196954
rect 16102 196718 16134 196954
rect 15514 176954 16134 196718
rect 15514 176718 15546 176954
rect 15782 176718 15866 176954
rect 16102 176718 16134 176954
rect 15514 156954 16134 176718
rect 15514 156718 15546 156954
rect 15782 156718 15866 156954
rect 16102 156718 16134 156954
rect 15514 136954 16134 156718
rect 15514 136718 15546 136954
rect 15782 136718 15866 136954
rect 16102 136718 16134 136954
rect 15514 116954 16134 136718
rect 15514 116718 15546 116954
rect 15782 116718 15866 116954
rect 16102 116718 16134 116954
rect 15514 96954 16134 116718
rect 15514 96718 15546 96954
rect 15782 96718 15866 96954
rect 16102 96718 16134 96954
rect 15514 76954 16134 96718
rect 15514 76718 15546 76954
rect 15782 76718 15866 76954
rect 16102 76718 16134 76954
rect 15514 56954 16134 76718
rect 15514 56718 15546 56954
rect 15782 56718 15866 56954
rect 16102 56718 16134 56954
rect 15514 36954 16134 56718
rect 15514 36718 15546 36954
rect 15782 36718 15866 36954
rect 16102 36718 16134 36954
rect 15514 16954 16134 36718
rect 15514 16718 15546 16954
rect 15782 16718 15866 16954
rect 16102 16718 16134 16954
rect 15514 -3226 16134 16718
rect 15514 -3462 15546 -3226
rect 15782 -3462 15866 -3226
rect 16102 -3462 16134 -3226
rect 15514 -3546 16134 -3462
rect 15514 -3782 15546 -3546
rect 15782 -3782 15866 -3546
rect 16102 -3782 16134 -3546
rect 15514 -3814 16134 -3782
rect 19234 700614 19854 709082
rect 19234 700378 19266 700614
rect 19502 700378 19586 700614
rect 19822 700378 19854 700614
rect 19234 680614 19854 700378
rect 19234 680378 19266 680614
rect 19502 680378 19586 680614
rect 19822 680378 19854 680614
rect 19234 660614 19854 680378
rect 19234 660378 19266 660614
rect 19502 660378 19586 660614
rect 19822 660378 19854 660614
rect 19234 640614 19854 660378
rect 19234 640378 19266 640614
rect 19502 640378 19586 640614
rect 19822 640378 19854 640614
rect 19234 620614 19854 640378
rect 19234 620378 19266 620614
rect 19502 620378 19586 620614
rect 19822 620378 19854 620614
rect 19234 600614 19854 620378
rect 19234 600378 19266 600614
rect 19502 600378 19586 600614
rect 19822 600378 19854 600614
rect 19234 580614 19854 600378
rect 19234 580378 19266 580614
rect 19502 580378 19586 580614
rect 19822 580378 19854 580614
rect 19234 560614 19854 580378
rect 19234 560378 19266 560614
rect 19502 560378 19586 560614
rect 19822 560378 19854 560614
rect 19234 540614 19854 560378
rect 19234 540378 19266 540614
rect 19502 540378 19586 540614
rect 19822 540378 19854 540614
rect 19234 520614 19854 540378
rect 19234 520378 19266 520614
rect 19502 520378 19586 520614
rect 19822 520378 19854 520614
rect 19234 500614 19854 520378
rect 19234 500378 19266 500614
rect 19502 500378 19586 500614
rect 19822 500378 19854 500614
rect 19234 480614 19854 500378
rect 19234 480378 19266 480614
rect 19502 480378 19586 480614
rect 19822 480378 19854 480614
rect 19234 460614 19854 480378
rect 19234 460378 19266 460614
rect 19502 460378 19586 460614
rect 19822 460378 19854 460614
rect 19234 440614 19854 460378
rect 19234 440378 19266 440614
rect 19502 440378 19586 440614
rect 19822 440378 19854 440614
rect 19234 420614 19854 440378
rect 19234 420378 19266 420614
rect 19502 420378 19586 420614
rect 19822 420378 19854 420614
rect 19234 400614 19854 420378
rect 19234 400378 19266 400614
rect 19502 400378 19586 400614
rect 19822 400378 19854 400614
rect 19234 380614 19854 400378
rect 19234 380378 19266 380614
rect 19502 380378 19586 380614
rect 19822 380378 19854 380614
rect 19234 360614 19854 380378
rect 19234 360378 19266 360614
rect 19502 360378 19586 360614
rect 19822 360378 19854 360614
rect 19234 340614 19854 360378
rect 19234 340378 19266 340614
rect 19502 340378 19586 340614
rect 19822 340378 19854 340614
rect 19234 320614 19854 340378
rect 19234 320378 19266 320614
rect 19502 320378 19586 320614
rect 19822 320378 19854 320614
rect 19234 300614 19854 320378
rect 19234 300378 19266 300614
rect 19502 300378 19586 300614
rect 19822 300378 19854 300614
rect 19234 280614 19854 300378
rect 19234 280378 19266 280614
rect 19502 280378 19586 280614
rect 19822 280378 19854 280614
rect 19234 260614 19854 280378
rect 19234 260378 19266 260614
rect 19502 260378 19586 260614
rect 19822 260378 19854 260614
rect 19234 240614 19854 260378
rect 19234 240378 19266 240614
rect 19502 240378 19586 240614
rect 19822 240378 19854 240614
rect 19234 220614 19854 240378
rect 19234 220378 19266 220614
rect 19502 220378 19586 220614
rect 19822 220378 19854 220614
rect 19234 200614 19854 220378
rect 19234 200378 19266 200614
rect 19502 200378 19586 200614
rect 19822 200378 19854 200614
rect 19234 180614 19854 200378
rect 19234 180378 19266 180614
rect 19502 180378 19586 180614
rect 19822 180378 19854 180614
rect 19234 160614 19854 180378
rect 19234 160378 19266 160614
rect 19502 160378 19586 160614
rect 19822 160378 19854 160614
rect 19234 140614 19854 160378
rect 19234 140378 19266 140614
rect 19502 140378 19586 140614
rect 19822 140378 19854 140614
rect 19234 120614 19854 140378
rect 19234 120378 19266 120614
rect 19502 120378 19586 120614
rect 19822 120378 19854 120614
rect 19234 100614 19854 120378
rect 19234 100378 19266 100614
rect 19502 100378 19586 100614
rect 19822 100378 19854 100614
rect 19234 80614 19854 100378
rect 19234 80378 19266 80614
rect 19502 80378 19586 80614
rect 19822 80378 19854 80614
rect 19234 60614 19854 80378
rect 19234 60378 19266 60614
rect 19502 60378 19586 60614
rect 19822 60378 19854 60614
rect 19234 40614 19854 60378
rect 19234 40378 19266 40614
rect 19502 40378 19586 40614
rect 19822 40378 19854 40614
rect 19234 20614 19854 40378
rect 19234 20378 19266 20614
rect 19502 20378 19586 20614
rect 19822 20378 19854 20614
rect 19234 -5146 19854 20378
rect 21794 704838 22414 705830
rect 21794 704602 21826 704838
rect 22062 704602 22146 704838
rect 22382 704602 22414 704838
rect 21794 704518 22414 704602
rect 21794 704282 21826 704518
rect 22062 704282 22146 704518
rect 22382 704282 22414 704518
rect 21794 683294 22414 704282
rect 21794 683058 21826 683294
rect 22062 683058 22146 683294
rect 22382 683058 22414 683294
rect 21794 663294 22414 683058
rect 21794 663058 21826 663294
rect 22062 663058 22146 663294
rect 22382 663058 22414 663294
rect 21794 643294 22414 663058
rect 21794 643058 21826 643294
rect 22062 643058 22146 643294
rect 22382 643058 22414 643294
rect 21794 623294 22414 643058
rect 21794 623058 21826 623294
rect 22062 623058 22146 623294
rect 22382 623058 22414 623294
rect 21794 603294 22414 623058
rect 21794 603058 21826 603294
rect 22062 603058 22146 603294
rect 22382 603058 22414 603294
rect 21794 583294 22414 603058
rect 21794 583058 21826 583294
rect 22062 583058 22146 583294
rect 22382 583058 22414 583294
rect 21794 563294 22414 583058
rect 21794 563058 21826 563294
rect 22062 563058 22146 563294
rect 22382 563058 22414 563294
rect 21794 543294 22414 563058
rect 21794 543058 21826 543294
rect 22062 543058 22146 543294
rect 22382 543058 22414 543294
rect 21794 523294 22414 543058
rect 21794 523058 21826 523294
rect 22062 523058 22146 523294
rect 22382 523058 22414 523294
rect 21794 503294 22414 523058
rect 21794 503058 21826 503294
rect 22062 503058 22146 503294
rect 22382 503058 22414 503294
rect 21794 483294 22414 503058
rect 21794 483058 21826 483294
rect 22062 483058 22146 483294
rect 22382 483058 22414 483294
rect 21794 463294 22414 483058
rect 21794 463058 21826 463294
rect 22062 463058 22146 463294
rect 22382 463058 22414 463294
rect 21794 443294 22414 463058
rect 21794 443058 21826 443294
rect 22062 443058 22146 443294
rect 22382 443058 22414 443294
rect 21794 423294 22414 443058
rect 21794 423058 21826 423294
rect 22062 423058 22146 423294
rect 22382 423058 22414 423294
rect 21794 403294 22414 423058
rect 21794 403058 21826 403294
rect 22062 403058 22146 403294
rect 22382 403058 22414 403294
rect 21794 383294 22414 403058
rect 21794 383058 21826 383294
rect 22062 383058 22146 383294
rect 22382 383058 22414 383294
rect 21794 363294 22414 383058
rect 21794 363058 21826 363294
rect 22062 363058 22146 363294
rect 22382 363058 22414 363294
rect 21794 343294 22414 363058
rect 21794 343058 21826 343294
rect 22062 343058 22146 343294
rect 22382 343058 22414 343294
rect 21794 323294 22414 343058
rect 21794 323058 21826 323294
rect 22062 323058 22146 323294
rect 22382 323058 22414 323294
rect 21794 303294 22414 323058
rect 21794 303058 21826 303294
rect 22062 303058 22146 303294
rect 22382 303058 22414 303294
rect 21794 283294 22414 303058
rect 21794 283058 21826 283294
rect 22062 283058 22146 283294
rect 22382 283058 22414 283294
rect 21794 263294 22414 283058
rect 21794 263058 21826 263294
rect 22062 263058 22146 263294
rect 22382 263058 22414 263294
rect 21794 243294 22414 263058
rect 21794 243058 21826 243294
rect 22062 243058 22146 243294
rect 22382 243058 22414 243294
rect 21794 223294 22414 243058
rect 21794 223058 21826 223294
rect 22062 223058 22146 223294
rect 22382 223058 22414 223294
rect 21794 203294 22414 223058
rect 21794 203058 21826 203294
rect 22062 203058 22146 203294
rect 22382 203058 22414 203294
rect 21794 183294 22414 203058
rect 21794 183058 21826 183294
rect 22062 183058 22146 183294
rect 22382 183058 22414 183294
rect 21794 163294 22414 183058
rect 21794 163058 21826 163294
rect 22062 163058 22146 163294
rect 22382 163058 22414 163294
rect 21794 143294 22414 163058
rect 21794 143058 21826 143294
rect 22062 143058 22146 143294
rect 22382 143058 22414 143294
rect 21794 123294 22414 143058
rect 21794 123058 21826 123294
rect 22062 123058 22146 123294
rect 22382 123058 22414 123294
rect 21794 103294 22414 123058
rect 21794 103058 21826 103294
rect 22062 103058 22146 103294
rect 22382 103058 22414 103294
rect 21794 83294 22414 103058
rect 21794 83058 21826 83294
rect 22062 83058 22146 83294
rect 22382 83058 22414 83294
rect 21794 63294 22414 83058
rect 21794 63058 21826 63294
rect 22062 63058 22146 63294
rect 22382 63058 22414 63294
rect 21794 43294 22414 63058
rect 21794 43058 21826 43294
rect 22062 43058 22146 43294
rect 22382 43058 22414 43294
rect 21794 23294 22414 43058
rect 21794 23058 21826 23294
rect 22062 23058 22146 23294
rect 22382 23058 22414 23294
rect 21794 3294 22414 23058
rect 21794 3058 21826 3294
rect 22062 3058 22146 3294
rect 22382 3058 22414 3294
rect 21794 -346 22414 3058
rect 21794 -582 21826 -346
rect 22062 -582 22146 -346
rect 22382 -582 22414 -346
rect 21794 -666 22414 -582
rect 21794 -902 21826 -666
rect 22062 -902 22146 -666
rect 22382 -902 22414 -666
rect 21794 -1894 22414 -902
rect 22954 684274 23574 711002
rect 32954 710598 33574 711590
rect 32954 710362 32986 710598
rect 33222 710362 33306 710598
rect 33542 710362 33574 710598
rect 32954 710278 33574 710362
rect 32954 710042 32986 710278
rect 33222 710042 33306 710278
rect 33542 710042 33574 710278
rect 29234 708678 29854 709670
rect 29234 708442 29266 708678
rect 29502 708442 29586 708678
rect 29822 708442 29854 708678
rect 29234 708358 29854 708442
rect 29234 708122 29266 708358
rect 29502 708122 29586 708358
rect 29822 708122 29854 708358
rect 22954 684038 22986 684274
rect 23222 684038 23306 684274
rect 23542 684038 23574 684274
rect 22954 664274 23574 684038
rect 22954 664038 22986 664274
rect 23222 664038 23306 664274
rect 23542 664038 23574 664274
rect 22954 644274 23574 664038
rect 22954 644038 22986 644274
rect 23222 644038 23306 644274
rect 23542 644038 23574 644274
rect 22954 624274 23574 644038
rect 22954 624038 22986 624274
rect 23222 624038 23306 624274
rect 23542 624038 23574 624274
rect 22954 604274 23574 624038
rect 22954 604038 22986 604274
rect 23222 604038 23306 604274
rect 23542 604038 23574 604274
rect 22954 584274 23574 604038
rect 22954 584038 22986 584274
rect 23222 584038 23306 584274
rect 23542 584038 23574 584274
rect 22954 564274 23574 584038
rect 22954 564038 22986 564274
rect 23222 564038 23306 564274
rect 23542 564038 23574 564274
rect 22954 544274 23574 564038
rect 22954 544038 22986 544274
rect 23222 544038 23306 544274
rect 23542 544038 23574 544274
rect 22954 524274 23574 544038
rect 22954 524038 22986 524274
rect 23222 524038 23306 524274
rect 23542 524038 23574 524274
rect 22954 504274 23574 524038
rect 22954 504038 22986 504274
rect 23222 504038 23306 504274
rect 23542 504038 23574 504274
rect 22954 484274 23574 504038
rect 22954 484038 22986 484274
rect 23222 484038 23306 484274
rect 23542 484038 23574 484274
rect 22954 464274 23574 484038
rect 22954 464038 22986 464274
rect 23222 464038 23306 464274
rect 23542 464038 23574 464274
rect 22954 444274 23574 464038
rect 22954 444038 22986 444274
rect 23222 444038 23306 444274
rect 23542 444038 23574 444274
rect 22954 424274 23574 444038
rect 22954 424038 22986 424274
rect 23222 424038 23306 424274
rect 23542 424038 23574 424274
rect 22954 404274 23574 424038
rect 22954 404038 22986 404274
rect 23222 404038 23306 404274
rect 23542 404038 23574 404274
rect 22954 384274 23574 404038
rect 22954 384038 22986 384274
rect 23222 384038 23306 384274
rect 23542 384038 23574 384274
rect 22954 364274 23574 384038
rect 22954 364038 22986 364274
rect 23222 364038 23306 364274
rect 23542 364038 23574 364274
rect 22954 344274 23574 364038
rect 22954 344038 22986 344274
rect 23222 344038 23306 344274
rect 23542 344038 23574 344274
rect 22954 324274 23574 344038
rect 22954 324038 22986 324274
rect 23222 324038 23306 324274
rect 23542 324038 23574 324274
rect 22954 304274 23574 324038
rect 22954 304038 22986 304274
rect 23222 304038 23306 304274
rect 23542 304038 23574 304274
rect 22954 284274 23574 304038
rect 22954 284038 22986 284274
rect 23222 284038 23306 284274
rect 23542 284038 23574 284274
rect 22954 264274 23574 284038
rect 22954 264038 22986 264274
rect 23222 264038 23306 264274
rect 23542 264038 23574 264274
rect 22954 244274 23574 264038
rect 22954 244038 22986 244274
rect 23222 244038 23306 244274
rect 23542 244038 23574 244274
rect 22954 224274 23574 244038
rect 22954 224038 22986 224274
rect 23222 224038 23306 224274
rect 23542 224038 23574 224274
rect 22954 204274 23574 224038
rect 22954 204038 22986 204274
rect 23222 204038 23306 204274
rect 23542 204038 23574 204274
rect 22954 184274 23574 204038
rect 22954 184038 22986 184274
rect 23222 184038 23306 184274
rect 23542 184038 23574 184274
rect 22954 164274 23574 184038
rect 22954 164038 22986 164274
rect 23222 164038 23306 164274
rect 23542 164038 23574 164274
rect 22954 144274 23574 164038
rect 22954 144038 22986 144274
rect 23222 144038 23306 144274
rect 23542 144038 23574 144274
rect 22954 124274 23574 144038
rect 22954 124038 22986 124274
rect 23222 124038 23306 124274
rect 23542 124038 23574 124274
rect 22954 104274 23574 124038
rect 22954 104038 22986 104274
rect 23222 104038 23306 104274
rect 23542 104038 23574 104274
rect 22954 84274 23574 104038
rect 22954 84038 22986 84274
rect 23222 84038 23306 84274
rect 23542 84038 23574 84274
rect 22954 64274 23574 84038
rect 22954 64038 22986 64274
rect 23222 64038 23306 64274
rect 23542 64038 23574 64274
rect 22954 44274 23574 64038
rect 22954 44038 22986 44274
rect 23222 44038 23306 44274
rect 23542 44038 23574 44274
rect 22954 24274 23574 44038
rect 22954 24038 22986 24274
rect 23222 24038 23306 24274
rect 23542 24038 23574 24274
rect 19234 -5382 19266 -5146
rect 19502 -5382 19586 -5146
rect 19822 -5382 19854 -5146
rect 19234 -5466 19854 -5382
rect 19234 -5702 19266 -5466
rect 19502 -5702 19586 -5466
rect 19822 -5702 19854 -5466
rect 19234 -5734 19854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 22954 -7066 23574 24038
rect 25514 706758 26134 707750
rect 25514 706522 25546 706758
rect 25782 706522 25866 706758
rect 26102 706522 26134 706758
rect 25514 706438 26134 706522
rect 25514 706202 25546 706438
rect 25782 706202 25866 706438
rect 26102 706202 26134 706438
rect 25514 686954 26134 706202
rect 25514 686718 25546 686954
rect 25782 686718 25866 686954
rect 26102 686718 26134 686954
rect 25514 666954 26134 686718
rect 29234 690614 29854 708122
rect 29234 690378 29266 690614
rect 29502 690378 29586 690614
rect 29822 690378 29854 690614
rect 29234 675308 29854 690378
rect 31794 705798 32414 705830
rect 31794 705562 31826 705798
rect 32062 705562 32146 705798
rect 32382 705562 32414 705798
rect 31794 705478 32414 705562
rect 31794 705242 31826 705478
rect 32062 705242 32146 705478
rect 32382 705242 32414 705478
rect 31794 693294 32414 705242
rect 31794 693058 31826 693294
rect 32062 693058 32146 693294
rect 32382 693058 32414 693294
rect 31794 675308 32414 693058
rect 32954 694274 33574 710042
rect 42954 711558 43574 711590
rect 42954 711322 42986 711558
rect 43222 711322 43306 711558
rect 43542 711322 43574 711558
rect 42954 711238 43574 711322
rect 42954 711002 42986 711238
rect 43222 711002 43306 711238
rect 43542 711002 43574 711238
rect 39234 709638 39854 709670
rect 39234 709402 39266 709638
rect 39502 709402 39586 709638
rect 39822 709402 39854 709638
rect 39234 709318 39854 709402
rect 39234 709082 39266 709318
rect 39502 709082 39586 709318
rect 39822 709082 39854 709318
rect 32954 694038 32986 694274
rect 33222 694038 33306 694274
rect 33542 694038 33574 694274
rect 32954 675308 33574 694038
rect 35514 707718 36134 707750
rect 35514 707482 35546 707718
rect 35782 707482 35866 707718
rect 36102 707482 36134 707718
rect 35514 707398 36134 707482
rect 35514 707162 35546 707398
rect 35782 707162 35866 707398
rect 36102 707162 36134 707398
rect 35514 696954 36134 707162
rect 35514 696718 35546 696954
rect 35782 696718 35866 696954
rect 36102 696718 36134 696954
rect 35514 676954 36134 696718
rect 35514 676718 35546 676954
rect 35782 676718 35866 676954
rect 36102 676718 36134 676954
rect 35514 675308 36134 676718
rect 39234 700614 39854 709082
rect 39234 700378 39266 700614
rect 39502 700378 39586 700614
rect 39822 700378 39854 700614
rect 39234 680614 39854 700378
rect 39234 680378 39266 680614
rect 39502 680378 39586 680614
rect 39822 680378 39854 680614
rect 39234 675308 39854 680378
rect 41794 704838 42414 705830
rect 41794 704602 41826 704838
rect 42062 704602 42146 704838
rect 42382 704602 42414 704838
rect 41794 704518 42414 704602
rect 41794 704282 41826 704518
rect 42062 704282 42146 704518
rect 42382 704282 42414 704518
rect 41794 683294 42414 704282
rect 41794 683058 41826 683294
rect 42062 683058 42146 683294
rect 42382 683058 42414 683294
rect 41794 675308 42414 683058
rect 42954 684274 43574 711002
rect 52954 710598 53574 711590
rect 52954 710362 52986 710598
rect 53222 710362 53306 710598
rect 53542 710362 53574 710598
rect 52954 710278 53574 710362
rect 52954 710042 52986 710278
rect 53222 710042 53306 710278
rect 53542 710042 53574 710278
rect 49234 708678 49854 709670
rect 49234 708442 49266 708678
rect 49502 708442 49586 708678
rect 49822 708442 49854 708678
rect 49234 708358 49854 708442
rect 49234 708122 49266 708358
rect 49502 708122 49586 708358
rect 49822 708122 49854 708358
rect 42954 684038 42986 684274
rect 43222 684038 43306 684274
rect 43542 684038 43574 684274
rect 42954 675308 43574 684038
rect 45514 706758 46134 707750
rect 45514 706522 45546 706758
rect 45782 706522 45866 706758
rect 46102 706522 46134 706758
rect 45514 706438 46134 706522
rect 45514 706202 45546 706438
rect 45782 706202 45866 706438
rect 46102 706202 46134 706438
rect 45514 686954 46134 706202
rect 45514 686718 45546 686954
rect 45782 686718 45866 686954
rect 46102 686718 46134 686954
rect 45514 675308 46134 686718
rect 49234 690614 49854 708122
rect 49234 690378 49266 690614
rect 49502 690378 49586 690614
rect 49822 690378 49854 690614
rect 49234 675308 49854 690378
rect 51794 705798 52414 705830
rect 51794 705562 51826 705798
rect 52062 705562 52146 705798
rect 52382 705562 52414 705798
rect 51794 705478 52414 705562
rect 51794 705242 51826 705478
rect 52062 705242 52146 705478
rect 52382 705242 52414 705478
rect 51794 693294 52414 705242
rect 51794 693058 51826 693294
rect 52062 693058 52146 693294
rect 52382 693058 52414 693294
rect 51794 675308 52414 693058
rect 52954 694274 53574 710042
rect 62954 711558 63574 711590
rect 62954 711322 62986 711558
rect 63222 711322 63306 711558
rect 63542 711322 63574 711558
rect 62954 711238 63574 711322
rect 62954 711002 62986 711238
rect 63222 711002 63306 711238
rect 63542 711002 63574 711238
rect 59234 709638 59854 709670
rect 59234 709402 59266 709638
rect 59502 709402 59586 709638
rect 59822 709402 59854 709638
rect 59234 709318 59854 709402
rect 59234 709082 59266 709318
rect 59502 709082 59586 709318
rect 59822 709082 59854 709318
rect 52954 694038 52986 694274
rect 53222 694038 53306 694274
rect 53542 694038 53574 694274
rect 52954 675308 53574 694038
rect 55514 707718 56134 707750
rect 55514 707482 55546 707718
rect 55782 707482 55866 707718
rect 56102 707482 56134 707718
rect 55514 707398 56134 707482
rect 55514 707162 55546 707398
rect 55782 707162 55866 707398
rect 56102 707162 56134 707398
rect 55514 696954 56134 707162
rect 55514 696718 55546 696954
rect 55782 696718 55866 696954
rect 56102 696718 56134 696954
rect 55514 676954 56134 696718
rect 55514 676718 55546 676954
rect 55782 676718 55866 676954
rect 56102 676718 56134 676954
rect 55514 675308 56134 676718
rect 59234 700614 59854 709082
rect 59234 700378 59266 700614
rect 59502 700378 59586 700614
rect 59822 700378 59854 700614
rect 59234 680614 59854 700378
rect 59234 680378 59266 680614
rect 59502 680378 59586 680614
rect 59822 680378 59854 680614
rect 59234 675308 59854 680378
rect 61794 704838 62414 705830
rect 61794 704602 61826 704838
rect 62062 704602 62146 704838
rect 62382 704602 62414 704838
rect 61794 704518 62414 704602
rect 61794 704282 61826 704518
rect 62062 704282 62146 704518
rect 62382 704282 62414 704518
rect 61794 683294 62414 704282
rect 61794 683058 61826 683294
rect 62062 683058 62146 683294
rect 62382 683058 62414 683294
rect 61794 675308 62414 683058
rect 62954 684274 63574 711002
rect 72954 710598 73574 711590
rect 72954 710362 72986 710598
rect 73222 710362 73306 710598
rect 73542 710362 73574 710598
rect 72954 710278 73574 710362
rect 72954 710042 72986 710278
rect 73222 710042 73306 710278
rect 73542 710042 73574 710278
rect 69234 708678 69854 709670
rect 69234 708442 69266 708678
rect 69502 708442 69586 708678
rect 69822 708442 69854 708678
rect 69234 708358 69854 708442
rect 69234 708122 69266 708358
rect 69502 708122 69586 708358
rect 69822 708122 69854 708358
rect 62954 684038 62986 684274
rect 63222 684038 63306 684274
rect 63542 684038 63574 684274
rect 62954 675308 63574 684038
rect 65514 706758 66134 707750
rect 65514 706522 65546 706758
rect 65782 706522 65866 706758
rect 66102 706522 66134 706758
rect 65514 706438 66134 706522
rect 65514 706202 65546 706438
rect 65782 706202 65866 706438
rect 66102 706202 66134 706438
rect 65514 686954 66134 706202
rect 65514 686718 65546 686954
rect 65782 686718 65866 686954
rect 66102 686718 66134 686954
rect 65514 675308 66134 686718
rect 69234 690614 69854 708122
rect 69234 690378 69266 690614
rect 69502 690378 69586 690614
rect 69822 690378 69854 690614
rect 69234 675308 69854 690378
rect 71794 705798 72414 705830
rect 71794 705562 71826 705798
rect 72062 705562 72146 705798
rect 72382 705562 72414 705798
rect 71794 705478 72414 705562
rect 71794 705242 71826 705478
rect 72062 705242 72146 705478
rect 72382 705242 72414 705478
rect 71794 693294 72414 705242
rect 71794 693058 71826 693294
rect 72062 693058 72146 693294
rect 72382 693058 72414 693294
rect 71794 675308 72414 693058
rect 72954 694274 73574 710042
rect 82954 711558 83574 711590
rect 82954 711322 82986 711558
rect 83222 711322 83306 711558
rect 83542 711322 83574 711558
rect 82954 711238 83574 711322
rect 82954 711002 82986 711238
rect 83222 711002 83306 711238
rect 83542 711002 83574 711238
rect 79234 709638 79854 709670
rect 79234 709402 79266 709638
rect 79502 709402 79586 709638
rect 79822 709402 79854 709638
rect 79234 709318 79854 709402
rect 79234 709082 79266 709318
rect 79502 709082 79586 709318
rect 79822 709082 79854 709318
rect 72954 694038 72986 694274
rect 73222 694038 73306 694274
rect 73542 694038 73574 694274
rect 72954 675308 73574 694038
rect 75514 707718 76134 707750
rect 75514 707482 75546 707718
rect 75782 707482 75866 707718
rect 76102 707482 76134 707718
rect 75514 707398 76134 707482
rect 75514 707162 75546 707398
rect 75782 707162 75866 707398
rect 76102 707162 76134 707398
rect 75514 696954 76134 707162
rect 75514 696718 75546 696954
rect 75782 696718 75866 696954
rect 76102 696718 76134 696954
rect 75514 676954 76134 696718
rect 75514 676718 75546 676954
rect 75782 676718 75866 676954
rect 76102 676718 76134 676954
rect 75514 675308 76134 676718
rect 79234 700614 79854 709082
rect 79234 700378 79266 700614
rect 79502 700378 79586 700614
rect 79822 700378 79854 700614
rect 79234 680614 79854 700378
rect 79234 680378 79266 680614
rect 79502 680378 79586 680614
rect 79822 680378 79854 680614
rect 79234 675308 79854 680378
rect 81794 704838 82414 705830
rect 81794 704602 81826 704838
rect 82062 704602 82146 704838
rect 82382 704602 82414 704838
rect 81794 704518 82414 704602
rect 81794 704282 81826 704518
rect 82062 704282 82146 704518
rect 82382 704282 82414 704518
rect 81794 683294 82414 704282
rect 81794 683058 81826 683294
rect 82062 683058 82146 683294
rect 82382 683058 82414 683294
rect 81794 675308 82414 683058
rect 82954 684274 83574 711002
rect 92954 710598 93574 711590
rect 92954 710362 92986 710598
rect 93222 710362 93306 710598
rect 93542 710362 93574 710598
rect 92954 710278 93574 710362
rect 92954 710042 92986 710278
rect 93222 710042 93306 710278
rect 93542 710042 93574 710278
rect 89234 708678 89854 709670
rect 89234 708442 89266 708678
rect 89502 708442 89586 708678
rect 89822 708442 89854 708678
rect 89234 708358 89854 708442
rect 89234 708122 89266 708358
rect 89502 708122 89586 708358
rect 89822 708122 89854 708358
rect 82954 684038 82986 684274
rect 83222 684038 83306 684274
rect 83542 684038 83574 684274
rect 82954 675308 83574 684038
rect 85514 706758 86134 707750
rect 85514 706522 85546 706758
rect 85782 706522 85866 706758
rect 86102 706522 86134 706758
rect 85514 706438 86134 706522
rect 85514 706202 85546 706438
rect 85782 706202 85866 706438
rect 86102 706202 86134 706438
rect 85514 686954 86134 706202
rect 85514 686718 85546 686954
rect 85782 686718 85866 686954
rect 86102 686718 86134 686954
rect 85514 675308 86134 686718
rect 89234 690614 89854 708122
rect 89234 690378 89266 690614
rect 89502 690378 89586 690614
rect 89822 690378 89854 690614
rect 89234 675308 89854 690378
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 693294 92414 705242
rect 91794 693058 91826 693294
rect 92062 693058 92146 693294
rect 92382 693058 92414 693294
rect 91794 675308 92414 693058
rect 92954 694274 93574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 92954 694038 92986 694274
rect 93222 694038 93306 694274
rect 93542 694038 93574 694274
rect 92954 675308 93574 694038
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 95514 696954 96134 707162
rect 95514 696718 95546 696954
rect 95782 696718 95866 696954
rect 96102 696718 96134 696954
rect 95514 676954 96134 696718
rect 95514 676718 95546 676954
rect 95782 676718 95866 676954
rect 96102 676718 96134 676954
rect 95514 675308 96134 676718
rect 99234 700614 99854 709082
rect 99234 700378 99266 700614
rect 99502 700378 99586 700614
rect 99822 700378 99854 700614
rect 99234 680614 99854 700378
rect 99234 680378 99266 680614
rect 99502 680378 99586 680614
rect 99822 680378 99854 680614
rect 99234 675308 99854 680378
rect 101794 704838 102414 705830
rect 101794 704602 101826 704838
rect 102062 704602 102146 704838
rect 102382 704602 102414 704838
rect 101794 704518 102414 704602
rect 101794 704282 101826 704518
rect 102062 704282 102146 704518
rect 102382 704282 102414 704518
rect 101794 683294 102414 704282
rect 101794 683058 101826 683294
rect 102062 683058 102146 683294
rect 102382 683058 102414 683294
rect 101794 675308 102414 683058
rect 102954 684274 103574 711002
rect 112954 710598 113574 711590
rect 112954 710362 112986 710598
rect 113222 710362 113306 710598
rect 113542 710362 113574 710598
rect 112954 710278 113574 710362
rect 112954 710042 112986 710278
rect 113222 710042 113306 710278
rect 113542 710042 113574 710278
rect 109234 708678 109854 709670
rect 109234 708442 109266 708678
rect 109502 708442 109586 708678
rect 109822 708442 109854 708678
rect 109234 708358 109854 708442
rect 109234 708122 109266 708358
rect 109502 708122 109586 708358
rect 109822 708122 109854 708358
rect 102954 684038 102986 684274
rect 103222 684038 103306 684274
rect 103542 684038 103574 684274
rect 102954 675308 103574 684038
rect 105514 706758 106134 707750
rect 105514 706522 105546 706758
rect 105782 706522 105866 706758
rect 106102 706522 106134 706758
rect 105514 706438 106134 706522
rect 105514 706202 105546 706438
rect 105782 706202 105866 706438
rect 106102 706202 106134 706438
rect 105514 686954 106134 706202
rect 105514 686718 105546 686954
rect 105782 686718 105866 686954
rect 106102 686718 106134 686954
rect 105514 675308 106134 686718
rect 109234 690614 109854 708122
rect 109234 690378 109266 690614
rect 109502 690378 109586 690614
rect 109822 690378 109854 690614
rect 109234 675308 109854 690378
rect 111794 705798 112414 705830
rect 111794 705562 111826 705798
rect 112062 705562 112146 705798
rect 112382 705562 112414 705798
rect 111794 705478 112414 705562
rect 111794 705242 111826 705478
rect 112062 705242 112146 705478
rect 112382 705242 112414 705478
rect 111794 693294 112414 705242
rect 111794 693058 111826 693294
rect 112062 693058 112146 693294
rect 112382 693058 112414 693294
rect 111794 675308 112414 693058
rect 112954 694274 113574 710042
rect 122954 711558 123574 711590
rect 122954 711322 122986 711558
rect 123222 711322 123306 711558
rect 123542 711322 123574 711558
rect 122954 711238 123574 711322
rect 122954 711002 122986 711238
rect 123222 711002 123306 711238
rect 123542 711002 123574 711238
rect 119234 709638 119854 709670
rect 119234 709402 119266 709638
rect 119502 709402 119586 709638
rect 119822 709402 119854 709638
rect 119234 709318 119854 709402
rect 119234 709082 119266 709318
rect 119502 709082 119586 709318
rect 119822 709082 119854 709318
rect 112954 694038 112986 694274
rect 113222 694038 113306 694274
rect 113542 694038 113574 694274
rect 112954 675308 113574 694038
rect 115514 707718 116134 707750
rect 115514 707482 115546 707718
rect 115782 707482 115866 707718
rect 116102 707482 116134 707718
rect 115514 707398 116134 707482
rect 115514 707162 115546 707398
rect 115782 707162 115866 707398
rect 116102 707162 116134 707398
rect 115514 696954 116134 707162
rect 115514 696718 115546 696954
rect 115782 696718 115866 696954
rect 116102 696718 116134 696954
rect 115514 676954 116134 696718
rect 115514 676718 115546 676954
rect 115782 676718 115866 676954
rect 116102 676718 116134 676954
rect 115514 675308 116134 676718
rect 119234 700614 119854 709082
rect 119234 700378 119266 700614
rect 119502 700378 119586 700614
rect 119822 700378 119854 700614
rect 119234 680614 119854 700378
rect 119234 680378 119266 680614
rect 119502 680378 119586 680614
rect 119822 680378 119854 680614
rect 119234 675308 119854 680378
rect 121794 704838 122414 705830
rect 121794 704602 121826 704838
rect 122062 704602 122146 704838
rect 122382 704602 122414 704838
rect 121794 704518 122414 704602
rect 121794 704282 121826 704518
rect 122062 704282 122146 704518
rect 122382 704282 122414 704518
rect 121794 683294 122414 704282
rect 121794 683058 121826 683294
rect 122062 683058 122146 683294
rect 122382 683058 122414 683294
rect 121794 675308 122414 683058
rect 122954 684274 123574 711002
rect 132954 710598 133574 711590
rect 132954 710362 132986 710598
rect 133222 710362 133306 710598
rect 133542 710362 133574 710598
rect 132954 710278 133574 710362
rect 132954 710042 132986 710278
rect 133222 710042 133306 710278
rect 133542 710042 133574 710278
rect 129234 708678 129854 709670
rect 129234 708442 129266 708678
rect 129502 708442 129586 708678
rect 129822 708442 129854 708678
rect 129234 708358 129854 708442
rect 129234 708122 129266 708358
rect 129502 708122 129586 708358
rect 129822 708122 129854 708358
rect 122954 684038 122986 684274
rect 123222 684038 123306 684274
rect 123542 684038 123574 684274
rect 122954 675308 123574 684038
rect 125514 706758 126134 707750
rect 125514 706522 125546 706758
rect 125782 706522 125866 706758
rect 126102 706522 126134 706758
rect 125514 706438 126134 706522
rect 125514 706202 125546 706438
rect 125782 706202 125866 706438
rect 126102 706202 126134 706438
rect 125514 686954 126134 706202
rect 125514 686718 125546 686954
rect 125782 686718 125866 686954
rect 126102 686718 126134 686954
rect 125514 675308 126134 686718
rect 129234 690614 129854 708122
rect 129234 690378 129266 690614
rect 129502 690378 129586 690614
rect 129822 690378 129854 690614
rect 129234 675308 129854 690378
rect 131794 705798 132414 705830
rect 131794 705562 131826 705798
rect 132062 705562 132146 705798
rect 132382 705562 132414 705798
rect 131794 705478 132414 705562
rect 131794 705242 131826 705478
rect 132062 705242 132146 705478
rect 132382 705242 132414 705478
rect 131794 693294 132414 705242
rect 131794 693058 131826 693294
rect 132062 693058 132146 693294
rect 132382 693058 132414 693294
rect 131794 675308 132414 693058
rect 132954 694274 133574 710042
rect 142954 711558 143574 711590
rect 142954 711322 142986 711558
rect 143222 711322 143306 711558
rect 143542 711322 143574 711558
rect 142954 711238 143574 711322
rect 142954 711002 142986 711238
rect 143222 711002 143306 711238
rect 143542 711002 143574 711238
rect 139234 709638 139854 709670
rect 139234 709402 139266 709638
rect 139502 709402 139586 709638
rect 139822 709402 139854 709638
rect 139234 709318 139854 709402
rect 139234 709082 139266 709318
rect 139502 709082 139586 709318
rect 139822 709082 139854 709318
rect 132954 694038 132986 694274
rect 133222 694038 133306 694274
rect 133542 694038 133574 694274
rect 132954 675308 133574 694038
rect 135514 707718 136134 707750
rect 135514 707482 135546 707718
rect 135782 707482 135866 707718
rect 136102 707482 136134 707718
rect 135514 707398 136134 707482
rect 135514 707162 135546 707398
rect 135782 707162 135866 707398
rect 136102 707162 136134 707398
rect 135514 696954 136134 707162
rect 135514 696718 135546 696954
rect 135782 696718 135866 696954
rect 136102 696718 136134 696954
rect 135514 676954 136134 696718
rect 135514 676718 135546 676954
rect 135782 676718 135866 676954
rect 136102 676718 136134 676954
rect 135514 675308 136134 676718
rect 139234 700614 139854 709082
rect 139234 700378 139266 700614
rect 139502 700378 139586 700614
rect 139822 700378 139854 700614
rect 139234 680614 139854 700378
rect 139234 680378 139266 680614
rect 139502 680378 139586 680614
rect 139822 680378 139854 680614
rect 139234 675308 139854 680378
rect 141794 704838 142414 705830
rect 141794 704602 141826 704838
rect 142062 704602 142146 704838
rect 142382 704602 142414 704838
rect 141794 704518 142414 704602
rect 141794 704282 141826 704518
rect 142062 704282 142146 704518
rect 142382 704282 142414 704518
rect 141794 683294 142414 704282
rect 141794 683058 141826 683294
rect 142062 683058 142146 683294
rect 142382 683058 142414 683294
rect 141794 675308 142414 683058
rect 142954 684274 143574 711002
rect 152954 710598 153574 711590
rect 152954 710362 152986 710598
rect 153222 710362 153306 710598
rect 153542 710362 153574 710598
rect 152954 710278 153574 710362
rect 152954 710042 152986 710278
rect 153222 710042 153306 710278
rect 153542 710042 153574 710278
rect 149234 708678 149854 709670
rect 149234 708442 149266 708678
rect 149502 708442 149586 708678
rect 149822 708442 149854 708678
rect 149234 708358 149854 708442
rect 149234 708122 149266 708358
rect 149502 708122 149586 708358
rect 149822 708122 149854 708358
rect 142954 684038 142986 684274
rect 143222 684038 143306 684274
rect 143542 684038 143574 684274
rect 142954 675308 143574 684038
rect 145514 706758 146134 707750
rect 145514 706522 145546 706758
rect 145782 706522 145866 706758
rect 146102 706522 146134 706758
rect 145514 706438 146134 706522
rect 145514 706202 145546 706438
rect 145782 706202 145866 706438
rect 146102 706202 146134 706438
rect 145514 686954 146134 706202
rect 145514 686718 145546 686954
rect 145782 686718 145866 686954
rect 146102 686718 146134 686954
rect 145514 675308 146134 686718
rect 149234 690614 149854 708122
rect 149234 690378 149266 690614
rect 149502 690378 149586 690614
rect 149822 690378 149854 690614
rect 149234 675308 149854 690378
rect 151794 705798 152414 705830
rect 151794 705562 151826 705798
rect 152062 705562 152146 705798
rect 152382 705562 152414 705798
rect 151794 705478 152414 705562
rect 151794 705242 151826 705478
rect 152062 705242 152146 705478
rect 152382 705242 152414 705478
rect 151794 693294 152414 705242
rect 151794 693058 151826 693294
rect 152062 693058 152146 693294
rect 152382 693058 152414 693294
rect 151794 675308 152414 693058
rect 152954 694274 153574 710042
rect 162954 711558 163574 711590
rect 162954 711322 162986 711558
rect 163222 711322 163306 711558
rect 163542 711322 163574 711558
rect 162954 711238 163574 711322
rect 162954 711002 162986 711238
rect 163222 711002 163306 711238
rect 163542 711002 163574 711238
rect 159234 709638 159854 709670
rect 159234 709402 159266 709638
rect 159502 709402 159586 709638
rect 159822 709402 159854 709638
rect 159234 709318 159854 709402
rect 159234 709082 159266 709318
rect 159502 709082 159586 709318
rect 159822 709082 159854 709318
rect 152954 694038 152986 694274
rect 153222 694038 153306 694274
rect 153542 694038 153574 694274
rect 152954 675308 153574 694038
rect 155514 707718 156134 707750
rect 155514 707482 155546 707718
rect 155782 707482 155866 707718
rect 156102 707482 156134 707718
rect 155514 707398 156134 707482
rect 155514 707162 155546 707398
rect 155782 707162 155866 707398
rect 156102 707162 156134 707398
rect 155514 696954 156134 707162
rect 155514 696718 155546 696954
rect 155782 696718 155866 696954
rect 156102 696718 156134 696954
rect 155514 676954 156134 696718
rect 155514 676718 155546 676954
rect 155782 676718 155866 676954
rect 156102 676718 156134 676954
rect 155514 675308 156134 676718
rect 159234 700614 159854 709082
rect 159234 700378 159266 700614
rect 159502 700378 159586 700614
rect 159822 700378 159854 700614
rect 159234 680614 159854 700378
rect 159234 680378 159266 680614
rect 159502 680378 159586 680614
rect 159822 680378 159854 680614
rect 159234 675308 159854 680378
rect 161794 704838 162414 705830
rect 161794 704602 161826 704838
rect 162062 704602 162146 704838
rect 162382 704602 162414 704838
rect 161794 704518 162414 704602
rect 161794 704282 161826 704518
rect 162062 704282 162146 704518
rect 162382 704282 162414 704518
rect 161794 683294 162414 704282
rect 161794 683058 161826 683294
rect 162062 683058 162146 683294
rect 162382 683058 162414 683294
rect 161794 675308 162414 683058
rect 162954 684274 163574 711002
rect 172954 710598 173574 711590
rect 172954 710362 172986 710598
rect 173222 710362 173306 710598
rect 173542 710362 173574 710598
rect 172954 710278 173574 710362
rect 172954 710042 172986 710278
rect 173222 710042 173306 710278
rect 173542 710042 173574 710278
rect 169234 708678 169854 709670
rect 169234 708442 169266 708678
rect 169502 708442 169586 708678
rect 169822 708442 169854 708678
rect 169234 708358 169854 708442
rect 169234 708122 169266 708358
rect 169502 708122 169586 708358
rect 169822 708122 169854 708358
rect 162954 684038 162986 684274
rect 163222 684038 163306 684274
rect 163542 684038 163574 684274
rect 162954 675308 163574 684038
rect 165514 706758 166134 707750
rect 165514 706522 165546 706758
rect 165782 706522 165866 706758
rect 166102 706522 166134 706758
rect 165514 706438 166134 706522
rect 165514 706202 165546 706438
rect 165782 706202 165866 706438
rect 166102 706202 166134 706438
rect 165514 686954 166134 706202
rect 165514 686718 165546 686954
rect 165782 686718 165866 686954
rect 166102 686718 166134 686954
rect 165514 675308 166134 686718
rect 169234 690614 169854 708122
rect 169234 690378 169266 690614
rect 169502 690378 169586 690614
rect 169822 690378 169854 690614
rect 35755 674932 35821 674933
rect 35755 674868 35756 674932
rect 35820 674868 35821 674932
rect 35755 674867 35821 674868
rect 46795 674932 46861 674933
rect 46795 674868 46796 674932
rect 46860 674868 46861 674932
rect 46795 674867 46861 674868
rect 48083 674932 48149 674933
rect 48083 674868 48084 674932
rect 48148 674868 48149 674932
rect 48083 674867 48149 674868
rect 35758 673470 35818 674867
rect 35720 673410 35818 673470
rect 46798 673470 46858 674867
rect 48086 673470 48146 674867
rect 46798 673410 46932 673470
rect 48086 673410 48156 673470
rect 35720 673202 35780 673410
rect 46872 673202 46932 673410
rect 48096 673202 48156 673410
rect 25514 666718 25546 666954
rect 25782 666718 25866 666954
rect 26102 666718 26134 666954
rect 25514 646954 26134 666718
rect 169234 670614 169854 690378
rect 169234 670378 169266 670614
rect 169502 670378 169586 670614
rect 169822 670378 169854 670614
rect 30952 663294 31300 663456
rect 30952 663058 31008 663294
rect 31244 663058 31300 663294
rect 30952 662896 31300 663058
rect 165320 663294 165668 663456
rect 165320 663058 165376 663294
rect 165612 663058 165668 663294
rect 165320 662896 165668 663058
rect 30272 653294 30620 653456
rect 30272 653058 30328 653294
rect 30564 653058 30620 653294
rect 30272 652896 30620 653058
rect 166000 653294 166348 653456
rect 166000 653058 166056 653294
rect 166292 653058 166348 653294
rect 166000 652896 166348 653058
rect 25514 646718 25546 646954
rect 25782 646718 25866 646954
rect 26102 646718 26134 646954
rect 25514 626954 26134 646718
rect 169234 650614 169854 670378
rect 169234 650378 169266 650614
rect 169502 650378 169586 650614
rect 169822 650378 169854 650614
rect 30952 643294 31300 643456
rect 30952 643058 31008 643294
rect 31244 643058 31300 643294
rect 30952 642896 31300 643058
rect 165320 643294 165668 643456
rect 165320 643058 165376 643294
rect 165612 643058 165668 643294
rect 165320 642896 165668 643058
rect 30272 633294 30620 633456
rect 30272 633058 30328 633294
rect 30564 633058 30620 633294
rect 30272 632896 30620 633058
rect 166000 633294 166348 633456
rect 166000 633058 166056 633294
rect 166292 633058 166348 633294
rect 166000 632896 166348 633058
rect 25514 626718 25546 626954
rect 25782 626718 25866 626954
rect 26102 626718 26134 626954
rect 25514 606954 26134 626718
rect 169234 630614 169854 650378
rect 169234 630378 169266 630614
rect 169502 630378 169586 630614
rect 169822 630378 169854 630614
rect 30952 623294 31300 623456
rect 30952 623058 31008 623294
rect 31244 623058 31300 623294
rect 30952 622896 31300 623058
rect 165320 623294 165668 623456
rect 165320 623058 165376 623294
rect 165612 623058 165668 623294
rect 165320 622896 165668 623058
rect 30272 613294 30620 613456
rect 30272 613058 30328 613294
rect 30564 613058 30620 613294
rect 30272 612896 30620 613058
rect 166000 613294 166348 613456
rect 166000 613058 166056 613294
rect 166292 613058 166348 613294
rect 166000 612896 166348 613058
rect 25514 606718 25546 606954
rect 25782 606718 25866 606954
rect 26102 606718 26134 606954
rect 25514 586954 26134 606718
rect 169234 610614 169854 630378
rect 169234 610378 169266 610614
rect 169502 610378 169586 610614
rect 169822 610378 169854 610614
rect 30952 603294 31300 603456
rect 30952 603058 31008 603294
rect 31244 603058 31300 603294
rect 30952 602896 31300 603058
rect 165320 603294 165668 603456
rect 165320 603058 165376 603294
rect 165612 603058 165668 603294
rect 165320 602896 165668 603058
rect 30272 593294 30620 593456
rect 30272 593058 30328 593294
rect 30564 593058 30620 593294
rect 30272 592896 30620 593058
rect 166000 593294 166348 593456
rect 166000 593058 166056 593294
rect 166292 593058 166348 593294
rect 166000 592896 166348 593058
rect 169234 590614 169854 610378
rect 169234 590378 169266 590614
rect 169502 590378 169586 590614
rect 169822 590378 169854 590614
rect 43200 589250 43260 590106
rect 43118 589190 43260 589250
rect 43336 589250 43396 590106
rect 60608 589290 60668 590106
rect 63192 589290 63252 590106
rect 65640 589290 65700 590106
rect 43336 589190 43730 589250
rect 43118 588165 43178 589190
rect 43115 588164 43181 588165
rect 43115 588100 43116 588164
rect 43180 588100 43181 588164
rect 43115 588099 43181 588100
rect 25514 586718 25546 586954
rect 25782 586718 25866 586954
rect 26102 586718 26134 586954
rect 25514 566954 26134 586718
rect 25514 566718 25546 566954
rect 25782 566718 25866 566954
rect 26102 566718 26134 566954
rect 25514 546954 26134 566718
rect 29234 570614 29854 588000
rect 29234 570378 29266 570614
rect 29502 570378 29586 570614
rect 29822 570378 29854 570614
rect 29234 563308 29854 570378
rect 31794 573294 32414 588000
rect 31794 573058 31826 573294
rect 32062 573058 32146 573294
rect 32382 573058 32414 573294
rect 31794 563308 32414 573058
rect 32954 574274 33574 588000
rect 32954 574038 32986 574274
rect 33222 574038 33306 574274
rect 33542 574038 33574 574274
rect 32954 563308 33574 574038
rect 35514 576954 36134 588000
rect 35514 576718 35546 576954
rect 35782 576718 35866 576954
rect 36102 576718 36134 576954
rect 35514 563308 36134 576718
rect 39234 580614 39854 588000
rect 39234 580378 39266 580614
rect 39502 580378 39586 580614
rect 39822 580378 39854 580614
rect 39234 563308 39854 580378
rect 41794 583294 42414 588000
rect 41794 583058 41826 583294
rect 42062 583058 42146 583294
rect 42382 583058 42414 583294
rect 41794 563308 42414 583058
rect 42954 584274 43574 588000
rect 43670 587893 43730 589190
rect 60598 589230 60668 589290
rect 63174 589230 63252 589290
rect 64646 589230 65700 589290
rect 68088 589290 68148 590106
rect 70672 589290 70732 590106
rect 73120 589290 73180 590106
rect 68088 589230 68202 589290
rect 70672 589230 70778 589290
rect 43667 587892 43733 587893
rect 43667 587828 43668 587892
rect 43732 587828 43733 587892
rect 43667 587827 43733 587828
rect 42954 584038 42986 584274
rect 43222 584038 43306 584274
rect 43542 584038 43574 584274
rect 42954 564274 43574 584038
rect 42954 564038 42986 564274
rect 43222 564038 43306 564274
rect 43542 564038 43574 564274
rect 42954 563308 43574 564038
rect 45514 586954 46134 588000
rect 45514 586718 45546 586954
rect 45782 586718 45866 586954
rect 46102 586718 46134 586954
rect 45514 566954 46134 586718
rect 45514 566718 45546 566954
rect 45782 566718 45866 566954
rect 46102 566718 46134 566954
rect 45514 563308 46134 566718
rect 49234 570614 49854 588000
rect 49234 570378 49266 570614
rect 49502 570378 49586 570614
rect 49822 570378 49854 570614
rect 49234 563308 49854 570378
rect 51794 573294 52414 588000
rect 51794 573058 51826 573294
rect 52062 573058 52146 573294
rect 52382 573058 52414 573294
rect 51794 563308 52414 573058
rect 52954 574274 53574 588000
rect 52954 574038 52986 574274
rect 53222 574038 53306 574274
rect 53542 574038 53574 574274
rect 52954 563308 53574 574038
rect 55514 576954 56134 588000
rect 55514 576718 55546 576954
rect 55782 576718 55866 576954
rect 56102 576718 56134 576954
rect 55514 563308 56134 576718
rect 59234 580614 59854 588000
rect 60598 587893 60658 589230
rect 63174 588165 63234 589230
rect 63171 588164 63237 588165
rect 63171 588100 63172 588164
rect 63236 588100 63237 588164
rect 63171 588099 63237 588100
rect 60595 587892 60661 587893
rect 60595 587828 60596 587892
rect 60660 587828 60661 587892
rect 60595 587827 60661 587828
rect 59234 580378 59266 580614
rect 59502 580378 59586 580614
rect 59822 580378 59854 580614
rect 59234 563308 59854 580378
rect 61794 583294 62414 588000
rect 61794 583058 61826 583294
rect 62062 583058 62146 583294
rect 62382 583058 62414 583294
rect 61794 563308 62414 583058
rect 62954 584274 63574 588000
rect 64646 586530 64706 589230
rect 65514 586954 66134 588000
rect 68142 587893 68202 589230
rect 68139 587892 68205 587893
rect 68139 587828 68140 587892
rect 68204 587828 68205 587892
rect 68139 587827 68205 587828
rect 65514 586718 65546 586954
rect 65782 586718 65866 586954
rect 66102 586718 66134 586954
rect 64827 586532 64893 586533
rect 64827 586530 64828 586532
rect 64646 586470 64828 586530
rect 64827 586468 64828 586470
rect 64892 586468 64893 586532
rect 64827 586467 64893 586468
rect 62954 584038 62986 584274
rect 63222 584038 63306 584274
rect 63542 584038 63574 584274
rect 62954 564274 63574 584038
rect 62954 564038 62986 564274
rect 63222 564038 63306 564274
rect 63542 564038 63574 564274
rect 62954 563308 63574 564038
rect 65514 566954 66134 586718
rect 65514 566718 65546 566954
rect 65782 566718 65866 566954
rect 66102 566718 66134 566954
rect 65514 563308 66134 566718
rect 69234 570614 69854 588000
rect 70718 586669 70778 589230
rect 73110 589230 73180 589290
rect 75568 589250 75628 590106
rect 73110 588165 73170 589230
rect 75318 589190 75628 589250
rect 78016 589250 78076 590106
rect 80600 589250 80660 590106
rect 83048 589250 83108 590106
rect 85632 589250 85692 590106
rect 78016 589190 78138 589250
rect 80600 589190 80714 589250
rect 73107 588164 73173 588165
rect 73107 588100 73108 588164
rect 73172 588100 73173 588164
rect 73107 588099 73173 588100
rect 70715 586668 70781 586669
rect 70715 586604 70716 586668
rect 70780 586604 70781 586668
rect 70715 586603 70781 586604
rect 69234 570378 69266 570614
rect 69502 570378 69586 570614
rect 69822 570378 69854 570614
rect 69234 563308 69854 570378
rect 71794 573294 72414 588000
rect 71794 573058 71826 573294
rect 72062 573058 72146 573294
rect 72382 573058 72414 573294
rect 71794 563308 72414 573058
rect 72954 574274 73574 588000
rect 75318 586669 75378 589190
rect 75315 586668 75381 586669
rect 75315 586604 75316 586668
rect 75380 586604 75381 586668
rect 75315 586603 75381 586604
rect 72954 574038 72986 574274
rect 73222 574038 73306 574274
rect 73542 574038 73574 574274
rect 72954 563308 73574 574038
rect 75514 576954 76134 588000
rect 78078 586669 78138 589190
rect 78075 586668 78141 586669
rect 78075 586604 78076 586668
rect 78140 586604 78141 586668
rect 78075 586603 78141 586604
rect 75514 576718 75546 576954
rect 75782 576718 75866 576954
rect 76102 576718 76134 576954
rect 75514 563308 76134 576718
rect 79234 580614 79854 588000
rect 80654 586669 80714 589190
rect 83046 589190 83108 589250
rect 85622 589190 85692 589250
rect 88080 589250 88140 590106
rect 90664 589250 90724 590106
rect 93112 589250 93172 590106
rect 95560 589250 95620 590106
rect 88080 589190 88258 589250
rect 83046 588165 83106 589190
rect 85622 588165 85682 589190
rect 83043 588164 83109 588165
rect 83043 588100 83044 588164
rect 83108 588100 83109 588164
rect 83043 588099 83109 588100
rect 85619 588164 85685 588165
rect 85619 588100 85620 588164
rect 85684 588100 85685 588164
rect 85619 588099 85685 588100
rect 80651 586668 80717 586669
rect 80651 586604 80652 586668
rect 80716 586604 80717 586668
rect 80651 586603 80717 586604
rect 79234 580378 79266 580614
rect 79502 580378 79586 580614
rect 79822 580378 79854 580614
rect 79234 563308 79854 580378
rect 81794 583294 82414 588000
rect 81794 583058 81826 583294
rect 82062 583058 82146 583294
rect 82382 583058 82414 583294
rect 81794 563308 82414 583058
rect 82954 584274 83574 588000
rect 82954 584038 82986 584274
rect 83222 584038 83306 584274
rect 83542 584038 83574 584274
rect 82954 564274 83574 584038
rect 82954 564038 82986 564274
rect 83222 564038 83306 564274
rect 83542 564038 83574 564274
rect 82954 563308 83574 564038
rect 85514 586954 86134 588000
rect 88198 587893 88258 589190
rect 90590 589190 90724 589250
rect 92798 589190 93172 589250
rect 95558 589190 95620 589250
rect 98280 589250 98340 590106
rect 100592 589250 100652 590106
rect 98280 589190 98378 589250
rect 88195 587892 88261 587893
rect 88195 587828 88196 587892
rect 88260 587828 88261 587892
rect 88195 587827 88261 587828
rect 85514 586718 85546 586954
rect 85782 586718 85866 586954
rect 86102 586718 86134 586954
rect 85514 566954 86134 586718
rect 85514 566718 85546 566954
rect 85782 566718 85866 566954
rect 86102 566718 86134 566954
rect 85514 563308 86134 566718
rect 89234 570614 89854 588000
rect 90590 586669 90650 589190
rect 90587 586668 90653 586669
rect 90587 586604 90588 586668
rect 90652 586604 90653 586668
rect 90587 586603 90653 586604
rect 89234 570378 89266 570614
rect 89502 570378 89586 570614
rect 89822 570378 89854 570614
rect 89234 563308 89854 570378
rect 91794 573294 92414 588000
rect 92798 586669 92858 589190
rect 95558 588165 95618 589190
rect 95555 588164 95621 588165
rect 95555 588100 95556 588164
rect 95620 588100 95621 588164
rect 95555 588099 95621 588100
rect 92795 586668 92861 586669
rect 92795 586604 92796 586668
rect 92860 586604 92861 586668
rect 92795 586603 92861 586604
rect 91794 573058 91826 573294
rect 92062 573058 92146 573294
rect 92382 573058 92414 573294
rect 91794 563308 92414 573058
rect 92954 574274 93574 588000
rect 92954 574038 92986 574274
rect 93222 574038 93306 574274
rect 93542 574038 93574 574274
rect 92954 563308 93574 574038
rect 95514 576954 96134 588000
rect 98318 587893 98378 589190
rect 100526 589190 100652 589250
rect 103040 589250 103100 590106
rect 105624 589290 105684 590106
rect 107392 589290 107452 590106
rect 108072 589290 108132 590106
rect 108480 589290 108540 590106
rect 109568 589290 109628 590106
rect 110520 589290 110580 590106
rect 103040 589190 103162 589250
rect 98315 587892 98381 587893
rect 98315 587828 98316 587892
rect 98380 587828 98381 587892
rect 98315 587827 98381 587828
rect 95514 576718 95546 576954
rect 95782 576718 95866 576954
rect 96102 576718 96134 576954
rect 95514 563308 96134 576718
rect 99234 580614 99854 588000
rect 100526 587893 100586 589190
rect 103102 588165 103162 589190
rect 105310 589230 105684 589290
rect 107334 589230 107452 589290
rect 108070 589230 108132 589290
rect 108438 589230 108540 589290
rect 109542 589230 109628 589290
rect 110462 589230 110580 589290
rect 110792 589290 110852 590106
rect 112152 589290 112212 590106
rect 110792 589230 110890 589290
rect 103099 588164 103165 588165
rect 103099 588100 103100 588164
rect 103164 588100 103165 588164
rect 103099 588099 103165 588100
rect 100523 587892 100589 587893
rect 100523 587828 100524 587892
rect 100588 587828 100589 587892
rect 100523 587827 100589 587828
rect 99234 580378 99266 580614
rect 99502 580378 99586 580614
rect 99822 580378 99854 580614
rect 99234 563308 99854 580378
rect 101794 583294 102414 588000
rect 101794 583058 101826 583294
rect 102062 583058 102146 583294
rect 102382 583058 102414 583294
rect 101794 563308 102414 583058
rect 102954 584274 103574 588000
rect 105310 587893 105370 589230
rect 105307 587892 105373 587893
rect 105307 587828 105308 587892
rect 105372 587828 105373 587892
rect 105307 587827 105373 587828
rect 102954 584038 102986 584274
rect 103222 584038 103306 584274
rect 103542 584038 103574 584274
rect 102954 564274 103574 584038
rect 102954 564038 102986 564274
rect 103222 564038 103306 564274
rect 103542 564038 103574 564274
rect 102954 563308 103574 564038
rect 105514 586954 106134 588000
rect 107334 587893 107394 589230
rect 107331 587892 107397 587893
rect 107331 587828 107332 587892
rect 107396 587828 107397 587892
rect 107331 587827 107397 587828
rect 105514 586718 105546 586954
rect 105782 586718 105866 586954
rect 106102 586718 106134 586954
rect 105514 566954 106134 586718
rect 108070 586669 108130 589230
rect 108438 587893 108498 589230
rect 109542 588165 109602 589230
rect 109539 588164 109605 588165
rect 109539 588100 109540 588164
rect 109604 588100 109605 588164
rect 109539 588099 109605 588100
rect 108435 587892 108501 587893
rect 108435 587828 108436 587892
rect 108500 587828 108501 587892
rect 108435 587827 108501 587828
rect 108067 586668 108133 586669
rect 108067 586604 108068 586668
rect 108132 586604 108133 586668
rect 108067 586603 108133 586604
rect 105514 566718 105546 566954
rect 105782 566718 105866 566954
rect 106102 566718 106134 566954
rect 105514 563308 106134 566718
rect 109234 570614 109854 588000
rect 110462 587893 110522 589230
rect 110830 587893 110890 589230
rect 112118 589230 112212 589290
rect 112968 589290 113028 590106
rect 113240 589290 113300 590106
rect 114328 589290 114388 590106
rect 115416 589290 115476 590106
rect 112968 589230 113098 589290
rect 113240 589230 113834 589290
rect 112118 588165 112178 589230
rect 113038 588165 113098 589230
rect 112115 588164 112181 588165
rect 112115 588100 112116 588164
rect 112180 588100 112181 588164
rect 112115 588099 112181 588100
rect 113035 588164 113101 588165
rect 113035 588100 113036 588164
rect 113100 588100 113101 588164
rect 113035 588099 113101 588100
rect 110459 587892 110525 587893
rect 110459 587828 110460 587892
rect 110524 587828 110525 587892
rect 110459 587827 110525 587828
rect 110827 587892 110893 587893
rect 110827 587828 110828 587892
rect 110892 587828 110893 587892
rect 110827 587827 110893 587828
rect 109234 570378 109266 570614
rect 109502 570378 109586 570614
rect 109822 570378 109854 570614
rect 109234 563308 109854 570378
rect 111794 573294 112414 588000
rect 111794 573058 111826 573294
rect 112062 573058 112146 573294
rect 112382 573058 112414 573294
rect 111794 563308 112414 573058
rect 112954 574274 113574 588000
rect 113774 587757 113834 589230
rect 114326 589230 114388 589290
rect 115246 589230 115476 589290
rect 115552 589290 115612 590106
rect 116776 589290 116836 590106
rect 117864 589290 117924 590106
rect 118272 589290 118332 590106
rect 118952 589290 119012 590106
rect 115552 589230 115674 589290
rect 114326 587893 114386 589230
rect 115246 587893 115306 589230
rect 115614 588165 115674 589230
rect 116718 589230 116836 589290
rect 117822 589230 117924 589290
rect 118190 589230 118332 589290
rect 118926 589230 119012 589290
rect 120176 589290 120236 590106
rect 120584 589290 120644 590106
rect 120176 589230 120274 589290
rect 115611 588164 115677 588165
rect 115611 588100 115612 588164
rect 115676 588100 115677 588164
rect 115611 588099 115677 588100
rect 114323 587892 114389 587893
rect 114323 587828 114324 587892
rect 114388 587828 114389 587892
rect 114323 587827 114389 587828
rect 115243 587892 115309 587893
rect 115243 587828 115244 587892
rect 115308 587828 115309 587892
rect 115243 587827 115309 587828
rect 113771 587756 113837 587757
rect 113771 587692 113772 587756
rect 113836 587692 113837 587756
rect 113771 587691 113837 587692
rect 112954 574038 112986 574274
rect 113222 574038 113306 574274
rect 113542 574038 113574 574274
rect 112954 563308 113574 574038
rect 115514 576954 116134 588000
rect 116718 587893 116778 589230
rect 116715 587892 116781 587893
rect 116715 587828 116716 587892
rect 116780 587828 116781 587892
rect 116715 587827 116781 587828
rect 117822 587077 117882 589230
rect 117819 587076 117885 587077
rect 117819 587012 117820 587076
rect 117884 587012 117885 587076
rect 117819 587011 117885 587012
rect 118190 586669 118250 589230
rect 118926 587893 118986 589230
rect 118923 587892 118989 587893
rect 118923 587828 118924 587892
rect 118988 587828 118989 587892
rect 118923 587827 118989 587828
rect 118187 586668 118253 586669
rect 118187 586604 118188 586668
rect 118252 586604 118253 586668
rect 118187 586603 118253 586604
rect 115514 576718 115546 576954
rect 115782 576718 115866 576954
rect 116102 576718 116134 576954
rect 115514 563308 116134 576718
rect 119234 580614 119854 588000
rect 120214 587893 120274 589230
rect 120582 589230 120644 589290
rect 121264 589290 121324 590106
rect 122624 589290 122684 590106
rect 123032 589290 123092 590106
rect 123712 589290 123772 590106
rect 121264 589230 121378 589290
rect 120211 587892 120277 587893
rect 120211 587828 120212 587892
rect 120276 587828 120277 587892
rect 120211 587827 120277 587828
rect 120582 587757 120642 589230
rect 121318 587893 121378 589230
rect 122606 589230 122684 589290
rect 122974 589230 123092 589290
rect 123710 589230 123772 589290
rect 124800 589290 124860 590106
rect 125480 589290 125540 590106
rect 124800 589230 124874 589290
rect 121315 587892 121381 587893
rect 121315 587828 121316 587892
rect 121380 587828 121381 587892
rect 121315 587827 121381 587828
rect 120579 587756 120645 587757
rect 120579 587692 120580 587756
rect 120644 587692 120645 587756
rect 120579 587691 120645 587692
rect 119234 580378 119266 580614
rect 119502 580378 119586 580614
rect 119822 580378 119854 580614
rect 119234 563308 119854 580378
rect 121794 583294 122414 588000
rect 122606 587893 122666 589230
rect 122974 588165 123034 589230
rect 122971 588164 123037 588165
rect 122971 588100 122972 588164
rect 123036 588100 123037 588164
rect 122971 588099 123037 588100
rect 122603 587892 122669 587893
rect 122603 587828 122604 587892
rect 122668 587828 122669 587892
rect 122603 587827 122669 587828
rect 121794 583058 121826 583294
rect 122062 583058 122146 583294
rect 122382 583058 122414 583294
rect 121794 563308 122414 583058
rect 122954 584274 123574 588000
rect 123710 587349 123770 589230
rect 124814 587893 124874 589230
rect 125366 589230 125540 589290
rect 125888 589290 125948 590106
rect 127112 589290 127172 590106
rect 128064 589290 128124 590106
rect 128472 589290 128532 590106
rect 129560 589290 129620 590106
rect 130512 589290 130572 590106
rect 130648 589290 130708 590106
rect 132008 589290 132068 590106
rect 132960 589290 133020 590106
rect 133096 589290 133156 590106
rect 125888 589230 126346 589290
rect 127112 589230 127266 589290
rect 128064 589230 128186 589290
rect 128472 589230 128554 589290
rect 129560 589230 129658 589290
rect 130512 589230 130578 589290
rect 130648 589230 130762 589290
rect 124811 587892 124877 587893
rect 124811 587828 124812 587892
rect 124876 587828 124877 587892
rect 124811 587827 124877 587828
rect 123707 587348 123773 587349
rect 123707 587284 123708 587348
rect 123772 587284 123773 587348
rect 123707 587283 123773 587284
rect 125366 586669 125426 589230
rect 125514 586954 126134 588000
rect 126286 587893 126346 589230
rect 126283 587892 126349 587893
rect 126283 587828 126284 587892
rect 126348 587828 126349 587892
rect 126283 587827 126349 587828
rect 127206 587485 127266 589230
rect 127203 587484 127269 587485
rect 127203 587420 127204 587484
rect 127268 587420 127269 587484
rect 127203 587419 127269 587420
rect 125514 586718 125546 586954
rect 125782 586718 125866 586954
rect 126102 586718 126134 586954
rect 125363 586668 125429 586669
rect 125363 586604 125364 586668
rect 125428 586604 125429 586668
rect 125363 586603 125429 586604
rect 122954 584038 122986 584274
rect 123222 584038 123306 584274
rect 123542 584038 123574 584274
rect 122954 564274 123574 584038
rect 122954 564038 122986 564274
rect 123222 564038 123306 564274
rect 123542 564038 123574 564274
rect 122954 563308 123574 564038
rect 125514 566954 126134 586718
rect 128126 586669 128186 589230
rect 128494 587893 128554 589230
rect 129598 588165 129658 589230
rect 129595 588164 129661 588165
rect 129595 588100 129596 588164
rect 129660 588100 129661 588164
rect 129595 588099 129661 588100
rect 128491 587892 128557 587893
rect 128491 587828 128492 587892
rect 128556 587828 128557 587892
rect 128491 587827 128557 587828
rect 128123 586668 128189 586669
rect 128123 586604 128124 586668
rect 128188 586604 128189 586668
rect 128123 586603 128189 586604
rect 125514 566718 125546 566954
rect 125782 566718 125866 566954
rect 126102 566718 126134 566954
rect 125514 563308 126134 566718
rect 129234 570614 129854 588000
rect 130518 587757 130578 589230
rect 130702 587893 130762 589230
rect 131622 589230 132068 589290
rect 132726 589230 133020 589290
rect 133094 589230 133156 589290
rect 134184 589290 134244 590106
rect 135272 589290 135332 590106
rect 135816 589290 135876 590106
rect 136496 589290 136556 590106
rect 137856 589290 137916 590106
rect 138264 589290 138324 590106
rect 134184 589230 134258 589290
rect 135272 589230 135362 589290
rect 135816 589230 136282 589290
rect 136496 589230 136650 589290
rect 137856 589230 137938 589290
rect 131622 587893 131682 589230
rect 130699 587892 130765 587893
rect 130699 587828 130700 587892
rect 130764 587828 130765 587892
rect 130699 587827 130765 587828
rect 131619 587892 131685 587893
rect 131619 587828 131620 587892
rect 131684 587828 131685 587892
rect 131619 587827 131685 587828
rect 130515 587756 130581 587757
rect 130515 587692 130516 587756
rect 130580 587692 130581 587756
rect 130515 587691 130581 587692
rect 129234 570378 129266 570614
rect 129502 570378 129586 570614
rect 129822 570378 129854 570614
rect 129234 563308 129854 570378
rect 131794 573294 132414 588000
rect 132726 587893 132786 589230
rect 133094 588165 133154 589230
rect 133091 588164 133157 588165
rect 133091 588100 133092 588164
rect 133156 588100 133157 588164
rect 133091 588099 133157 588100
rect 132723 587892 132789 587893
rect 132723 587828 132724 587892
rect 132788 587828 132789 587892
rect 132723 587827 132789 587828
rect 131794 573058 131826 573294
rect 132062 573058 132146 573294
rect 132382 573058 132414 573294
rect 131794 563308 132414 573058
rect 132954 574274 133574 588000
rect 134198 587757 134258 589230
rect 134195 587756 134261 587757
rect 134195 587692 134196 587756
rect 134260 587692 134261 587756
rect 134195 587691 134261 587692
rect 135302 587621 135362 589230
rect 135299 587620 135365 587621
rect 135299 587556 135300 587620
rect 135364 587556 135365 587620
rect 135299 587555 135365 587556
rect 132954 574038 132986 574274
rect 133222 574038 133306 574274
rect 133542 574038 133574 574274
rect 132954 563308 133574 574038
rect 135514 576954 136134 588000
rect 136222 587893 136282 589230
rect 136219 587892 136285 587893
rect 136219 587828 136220 587892
rect 136284 587828 136285 587892
rect 136219 587827 136285 587828
rect 136590 587077 136650 589230
rect 137878 587893 137938 589230
rect 138246 589230 138324 589290
rect 138944 589290 139004 590106
rect 140032 589290 140092 590106
rect 141120 589290 141180 590106
rect 138944 589230 139042 589290
rect 140032 589230 140146 589290
rect 138246 587893 138306 589230
rect 137875 587892 137941 587893
rect 137875 587828 137876 587892
rect 137940 587828 137941 587892
rect 137875 587827 137941 587828
rect 138243 587892 138309 587893
rect 138243 587828 138244 587892
rect 138308 587828 138309 587892
rect 138243 587827 138309 587828
rect 138982 587077 139042 589230
rect 136587 587076 136653 587077
rect 136587 587012 136588 587076
rect 136652 587012 136653 587076
rect 136587 587011 136653 587012
rect 138979 587076 139045 587077
rect 138979 587012 138980 587076
rect 139044 587012 139045 587076
rect 138979 587011 139045 587012
rect 135514 576718 135546 576954
rect 135782 576718 135866 576954
rect 136102 576718 136134 576954
rect 135514 563308 136134 576718
rect 139234 580614 139854 588000
rect 140086 587893 140146 589230
rect 141006 589230 141180 589290
rect 142344 589250 142404 590106
rect 143432 589250 143492 590106
rect 144792 589797 144852 590106
rect 146016 589797 146076 590106
rect 144789 589796 144855 589797
rect 144789 589732 144790 589796
rect 144854 589732 144855 589796
rect 144789 589731 144855 589732
rect 146013 589796 146079 589797
rect 146013 589732 146014 589796
rect 146078 589732 146079 589796
rect 146013 589731 146079 589732
rect 140083 587892 140149 587893
rect 140083 587828 140084 587892
rect 140148 587828 140149 587892
rect 140083 587827 140149 587828
rect 141006 586669 141066 589230
rect 142344 589190 142722 589250
rect 141003 586668 141069 586669
rect 141003 586604 141004 586668
rect 141068 586604 141069 586668
rect 141003 586603 141069 586604
rect 139234 580378 139266 580614
rect 139502 580378 139586 580614
rect 139822 580378 139854 580614
rect 139234 563308 139854 580378
rect 141794 583294 142414 588000
rect 142662 587893 142722 589190
rect 143398 589190 143492 589250
rect 146016 589250 146076 589731
rect 146968 589250 147028 590106
rect 148328 589250 148388 590106
rect 149416 589250 149476 590106
rect 150504 589250 150564 590106
rect 146016 589190 147138 589250
rect 148328 589190 148426 589250
rect 149416 589190 149530 589250
rect 150504 589190 150634 589250
rect 143398 588165 143458 589190
rect 143395 588164 143461 588165
rect 143395 588100 143396 588164
rect 143460 588100 143461 588164
rect 143395 588099 143461 588100
rect 142659 587892 142725 587893
rect 142659 587828 142660 587892
rect 142724 587828 142725 587892
rect 142659 587827 142725 587828
rect 141794 583058 141826 583294
rect 142062 583058 142146 583294
rect 142382 583058 142414 583294
rect 141794 563308 142414 583058
rect 142954 584274 143574 588000
rect 142954 584038 142986 584274
rect 143222 584038 143306 584274
rect 143542 584038 143574 584274
rect 142954 564274 143574 584038
rect 142954 564038 142986 564274
rect 143222 564038 143306 564274
rect 143542 564038 143574 564274
rect 142954 563308 143574 564038
rect 145514 586954 146134 588000
rect 147078 587893 147138 589190
rect 148366 587893 148426 589190
rect 149470 588165 149530 589190
rect 149467 588164 149533 588165
rect 149467 588100 149468 588164
rect 149532 588100 149533 588164
rect 149467 588099 149533 588100
rect 147075 587892 147141 587893
rect 147075 587828 147076 587892
rect 147140 587828 147141 587892
rect 147075 587827 147141 587828
rect 148363 587892 148429 587893
rect 148363 587828 148364 587892
rect 148428 587828 148429 587892
rect 148363 587827 148429 587828
rect 145514 586718 145546 586954
rect 145782 586718 145866 586954
rect 146102 586718 146134 586954
rect 145514 566954 146134 586718
rect 145514 566718 145546 566954
rect 145782 566718 145866 566954
rect 146102 566718 146134 566954
rect 145514 563308 146134 566718
rect 149234 570614 149854 588000
rect 150574 587893 150634 589190
rect 150571 587892 150637 587893
rect 150571 587828 150572 587892
rect 150636 587828 150637 587892
rect 150571 587827 150637 587828
rect 149234 570378 149266 570614
rect 149502 570378 149586 570614
rect 149822 570378 149854 570614
rect 149234 563308 149854 570378
rect 151794 573294 152414 588000
rect 151794 573058 151826 573294
rect 152062 573058 152146 573294
rect 152382 573058 152414 573294
rect 151794 563308 152414 573058
rect 152954 574274 153574 588000
rect 152954 574038 152986 574274
rect 153222 574038 153306 574274
rect 153542 574038 153574 574274
rect 152954 563308 153574 574038
rect 155514 576954 156134 588000
rect 155514 576718 155546 576954
rect 155782 576718 155866 576954
rect 156102 576718 156134 576954
rect 155514 563308 156134 576718
rect 159234 580614 159854 588000
rect 159234 580378 159266 580614
rect 159502 580378 159586 580614
rect 159822 580378 159854 580614
rect 159234 563308 159854 580378
rect 161794 583294 162414 588000
rect 161794 583058 161826 583294
rect 162062 583058 162146 583294
rect 162382 583058 162414 583294
rect 161794 563308 162414 583058
rect 162954 584274 163574 588000
rect 162954 584038 162986 584274
rect 163222 584038 163306 584274
rect 163542 584038 163574 584274
rect 162954 564274 163574 584038
rect 162954 564038 162986 564274
rect 163222 564038 163306 564274
rect 163542 564038 163574 564274
rect 162954 563308 163574 564038
rect 165514 586954 166134 588000
rect 166947 587756 167013 587757
rect 166947 587692 166948 587756
rect 167012 587692 167013 587756
rect 166947 587691 167013 587692
rect 165514 586718 165546 586954
rect 165782 586718 165866 586954
rect 166102 586718 166134 586954
rect 165514 566954 166134 586718
rect 165514 566718 165546 566954
rect 165782 566718 165866 566954
rect 166102 566718 166134 566954
rect 165514 563308 166134 566718
rect 35755 563140 35821 563141
rect 35755 563076 35756 563140
rect 35820 563076 35821 563140
rect 35755 563075 35821 563076
rect 46795 563140 46861 563141
rect 46795 563076 46796 563140
rect 46860 563076 46861 563140
rect 46795 563075 46861 563076
rect 35758 562050 35818 563075
rect 35720 561990 35818 562050
rect 46798 562050 46858 563075
rect 46798 561990 46932 562050
rect 35720 561202 35780 561990
rect 46872 561202 46932 561990
rect 48093 561780 48159 561781
rect 48093 561716 48094 561780
rect 48158 561716 48159 561780
rect 48093 561715 48159 561716
rect 48096 561202 48156 561715
rect 30272 553294 30620 553456
rect 30272 553058 30328 553294
rect 30564 553058 30620 553294
rect 30272 552896 30620 553058
rect 166000 553294 166348 553456
rect 166000 553058 166056 553294
rect 166292 553058 166348 553294
rect 166000 552896 166348 553058
rect 25514 546718 25546 546954
rect 25782 546718 25866 546954
rect 26102 546718 26134 546954
rect 25514 526954 26134 546718
rect 30952 543294 31300 543456
rect 30952 543058 31008 543294
rect 31244 543058 31300 543294
rect 30952 542896 31300 543058
rect 165320 543294 165668 543456
rect 165320 543058 165376 543294
rect 165612 543058 165668 543294
rect 165320 542896 165668 543058
rect 30272 533294 30620 533456
rect 30272 533058 30328 533294
rect 30564 533058 30620 533294
rect 30272 532896 30620 533058
rect 166000 533294 166348 533456
rect 166000 533058 166056 533294
rect 166292 533058 166348 533294
rect 166000 532896 166348 533058
rect 25514 526718 25546 526954
rect 25782 526718 25866 526954
rect 26102 526718 26134 526954
rect 25514 506954 26134 526718
rect 30952 523294 31300 523456
rect 30952 523058 31008 523294
rect 31244 523058 31300 523294
rect 30952 522896 31300 523058
rect 165320 523294 165668 523456
rect 165320 523058 165376 523294
rect 165612 523058 165668 523294
rect 165320 522896 165668 523058
rect 30272 513294 30620 513456
rect 30272 513058 30328 513294
rect 30564 513058 30620 513294
rect 30272 512896 30620 513058
rect 166000 513294 166348 513456
rect 166000 513058 166056 513294
rect 166292 513058 166348 513294
rect 166000 512896 166348 513058
rect 25514 506718 25546 506954
rect 25782 506718 25866 506954
rect 26102 506718 26134 506954
rect 25514 486954 26134 506718
rect 30952 503294 31300 503456
rect 30952 503058 31008 503294
rect 31244 503058 31300 503294
rect 30952 502896 31300 503058
rect 165320 503294 165668 503456
rect 165320 503058 165376 503294
rect 165612 503058 165668 503294
rect 165320 502896 165668 503058
rect 30272 493294 30620 493456
rect 30272 493058 30328 493294
rect 30564 493058 30620 493294
rect 30272 492896 30620 493058
rect 166000 493294 166348 493456
rect 166000 493058 166056 493294
rect 166292 493058 166348 493294
rect 166000 492896 166348 493058
rect 25514 486718 25546 486954
rect 25782 486718 25866 486954
rect 26102 486718 26134 486954
rect 25514 466954 26134 486718
rect 30952 483294 31300 483456
rect 30952 483058 31008 483294
rect 31244 483058 31300 483294
rect 30952 482896 31300 483058
rect 165320 483294 165668 483456
rect 165320 483058 165376 483294
rect 165612 483058 165668 483294
rect 165320 482896 165668 483058
rect 43200 477730 43260 478040
rect 42750 477670 43260 477730
rect 43336 477730 43396 478040
rect 60608 477730 60668 478040
rect 63192 477730 63252 478040
rect 43336 477670 43730 477730
rect 25514 466718 25546 466954
rect 25782 466718 25866 466954
rect 26102 466718 26134 466954
rect 25514 446954 26134 466718
rect 29234 470614 29854 476000
rect 29234 470378 29266 470614
rect 29502 470378 29586 470614
rect 29822 470378 29854 470614
rect 29234 451308 29854 470378
rect 31794 473294 32414 476000
rect 31794 473058 31826 473294
rect 32062 473058 32146 473294
rect 32382 473058 32414 473294
rect 31794 453294 32414 473058
rect 31794 453058 31826 453294
rect 32062 453058 32146 453294
rect 32382 453058 32414 453294
rect 31794 451308 32414 453058
rect 32954 474274 33574 476000
rect 32954 474038 32986 474274
rect 33222 474038 33306 474274
rect 33542 474038 33574 474274
rect 32954 454274 33574 474038
rect 32954 454038 32986 454274
rect 33222 454038 33306 454274
rect 33542 454038 33574 454274
rect 32954 451308 33574 454038
rect 35514 456954 36134 476000
rect 35514 456718 35546 456954
rect 35782 456718 35866 456954
rect 36102 456718 36134 456954
rect 35203 452572 35269 452573
rect 35203 452508 35204 452572
rect 35268 452508 35269 452572
rect 35203 452507 35269 452508
rect 35206 449850 35266 452507
rect 35514 451308 36134 456718
rect 39234 460614 39854 476000
rect 39234 460378 39266 460614
rect 39502 460378 39586 460614
rect 39822 460378 39854 460614
rect 39234 451308 39854 460378
rect 41794 463294 42414 476000
rect 42750 475557 42810 477670
rect 42747 475556 42813 475557
rect 42747 475492 42748 475556
rect 42812 475492 42813 475556
rect 42747 475491 42813 475492
rect 41794 463058 41826 463294
rect 42062 463058 42146 463294
rect 42382 463058 42414 463294
rect 41794 451308 42414 463058
rect 42954 464274 43574 476000
rect 43670 475421 43730 477670
rect 60598 477670 60668 477730
rect 63174 477670 63252 477730
rect 65640 477730 65700 478040
rect 68088 477730 68148 478040
rect 70672 477730 70732 478040
rect 73120 477730 73180 478040
rect 75568 477730 75628 478040
rect 65640 477670 65810 477730
rect 68088 477670 68202 477730
rect 70672 477670 70778 477730
rect 73120 477670 73722 477730
rect 43667 475420 43733 475421
rect 43667 475356 43668 475420
rect 43732 475356 43733 475420
rect 43667 475355 43733 475356
rect 42954 464038 42986 464274
rect 43222 464038 43306 464274
rect 43542 464038 43574 464274
rect 42954 451308 43574 464038
rect 45514 466954 46134 476000
rect 45514 466718 45546 466954
rect 45782 466718 45866 466954
rect 46102 466718 46134 466954
rect 45514 451308 46134 466718
rect 49234 470614 49854 476000
rect 49234 470378 49266 470614
rect 49502 470378 49586 470614
rect 49822 470378 49854 470614
rect 46795 451892 46861 451893
rect 46795 451828 46796 451892
rect 46860 451828 46861 451892
rect 46795 451827 46861 451828
rect 46798 449850 46858 451827
rect 48083 451348 48149 451349
rect 48083 451284 48084 451348
rect 48148 451284 48149 451348
rect 49234 451308 49854 470378
rect 51794 473294 52414 476000
rect 51794 473058 51826 473294
rect 52062 473058 52146 473294
rect 52382 473058 52414 473294
rect 51794 453294 52414 473058
rect 51794 453058 51826 453294
rect 52062 453058 52146 453294
rect 52382 453058 52414 453294
rect 51794 451308 52414 453058
rect 52954 474274 53574 476000
rect 52954 474038 52986 474274
rect 53222 474038 53306 474274
rect 53542 474038 53574 474274
rect 52954 454274 53574 474038
rect 52954 454038 52986 454274
rect 53222 454038 53306 454274
rect 53542 454038 53574 454274
rect 52954 451308 53574 454038
rect 55514 456954 56134 476000
rect 55514 456718 55546 456954
rect 55782 456718 55866 456954
rect 56102 456718 56134 456954
rect 55514 451308 56134 456718
rect 59234 460614 59854 476000
rect 60598 474877 60658 477670
rect 63174 476237 63234 477670
rect 65750 476237 65810 477670
rect 63171 476236 63237 476237
rect 63171 476172 63172 476236
rect 63236 476172 63237 476236
rect 63171 476171 63237 476172
rect 65747 476236 65813 476237
rect 65747 476172 65748 476236
rect 65812 476172 65813 476236
rect 65747 476171 65813 476172
rect 60595 474876 60661 474877
rect 60595 474812 60596 474876
rect 60660 474812 60661 474876
rect 60595 474811 60661 474812
rect 59234 460378 59266 460614
rect 59502 460378 59586 460614
rect 59822 460378 59854 460614
rect 59234 451308 59854 460378
rect 61794 463294 62414 476000
rect 61794 463058 61826 463294
rect 62062 463058 62146 463294
rect 62382 463058 62414 463294
rect 61794 451308 62414 463058
rect 62954 464274 63574 476000
rect 62954 464038 62986 464274
rect 63222 464038 63306 464274
rect 63542 464038 63574 464274
rect 62954 451308 63574 464038
rect 65514 466954 66134 476000
rect 68142 474877 68202 477670
rect 68139 474876 68205 474877
rect 68139 474812 68140 474876
rect 68204 474812 68205 474876
rect 68139 474811 68205 474812
rect 65514 466718 65546 466954
rect 65782 466718 65866 466954
rect 66102 466718 66134 466954
rect 65514 451308 66134 466718
rect 69234 470614 69854 476000
rect 70718 474877 70778 477670
rect 70715 474876 70781 474877
rect 70715 474812 70716 474876
rect 70780 474812 70781 474876
rect 70715 474811 70781 474812
rect 69234 470378 69266 470614
rect 69502 470378 69586 470614
rect 69822 470378 69854 470614
rect 69234 451308 69854 470378
rect 71794 473294 72414 476000
rect 71794 473058 71826 473294
rect 72062 473058 72146 473294
rect 72382 473058 72414 473294
rect 71794 453294 72414 473058
rect 71794 453058 71826 453294
rect 72062 453058 72146 453294
rect 72382 453058 72414 453294
rect 71794 451308 72414 453058
rect 72954 474274 73574 476000
rect 73662 474877 73722 477670
rect 75318 477670 75628 477730
rect 78016 477730 78076 478040
rect 80600 477730 80660 478040
rect 83048 477730 83108 478040
rect 85632 477730 85692 478040
rect 78016 477670 78138 477730
rect 80600 477670 80714 477730
rect 75318 474877 75378 477670
rect 73659 474876 73725 474877
rect 73659 474812 73660 474876
rect 73724 474812 73725 474876
rect 73659 474811 73725 474812
rect 75315 474876 75381 474877
rect 75315 474812 75316 474876
rect 75380 474812 75381 474876
rect 75315 474811 75381 474812
rect 72954 474038 72986 474274
rect 73222 474038 73306 474274
rect 73542 474038 73574 474274
rect 72954 454274 73574 474038
rect 72954 454038 72986 454274
rect 73222 454038 73306 454274
rect 73542 454038 73574 454274
rect 72954 451308 73574 454038
rect 75514 456954 76134 476000
rect 78078 474877 78138 477670
rect 78075 474876 78141 474877
rect 78075 474812 78076 474876
rect 78140 474812 78141 474876
rect 78075 474811 78141 474812
rect 75514 456718 75546 456954
rect 75782 456718 75866 456954
rect 76102 456718 76134 456954
rect 75514 451308 76134 456718
rect 79234 460614 79854 476000
rect 80654 474877 80714 477670
rect 83046 477670 83108 477730
rect 85622 477670 85692 477730
rect 88080 477730 88140 478040
rect 90664 477730 90724 478040
rect 93112 477730 93172 478040
rect 95560 477730 95620 478040
rect 88080 477670 88258 477730
rect 90664 477670 90834 477730
rect 93112 477670 93778 477730
rect 83046 476237 83106 477670
rect 85622 476237 85682 477670
rect 83043 476236 83109 476237
rect 83043 476172 83044 476236
rect 83108 476172 83109 476236
rect 83043 476171 83109 476172
rect 85619 476236 85685 476237
rect 85619 476172 85620 476236
rect 85684 476172 85685 476236
rect 85619 476171 85685 476172
rect 80651 474876 80717 474877
rect 80651 474812 80652 474876
rect 80716 474812 80717 474876
rect 80651 474811 80717 474812
rect 79234 460378 79266 460614
rect 79502 460378 79586 460614
rect 79822 460378 79854 460614
rect 79234 451308 79854 460378
rect 81794 463294 82414 476000
rect 81794 463058 81826 463294
rect 82062 463058 82146 463294
rect 82382 463058 82414 463294
rect 81794 451308 82414 463058
rect 82954 464274 83574 476000
rect 82954 464038 82986 464274
rect 83222 464038 83306 464274
rect 83542 464038 83574 464274
rect 82954 451308 83574 464038
rect 85514 466954 86134 476000
rect 88198 474877 88258 477670
rect 88195 474876 88261 474877
rect 88195 474812 88196 474876
rect 88260 474812 88261 474876
rect 88195 474811 88261 474812
rect 85514 466718 85546 466954
rect 85782 466718 85866 466954
rect 86102 466718 86134 466954
rect 85514 451308 86134 466718
rect 89234 470614 89854 476000
rect 90774 474877 90834 477670
rect 90771 474876 90837 474877
rect 90771 474812 90772 474876
rect 90836 474812 90837 474876
rect 90771 474811 90837 474812
rect 89234 470378 89266 470614
rect 89502 470378 89586 470614
rect 89822 470378 89854 470614
rect 89234 451308 89854 470378
rect 91794 473294 92414 476000
rect 91794 473058 91826 473294
rect 92062 473058 92146 473294
rect 92382 473058 92414 473294
rect 91794 453294 92414 473058
rect 91794 453058 91826 453294
rect 92062 453058 92146 453294
rect 92382 453058 92414 453294
rect 91794 451308 92414 453058
rect 92954 474274 93574 476000
rect 93718 474877 93778 477670
rect 95374 477670 95620 477730
rect 98280 477730 98340 478040
rect 100592 477730 100652 478040
rect 103040 477730 103100 478040
rect 98280 477670 98378 477730
rect 95374 476101 95434 477670
rect 95371 476100 95437 476101
rect 95371 476036 95372 476100
rect 95436 476036 95437 476100
rect 95371 476035 95437 476036
rect 93715 474876 93781 474877
rect 93715 474812 93716 474876
rect 93780 474812 93781 474876
rect 93715 474811 93781 474812
rect 92954 474038 92986 474274
rect 93222 474038 93306 474274
rect 93542 474038 93574 474274
rect 92954 454274 93574 474038
rect 92954 454038 92986 454274
rect 93222 454038 93306 454274
rect 93542 454038 93574 454274
rect 92954 451308 93574 454038
rect 95514 456954 96134 476000
rect 98318 474877 98378 477670
rect 100526 477670 100652 477730
rect 102734 477670 103100 477730
rect 105624 477730 105684 478040
rect 107392 477730 107452 478040
rect 108072 477730 108132 478040
rect 108480 477730 108540 478040
rect 105624 477670 105738 477730
rect 98315 474876 98381 474877
rect 98315 474812 98316 474876
rect 98380 474812 98381 474876
rect 98315 474811 98381 474812
rect 95514 456718 95546 456954
rect 95782 456718 95866 456954
rect 96102 456718 96134 456954
rect 95514 451308 96134 456718
rect 99234 460614 99854 476000
rect 100526 474877 100586 477670
rect 100523 474876 100589 474877
rect 100523 474812 100524 474876
rect 100588 474812 100589 474876
rect 100523 474811 100589 474812
rect 99234 460378 99266 460614
rect 99502 460378 99586 460614
rect 99822 460378 99854 460614
rect 99234 451308 99854 460378
rect 101794 463294 102414 476000
rect 102734 474877 102794 477670
rect 105678 476237 105738 477670
rect 107334 477670 107452 477730
rect 108070 477670 108132 477730
rect 108438 477670 108540 477730
rect 109568 477730 109628 478040
rect 110520 477730 110580 478040
rect 109568 477670 110154 477730
rect 105675 476236 105741 476237
rect 105675 476172 105676 476236
rect 105740 476172 105741 476236
rect 105675 476171 105741 476172
rect 102731 474876 102797 474877
rect 102731 474812 102732 474876
rect 102796 474812 102797 474876
rect 102731 474811 102797 474812
rect 101794 463058 101826 463294
rect 102062 463058 102146 463294
rect 102382 463058 102414 463294
rect 101794 451308 102414 463058
rect 102954 464274 103574 476000
rect 102954 464038 102986 464274
rect 103222 464038 103306 464274
rect 103542 464038 103574 464274
rect 102954 451308 103574 464038
rect 105514 466954 106134 476000
rect 107334 474877 107394 477670
rect 108070 475013 108130 477670
rect 108067 475012 108133 475013
rect 108067 474948 108068 475012
rect 108132 474948 108133 475012
rect 108067 474947 108133 474948
rect 108438 474877 108498 477670
rect 107331 474876 107397 474877
rect 107331 474812 107332 474876
rect 107396 474812 107397 474876
rect 107331 474811 107397 474812
rect 108435 474876 108501 474877
rect 108435 474812 108436 474876
rect 108500 474812 108501 474876
rect 108435 474811 108501 474812
rect 105514 466718 105546 466954
rect 105782 466718 105866 466954
rect 106102 466718 106134 466954
rect 105514 451308 106134 466718
rect 109234 470614 109854 476000
rect 110094 475013 110154 477670
rect 110462 477670 110580 477730
rect 110792 477730 110852 478040
rect 112152 477730 112212 478040
rect 112968 477730 113028 478040
rect 113240 477730 113300 478040
rect 114328 477730 114388 478040
rect 115416 477869 115476 478040
rect 115413 477868 115479 477869
rect 115413 477804 115414 477868
rect 115478 477804 115479 477868
rect 115413 477803 115479 477804
rect 115552 477730 115612 478040
rect 116776 477730 116836 478040
rect 117864 477730 117924 478040
rect 110792 477670 110890 477730
rect 112152 477670 112730 477730
rect 112968 477670 113098 477730
rect 113240 477670 113834 477730
rect 110462 475013 110522 477670
rect 110091 475012 110157 475013
rect 110091 474948 110092 475012
rect 110156 474948 110157 475012
rect 110091 474947 110157 474948
rect 110459 475012 110525 475013
rect 110459 474948 110460 475012
rect 110524 474948 110525 475012
rect 110459 474947 110525 474948
rect 110830 474877 110890 477670
rect 110827 474876 110893 474877
rect 110827 474812 110828 474876
rect 110892 474812 110893 474876
rect 110827 474811 110893 474812
rect 109234 470378 109266 470614
rect 109502 470378 109586 470614
rect 109822 470378 109854 470614
rect 109234 451308 109854 470378
rect 111794 473294 112414 476000
rect 112670 474877 112730 477670
rect 113038 476237 113098 477670
rect 113035 476236 113101 476237
rect 113035 476172 113036 476236
rect 113100 476172 113101 476236
rect 113035 476171 113101 476172
rect 112667 474876 112733 474877
rect 112667 474812 112668 474876
rect 112732 474812 112733 474876
rect 112667 474811 112733 474812
rect 111794 473058 111826 473294
rect 112062 473058 112146 473294
rect 112382 473058 112414 473294
rect 111794 453294 112414 473058
rect 111794 453058 111826 453294
rect 112062 453058 112146 453294
rect 112382 453058 112414 453294
rect 111794 451308 112414 453058
rect 112954 474274 113574 476000
rect 113774 475013 113834 477670
rect 114326 477670 114388 477730
rect 115246 477670 115612 477730
rect 116718 477670 116836 477730
rect 117822 477670 117924 477730
rect 118272 477730 118332 478040
rect 118952 477730 119012 478040
rect 118272 477670 118434 477730
rect 113771 475012 113837 475013
rect 113771 474948 113772 475012
rect 113836 474948 113837 475012
rect 113771 474947 113837 474948
rect 114326 474877 114386 477670
rect 115246 474877 115306 477670
rect 114323 474876 114389 474877
rect 114323 474812 114324 474876
rect 114388 474812 114389 474876
rect 114323 474811 114389 474812
rect 115243 474876 115309 474877
rect 115243 474812 115244 474876
rect 115308 474812 115309 474876
rect 115243 474811 115309 474812
rect 112954 474038 112986 474274
rect 113222 474038 113306 474274
rect 113542 474038 113574 474274
rect 112954 454274 113574 474038
rect 112954 454038 112986 454274
rect 113222 454038 113306 454274
rect 113542 454038 113574 454274
rect 112954 451308 113574 454038
rect 115514 456954 116134 476000
rect 116718 474877 116778 477670
rect 117822 475013 117882 477670
rect 117819 475012 117885 475013
rect 117819 474948 117820 475012
rect 117884 474948 117885 475012
rect 117819 474947 117885 474948
rect 118374 474877 118434 477670
rect 118926 477670 119012 477730
rect 120176 477730 120236 478040
rect 120584 477730 120644 478040
rect 120176 477670 120274 477730
rect 118926 474877 118986 477670
rect 116715 474876 116781 474877
rect 116715 474812 116716 474876
rect 116780 474812 116781 474876
rect 116715 474811 116781 474812
rect 118371 474876 118437 474877
rect 118371 474812 118372 474876
rect 118436 474812 118437 474876
rect 118371 474811 118437 474812
rect 118923 474876 118989 474877
rect 118923 474812 118924 474876
rect 118988 474812 118989 474876
rect 118923 474811 118989 474812
rect 115514 456718 115546 456954
rect 115782 456718 115866 456954
rect 116102 456718 116134 456954
rect 115514 451308 116134 456718
rect 119234 460614 119854 476000
rect 120214 475557 120274 477670
rect 120582 477670 120644 477730
rect 121264 477730 121324 478040
rect 122624 477869 122684 478040
rect 122621 477868 122687 477869
rect 122621 477804 122622 477868
rect 122686 477804 122687 477868
rect 123032 477866 123092 478040
rect 122621 477803 122687 477804
rect 122974 477806 123092 477866
rect 122974 477730 123034 477806
rect 123712 477730 123772 478040
rect 121264 477670 121378 477730
rect 120211 475556 120277 475557
rect 120211 475492 120212 475556
rect 120276 475492 120277 475556
rect 120211 475491 120277 475492
rect 120582 474877 120642 477670
rect 121318 475013 121378 477670
rect 122606 477670 123034 477730
rect 123710 477670 123772 477730
rect 124800 477730 124860 478040
rect 125480 477730 125540 478040
rect 124800 477670 124874 477730
rect 121315 475012 121381 475013
rect 121315 474948 121316 475012
rect 121380 474948 121381 475012
rect 121315 474947 121381 474948
rect 120579 474876 120645 474877
rect 120579 474812 120580 474876
rect 120644 474812 120645 474876
rect 120579 474811 120645 474812
rect 119234 460378 119266 460614
rect 119502 460378 119586 460614
rect 119822 460378 119854 460614
rect 119234 451308 119854 460378
rect 121794 463294 122414 476000
rect 122606 475829 122666 477670
rect 122603 475828 122669 475829
rect 122603 475764 122604 475828
rect 122668 475764 122669 475828
rect 122603 475763 122669 475764
rect 121794 463058 121826 463294
rect 122062 463058 122146 463294
rect 122382 463058 122414 463294
rect 121794 451308 122414 463058
rect 122954 464274 123574 476000
rect 123710 474877 123770 477670
rect 124814 475557 124874 477670
rect 125366 477670 125540 477730
rect 125888 477730 125948 478040
rect 127112 477730 127172 478040
rect 128064 477730 128124 478040
rect 128472 477730 128532 478040
rect 129560 477730 129620 478040
rect 130512 477730 130572 478040
rect 130648 477730 130708 478040
rect 132008 477730 132068 478040
rect 132960 477730 133020 478040
rect 133096 477730 133156 478040
rect 125888 477670 126346 477730
rect 127112 477670 127266 477730
rect 128064 477670 128186 477730
rect 128472 477670 128554 477730
rect 129560 477670 129658 477730
rect 130512 477670 130578 477730
rect 130648 477670 130762 477730
rect 124811 475556 124877 475557
rect 124811 475492 124812 475556
rect 124876 475492 124877 475556
rect 124811 475491 124877 475492
rect 125366 474877 125426 477670
rect 123707 474876 123773 474877
rect 123707 474812 123708 474876
rect 123772 474812 123773 474876
rect 123707 474811 123773 474812
rect 125363 474876 125429 474877
rect 125363 474812 125364 474876
rect 125428 474812 125429 474876
rect 125363 474811 125429 474812
rect 122954 464038 122986 464274
rect 123222 464038 123306 464274
rect 123542 464038 123574 464274
rect 122954 451308 123574 464038
rect 125514 466954 126134 476000
rect 126286 475285 126346 477670
rect 126283 475284 126349 475285
rect 126283 475220 126284 475284
rect 126348 475220 126349 475284
rect 126283 475219 126349 475220
rect 127206 475149 127266 477670
rect 127203 475148 127269 475149
rect 127203 475084 127204 475148
rect 127268 475084 127269 475148
rect 127203 475083 127269 475084
rect 128126 474877 128186 477670
rect 128494 475421 128554 477670
rect 129598 476237 129658 477670
rect 129595 476236 129661 476237
rect 129595 476172 129596 476236
rect 129660 476172 129661 476236
rect 129595 476171 129661 476172
rect 128491 475420 128557 475421
rect 128491 475356 128492 475420
rect 128556 475356 128557 475420
rect 128491 475355 128557 475356
rect 128123 474876 128189 474877
rect 128123 474812 128124 474876
rect 128188 474812 128189 474876
rect 128123 474811 128189 474812
rect 125514 466718 125546 466954
rect 125782 466718 125866 466954
rect 126102 466718 126134 466954
rect 125514 451308 126134 466718
rect 129234 470614 129854 476000
rect 130518 474877 130578 477670
rect 130702 475285 130762 477670
rect 131990 477670 132068 477730
rect 132726 477670 133020 477730
rect 133094 477670 133156 477730
rect 134184 477730 134244 478040
rect 135272 477730 135332 478040
rect 135816 477730 135876 478040
rect 136496 477730 136556 478040
rect 137856 477730 137916 478040
rect 138264 477730 138324 478040
rect 134184 477670 134258 477730
rect 135272 477670 135362 477730
rect 135816 477670 136282 477730
rect 136496 477670 136650 477730
rect 137856 477670 137938 477730
rect 131990 476237 132050 477670
rect 131987 476236 132053 476237
rect 131987 476172 131988 476236
rect 132052 476172 132053 476236
rect 131987 476171 132053 476172
rect 130699 475284 130765 475285
rect 130699 475220 130700 475284
rect 130764 475220 130765 475284
rect 130699 475219 130765 475220
rect 130515 474876 130581 474877
rect 130515 474812 130516 474876
rect 130580 474812 130581 474876
rect 130515 474811 130581 474812
rect 129234 470378 129266 470614
rect 129502 470378 129586 470614
rect 129822 470378 129854 470614
rect 129234 451308 129854 470378
rect 131794 473294 132414 476000
rect 132726 475149 132786 477670
rect 133094 476237 133154 477670
rect 133091 476236 133157 476237
rect 133091 476172 133092 476236
rect 133156 476172 133157 476236
rect 133091 476171 133157 476172
rect 132723 475148 132789 475149
rect 132723 475084 132724 475148
rect 132788 475084 132789 475148
rect 132723 475083 132789 475084
rect 131794 473058 131826 473294
rect 132062 473058 132146 473294
rect 132382 473058 132414 473294
rect 131794 453294 132414 473058
rect 131794 453058 131826 453294
rect 132062 453058 132146 453294
rect 132382 453058 132414 453294
rect 131794 451308 132414 453058
rect 132954 474274 133574 476000
rect 134198 474877 134258 477670
rect 135302 475013 135362 477670
rect 135299 475012 135365 475013
rect 135299 474948 135300 475012
rect 135364 474948 135365 475012
rect 135299 474947 135365 474948
rect 134195 474876 134261 474877
rect 134195 474812 134196 474876
rect 134260 474812 134261 474876
rect 134195 474811 134261 474812
rect 132954 474038 132986 474274
rect 133222 474038 133306 474274
rect 133542 474038 133574 474274
rect 132954 454274 133574 474038
rect 132954 454038 132986 454274
rect 133222 454038 133306 454274
rect 133542 454038 133574 454274
rect 132954 451308 133574 454038
rect 135514 456954 136134 476000
rect 136222 474877 136282 477670
rect 136590 474877 136650 477670
rect 137878 474877 137938 477670
rect 138246 477670 138324 477730
rect 138944 477730 139004 478040
rect 140032 477730 140092 478040
rect 141120 477730 141180 478040
rect 142344 477730 142404 478040
rect 143432 477730 143492 478040
rect 138944 477670 139042 477730
rect 140032 477670 140146 477730
rect 141120 477670 141250 477730
rect 142344 477670 142722 477730
rect 138246 475285 138306 477670
rect 138243 475284 138309 475285
rect 138243 475220 138244 475284
rect 138308 475220 138309 475284
rect 138243 475219 138309 475220
rect 138982 474877 139042 477670
rect 136219 474876 136285 474877
rect 136219 474812 136220 474876
rect 136284 474812 136285 474876
rect 136219 474811 136285 474812
rect 136587 474876 136653 474877
rect 136587 474812 136588 474876
rect 136652 474812 136653 474876
rect 136587 474811 136653 474812
rect 137875 474876 137941 474877
rect 137875 474812 137876 474876
rect 137940 474812 137941 474876
rect 137875 474811 137941 474812
rect 138979 474876 139045 474877
rect 138979 474812 138980 474876
rect 139044 474812 139045 474876
rect 138979 474811 139045 474812
rect 135514 456718 135546 456954
rect 135782 456718 135866 456954
rect 136102 456718 136134 456954
rect 135514 451308 136134 456718
rect 139234 460614 139854 476000
rect 140086 474877 140146 477670
rect 141190 475829 141250 477670
rect 141187 475828 141253 475829
rect 141187 475764 141188 475828
rect 141252 475764 141253 475828
rect 141187 475763 141253 475764
rect 140083 474876 140149 474877
rect 140083 474812 140084 474876
rect 140148 474812 140149 474876
rect 140083 474811 140149 474812
rect 139234 460378 139266 460614
rect 139502 460378 139586 460614
rect 139822 460378 139854 460614
rect 139234 451308 139854 460378
rect 141794 463294 142414 476000
rect 142662 474877 142722 477670
rect 143398 477670 143492 477730
rect 144792 477730 144852 478040
rect 146016 477730 146076 478040
rect 146968 477730 147028 478040
rect 148328 477730 148388 478040
rect 149416 477730 149476 478040
rect 150504 477730 150564 478040
rect 144792 477670 147138 477730
rect 148328 477670 148426 477730
rect 149416 477670 150082 477730
rect 150504 477670 150634 477730
rect 143398 476237 143458 477670
rect 143395 476236 143461 476237
rect 143395 476172 143396 476236
rect 143460 476172 143461 476236
rect 143395 476171 143461 476172
rect 147078 476101 147138 477670
rect 148366 476101 148426 477670
rect 147075 476100 147141 476101
rect 147075 476036 147076 476100
rect 147140 476036 147141 476100
rect 147075 476035 147141 476036
rect 148363 476100 148429 476101
rect 148363 476036 148364 476100
rect 148428 476036 148429 476100
rect 148363 476035 148429 476036
rect 142659 474876 142725 474877
rect 142659 474812 142660 474876
rect 142724 474812 142725 474876
rect 142659 474811 142725 474812
rect 141794 463058 141826 463294
rect 142062 463058 142146 463294
rect 142382 463058 142414 463294
rect 141794 451308 142414 463058
rect 142954 464274 143574 476000
rect 142954 464038 142986 464274
rect 143222 464038 143306 464274
rect 143542 464038 143574 464274
rect 142954 451308 143574 464038
rect 145514 466954 146134 476000
rect 145514 466718 145546 466954
rect 145782 466718 145866 466954
rect 146102 466718 146134 466954
rect 145514 451308 146134 466718
rect 149234 470614 149854 476000
rect 150022 474877 150082 477670
rect 150574 475557 150634 477670
rect 150571 475556 150637 475557
rect 150571 475492 150572 475556
rect 150636 475492 150637 475556
rect 150571 475491 150637 475492
rect 150019 474876 150085 474877
rect 150019 474812 150020 474876
rect 150084 474812 150085 474876
rect 150019 474811 150085 474812
rect 149234 470378 149266 470614
rect 149502 470378 149586 470614
rect 149822 470378 149854 470614
rect 149234 451308 149854 470378
rect 151794 473294 152414 476000
rect 151794 473058 151826 473294
rect 152062 473058 152146 473294
rect 152382 473058 152414 473294
rect 151794 453294 152414 473058
rect 151794 453058 151826 453294
rect 152062 453058 152146 453294
rect 152382 453058 152414 453294
rect 151794 451308 152414 453058
rect 152954 474274 153574 476000
rect 152954 474038 152986 474274
rect 153222 474038 153306 474274
rect 153542 474038 153574 474274
rect 152954 454274 153574 474038
rect 152954 454038 152986 454274
rect 153222 454038 153306 454274
rect 153542 454038 153574 454274
rect 152954 451308 153574 454038
rect 155514 456954 156134 476000
rect 155514 456718 155546 456954
rect 155782 456718 155866 456954
rect 156102 456718 156134 456954
rect 155514 451308 156134 456718
rect 159234 460614 159854 476000
rect 159234 460378 159266 460614
rect 159502 460378 159586 460614
rect 159822 460378 159854 460614
rect 159234 451308 159854 460378
rect 161794 463294 162414 476000
rect 161794 463058 161826 463294
rect 162062 463058 162146 463294
rect 162382 463058 162414 463294
rect 161794 451308 162414 463058
rect 162954 464274 163574 476000
rect 162954 464038 162986 464274
rect 163222 464038 163306 464274
rect 163542 464038 163574 464274
rect 162954 451308 163574 464038
rect 165514 466954 166134 476000
rect 165514 466718 165546 466954
rect 165782 466718 165866 466954
rect 166102 466718 166134 466954
rect 165514 451308 166134 466718
rect 48083 451283 48149 451284
rect 48086 449850 48146 451283
rect 35206 449790 35780 449850
rect 46798 449790 46932 449850
rect 48086 449790 48156 449850
rect 35720 449202 35780 449790
rect 46872 449202 46932 449790
rect 48096 449202 48156 449790
rect 25514 446718 25546 446954
rect 25782 446718 25866 446954
rect 26102 446718 26134 446954
rect 25514 426954 26134 446718
rect 30952 443294 31300 443456
rect 30952 443058 31008 443294
rect 31244 443058 31300 443294
rect 30952 442896 31300 443058
rect 165320 443294 165668 443456
rect 165320 443058 165376 443294
rect 165612 443058 165668 443294
rect 165320 442896 165668 443058
rect 30272 433294 30620 433456
rect 30272 433058 30328 433294
rect 30564 433058 30620 433294
rect 30272 432896 30620 433058
rect 166000 433294 166348 433456
rect 166000 433058 166056 433294
rect 166292 433058 166348 433294
rect 166000 432896 166348 433058
rect 25514 426718 25546 426954
rect 25782 426718 25866 426954
rect 26102 426718 26134 426954
rect 25514 406954 26134 426718
rect 166950 425645 167010 587691
rect 168419 584900 168485 584901
rect 168419 584836 168420 584900
rect 168484 584836 168485 584900
rect 168419 584835 168485 584836
rect 167131 584764 167197 584765
rect 167131 584700 167132 584764
rect 167196 584700 167197 584764
rect 167131 584699 167197 584700
rect 167134 476237 167194 584699
rect 167683 581636 167749 581637
rect 167683 581572 167684 581636
rect 167748 581572 167749 581636
rect 167683 581571 167749 581572
rect 167131 476236 167197 476237
rect 167131 476172 167132 476236
rect 167196 476172 167197 476236
rect 167131 476171 167197 476172
rect 167499 451892 167565 451893
rect 167499 451828 167500 451892
rect 167564 451828 167565 451892
rect 167499 451827 167565 451828
rect 167131 449988 167197 449989
rect 167131 449924 167132 449988
rect 167196 449924 167197 449988
rect 167131 449923 167197 449924
rect 166947 425644 167013 425645
rect 166947 425580 166948 425644
rect 167012 425580 167013 425644
rect 166947 425579 167013 425580
rect 30952 423294 31300 423456
rect 30952 423058 31008 423294
rect 31244 423058 31300 423294
rect 30952 422896 31300 423058
rect 165320 423294 165668 423456
rect 165320 423058 165376 423294
rect 165612 423058 165668 423294
rect 165320 422896 165668 423058
rect 30272 413294 30620 413456
rect 30272 413058 30328 413294
rect 30564 413058 30620 413294
rect 30272 412896 30620 413058
rect 166000 413294 166348 413456
rect 166000 413058 166056 413294
rect 166292 413058 166348 413294
rect 166000 412896 166348 413058
rect 25514 406718 25546 406954
rect 25782 406718 25866 406954
rect 26102 406718 26134 406954
rect 25514 386954 26134 406718
rect 30952 403294 31300 403456
rect 30952 403058 31008 403294
rect 31244 403058 31300 403294
rect 30952 402896 31300 403058
rect 165320 403294 165668 403456
rect 165320 403058 165376 403294
rect 165612 403058 165668 403294
rect 165320 402896 165668 403058
rect 30272 393294 30620 393456
rect 30272 393058 30328 393294
rect 30564 393058 30620 393294
rect 30272 392896 30620 393058
rect 166000 393294 166348 393456
rect 166000 393058 166056 393294
rect 166292 393058 166348 393294
rect 166000 392896 166348 393058
rect 25514 386718 25546 386954
rect 25782 386718 25866 386954
rect 26102 386718 26134 386954
rect 25514 366954 26134 386718
rect 30952 383294 31300 383456
rect 30952 383058 31008 383294
rect 31244 383058 31300 383294
rect 30952 382896 31300 383058
rect 165320 383294 165668 383456
rect 165320 383058 165376 383294
rect 165612 383058 165668 383294
rect 165320 382896 165668 383058
rect 30272 373294 30620 373456
rect 30272 373058 30328 373294
rect 30564 373058 30620 373294
rect 30272 372896 30620 373058
rect 166000 373294 166348 373456
rect 166000 373058 166056 373294
rect 166292 373058 166348 373294
rect 166000 372896 166348 373058
rect 25514 366718 25546 366954
rect 25782 366718 25866 366954
rect 26102 366718 26134 366954
rect 25514 346954 26134 366718
rect 43200 365530 43260 366106
rect 43118 365470 43260 365530
rect 43336 365530 43396 366106
rect 60608 365530 60668 366106
rect 63192 365530 63252 366106
rect 43336 365470 43546 365530
rect 43118 364309 43178 365470
rect 43115 364308 43181 364309
rect 43115 364244 43116 364308
rect 43180 364244 43181 364308
rect 43115 364243 43181 364244
rect 43486 364173 43546 365470
rect 60598 365470 60668 365530
rect 63174 365470 63252 365530
rect 65640 365530 65700 366106
rect 68088 365530 68148 366106
rect 70672 365530 70732 366106
rect 73120 365530 73180 366106
rect 65640 365470 65810 365530
rect 68088 365470 68202 365530
rect 70672 365470 70778 365530
rect 43483 364172 43549 364173
rect 43483 364108 43484 364172
rect 43548 364108 43549 364172
rect 43483 364107 43549 364108
rect 25514 346718 25546 346954
rect 25782 346718 25866 346954
rect 26102 346718 26134 346954
rect 25514 326954 26134 346718
rect 29234 350614 29854 364000
rect 29234 350378 29266 350614
rect 29502 350378 29586 350614
rect 29822 350378 29854 350614
rect 29234 339308 29854 350378
rect 31794 353294 32414 364000
rect 31794 353058 31826 353294
rect 32062 353058 32146 353294
rect 32382 353058 32414 353294
rect 31794 339308 32414 353058
rect 32954 354274 33574 364000
rect 32954 354038 32986 354274
rect 33222 354038 33306 354274
rect 33542 354038 33574 354274
rect 32954 339308 33574 354038
rect 35514 356954 36134 364000
rect 35514 356718 35546 356954
rect 35782 356718 35866 356954
rect 36102 356718 36134 356954
rect 35203 339556 35269 339557
rect 35203 339492 35204 339556
rect 35268 339492 35269 339556
rect 35203 339491 35269 339492
rect 35206 337650 35266 339491
rect 35514 339308 36134 356718
rect 39234 360614 39854 364000
rect 39234 360378 39266 360614
rect 39502 360378 39586 360614
rect 39822 360378 39854 360614
rect 39234 340614 39854 360378
rect 39234 340378 39266 340614
rect 39502 340378 39586 340614
rect 39822 340378 39854 340614
rect 39234 339308 39854 340378
rect 41794 363294 42414 364000
rect 41794 363058 41826 363294
rect 42062 363058 42146 363294
rect 42382 363058 42414 363294
rect 41794 343294 42414 363058
rect 41794 343058 41826 343294
rect 42062 343058 42146 343294
rect 42382 343058 42414 343294
rect 41794 339308 42414 343058
rect 42954 344274 43574 364000
rect 42954 344038 42986 344274
rect 43222 344038 43306 344274
rect 43542 344038 43574 344274
rect 42954 339308 43574 344038
rect 45514 346954 46134 364000
rect 45514 346718 45546 346954
rect 45782 346718 45866 346954
rect 46102 346718 46134 346954
rect 45514 339308 46134 346718
rect 49234 350614 49854 364000
rect 49234 350378 49266 350614
rect 49502 350378 49586 350614
rect 49822 350378 49854 350614
rect 48083 340780 48149 340781
rect 48083 340716 48084 340780
rect 48148 340716 48149 340780
rect 48083 340715 48149 340716
rect 46795 340236 46861 340237
rect 46795 340172 46796 340236
rect 46860 340172 46861 340236
rect 46795 340171 46861 340172
rect 46798 337650 46858 340171
rect 48086 337650 48146 340715
rect 49234 339308 49854 350378
rect 51794 353294 52414 364000
rect 51794 353058 51826 353294
rect 52062 353058 52146 353294
rect 52382 353058 52414 353294
rect 51794 339308 52414 353058
rect 52954 354274 53574 364000
rect 52954 354038 52986 354274
rect 53222 354038 53306 354274
rect 53542 354038 53574 354274
rect 52954 339308 53574 354038
rect 55514 356954 56134 364000
rect 55514 356718 55546 356954
rect 55782 356718 55866 356954
rect 56102 356718 56134 356954
rect 55514 339308 56134 356718
rect 59234 360614 59854 364000
rect 60598 363085 60658 365470
rect 63174 364173 63234 365470
rect 65750 364173 65810 365470
rect 63171 364172 63237 364173
rect 63171 364108 63172 364172
rect 63236 364108 63237 364172
rect 63171 364107 63237 364108
rect 65747 364172 65813 364173
rect 65747 364108 65748 364172
rect 65812 364108 65813 364172
rect 65747 364107 65813 364108
rect 61794 363294 62414 364000
rect 60595 363084 60661 363085
rect 60595 363020 60596 363084
rect 60660 363020 60661 363084
rect 60595 363019 60661 363020
rect 61794 363058 61826 363294
rect 62062 363058 62146 363294
rect 62382 363058 62414 363294
rect 59234 360378 59266 360614
rect 59502 360378 59586 360614
rect 59822 360378 59854 360614
rect 59234 340614 59854 360378
rect 59234 340378 59266 340614
rect 59502 340378 59586 340614
rect 59822 340378 59854 340614
rect 59234 339308 59854 340378
rect 61794 343294 62414 363058
rect 61794 343058 61826 343294
rect 62062 343058 62146 343294
rect 62382 343058 62414 343294
rect 61794 339308 62414 343058
rect 62954 344274 63574 364000
rect 62954 344038 62986 344274
rect 63222 344038 63306 344274
rect 63542 344038 63574 344274
rect 62954 339308 63574 344038
rect 65514 346954 66134 364000
rect 68142 363085 68202 365470
rect 68139 363084 68205 363085
rect 68139 363020 68140 363084
rect 68204 363020 68205 363084
rect 68139 363019 68205 363020
rect 65514 346718 65546 346954
rect 65782 346718 65866 346954
rect 66102 346718 66134 346954
rect 65514 339308 66134 346718
rect 69234 350614 69854 364000
rect 70718 363085 70778 365470
rect 73110 365470 73180 365530
rect 75568 365530 75628 366106
rect 78016 365530 78076 366106
rect 80600 365530 80660 366106
rect 83048 365530 83108 366106
rect 85632 365530 85692 366106
rect 75568 365470 75746 365530
rect 78016 365470 78138 365530
rect 80600 365470 80714 365530
rect 73110 364173 73170 365470
rect 75686 364173 75746 365470
rect 73107 364172 73173 364173
rect 73107 364108 73108 364172
rect 73172 364108 73173 364172
rect 73107 364107 73173 364108
rect 75683 364172 75749 364173
rect 75683 364108 75684 364172
rect 75748 364108 75749 364172
rect 75683 364107 75749 364108
rect 70715 363084 70781 363085
rect 70715 363020 70716 363084
rect 70780 363020 70781 363084
rect 70715 363019 70781 363020
rect 69234 350378 69266 350614
rect 69502 350378 69586 350614
rect 69822 350378 69854 350614
rect 69234 339308 69854 350378
rect 71794 353294 72414 364000
rect 71794 353058 71826 353294
rect 72062 353058 72146 353294
rect 72382 353058 72414 353294
rect 71794 339308 72414 353058
rect 72954 354274 73574 364000
rect 72954 354038 72986 354274
rect 73222 354038 73306 354274
rect 73542 354038 73574 354274
rect 72954 339308 73574 354038
rect 75514 356954 76134 364000
rect 78078 363085 78138 365470
rect 78075 363084 78141 363085
rect 78075 363020 78076 363084
rect 78140 363020 78141 363084
rect 78075 363019 78141 363020
rect 75514 356718 75546 356954
rect 75782 356718 75866 356954
rect 76102 356718 76134 356954
rect 75514 339308 76134 356718
rect 79234 360614 79854 364000
rect 80654 363085 80714 365470
rect 83046 365470 83108 365530
rect 85622 365470 85692 365530
rect 88080 365530 88140 366106
rect 90664 365530 90724 366106
rect 93112 365530 93172 366106
rect 95560 365530 95620 366106
rect 88080 365470 88258 365530
rect 90664 365470 90834 365530
rect 93112 365470 93226 365530
rect 83046 364173 83106 365470
rect 85622 364173 85682 365470
rect 83043 364172 83109 364173
rect 83043 364108 83044 364172
rect 83108 364108 83109 364172
rect 83043 364107 83109 364108
rect 85619 364172 85685 364173
rect 85619 364108 85620 364172
rect 85684 364108 85685 364172
rect 85619 364107 85685 364108
rect 81794 363294 82414 364000
rect 80651 363084 80717 363085
rect 80651 363020 80652 363084
rect 80716 363020 80717 363084
rect 80651 363019 80717 363020
rect 81794 363058 81826 363294
rect 82062 363058 82146 363294
rect 82382 363058 82414 363294
rect 79234 360378 79266 360614
rect 79502 360378 79586 360614
rect 79822 360378 79854 360614
rect 79234 340614 79854 360378
rect 79234 340378 79266 340614
rect 79502 340378 79586 340614
rect 79822 340378 79854 340614
rect 79234 339308 79854 340378
rect 81794 343294 82414 363058
rect 81794 343058 81826 343294
rect 82062 343058 82146 343294
rect 82382 343058 82414 343294
rect 81794 339308 82414 343058
rect 82954 344274 83574 364000
rect 82954 344038 82986 344274
rect 83222 344038 83306 344274
rect 83542 344038 83574 344274
rect 82954 339308 83574 344038
rect 85514 346954 86134 364000
rect 88198 363085 88258 365470
rect 88195 363084 88261 363085
rect 88195 363020 88196 363084
rect 88260 363020 88261 363084
rect 88195 363019 88261 363020
rect 85514 346718 85546 346954
rect 85782 346718 85866 346954
rect 86102 346718 86134 346954
rect 85514 339308 86134 346718
rect 89234 350614 89854 364000
rect 90774 363085 90834 365470
rect 93166 364173 93226 365470
rect 95558 365470 95620 365530
rect 98280 365530 98340 366106
rect 100592 365530 100652 366106
rect 98280 365470 98378 365530
rect 95558 364173 95618 365470
rect 93163 364172 93229 364173
rect 93163 364108 93164 364172
rect 93228 364108 93229 364172
rect 93163 364107 93229 364108
rect 95555 364172 95621 364173
rect 95555 364108 95556 364172
rect 95620 364108 95621 364172
rect 95555 364107 95621 364108
rect 90771 363084 90837 363085
rect 90771 363020 90772 363084
rect 90836 363020 90837 363084
rect 90771 363019 90837 363020
rect 89234 350378 89266 350614
rect 89502 350378 89586 350614
rect 89822 350378 89854 350614
rect 89234 339308 89854 350378
rect 91794 353294 92414 364000
rect 91794 353058 91826 353294
rect 92062 353058 92146 353294
rect 92382 353058 92414 353294
rect 91794 339308 92414 353058
rect 92954 354274 93574 364000
rect 92954 354038 92986 354274
rect 93222 354038 93306 354274
rect 93542 354038 93574 354274
rect 92954 339308 93574 354038
rect 95514 356954 96134 364000
rect 98318 363085 98378 365470
rect 100526 365470 100652 365530
rect 103040 365530 103100 366106
rect 105624 365530 105684 366106
rect 107392 365530 107452 366106
rect 108072 365530 108132 366106
rect 108480 365530 108540 366106
rect 109568 365530 109628 366106
rect 110520 365530 110580 366106
rect 103040 365470 103162 365530
rect 105624 365470 105738 365530
rect 98315 363084 98381 363085
rect 98315 363020 98316 363084
rect 98380 363020 98381 363084
rect 98315 363019 98381 363020
rect 95514 356718 95546 356954
rect 95782 356718 95866 356954
rect 96102 356718 96134 356954
rect 95514 339308 96134 356718
rect 99234 360614 99854 364000
rect 100526 363085 100586 365470
rect 103102 364173 103162 365470
rect 105678 364173 105738 365470
rect 107334 365470 107452 365530
rect 108070 365470 108132 365530
rect 108438 365470 108540 365530
rect 109542 365470 109628 365530
rect 110462 365470 110580 365530
rect 110792 365530 110852 366106
rect 112152 365530 112212 366106
rect 110792 365470 110890 365530
rect 103099 364172 103165 364173
rect 103099 364108 103100 364172
rect 103164 364108 103165 364172
rect 103099 364107 103165 364108
rect 105675 364172 105741 364173
rect 105675 364108 105676 364172
rect 105740 364108 105741 364172
rect 105675 364107 105741 364108
rect 101794 363294 102414 364000
rect 100523 363084 100589 363085
rect 100523 363020 100524 363084
rect 100588 363020 100589 363084
rect 100523 363019 100589 363020
rect 101794 363058 101826 363294
rect 102062 363058 102146 363294
rect 102382 363058 102414 363294
rect 99234 360378 99266 360614
rect 99502 360378 99586 360614
rect 99822 360378 99854 360614
rect 99234 340614 99854 360378
rect 99234 340378 99266 340614
rect 99502 340378 99586 340614
rect 99822 340378 99854 340614
rect 99234 339308 99854 340378
rect 101794 343294 102414 363058
rect 101794 343058 101826 343294
rect 102062 343058 102146 343294
rect 102382 343058 102414 343294
rect 101794 339308 102414 343058
rect 102954 344274 103574 364000
rect 102954 344038 102986 344274
rect 103222 344038 103306 344274
rect 103542 344038 103574 344274
rect 102954 339308 103574 344038
rect 105514 346954 106134 364000
rect 107334 363085 107394 365470
rect 108070 363357 108130 365470
rect 108067 363356 108133 363357
rect 108067 363292 108068 363356
rect 108132 363292 108133 363356
rect 108067 363291 108133 363292
rect 108438 363085 108498 365470
rect 109542 364173 109602 365470
rect 109539 364172 109605 364173
rect 109539 364108 109540 364172
rect 109604 364108 109605 364172
rect 109539 364107 109605 364108
rect 107331 363084 107397 363085
rect 107331 363020 107332 363084
rect 107396 363020 107397 363084
rect 107331 363019 107397 363020
rect 108435 363084 108501 363085
rect 108435 363020 108436 363084
rect 108500 363020 108501 363084
rect 108435 363019 108501 363020
rect 105514 346718 105546 346954
rect 105782 346718 105866 346954
rect 106102 346718 106134 346954
rect 105514 339308 106134 346718
rect 109234 350614 109854 364000
rect 110462 363221 110522 365470
rect 110459 363220 110525 363221
rect 110459 363156 110460 363220
rect 110524 363156 110525 363220
rect 110459 363155 110525 363156
rect 110830 363085 110890 365470
rect 112118 365470 112212 365530
rect 112968 365530 113028 366106
rect 113240 365530 113300 366106
rect 114328 365530 114388 366106
rect 112968 365470 113098 365530
rect 112118 364309 112178 365470
rect 112115 364308 112181 364309
rect 112115 364244 112116 364308
rect 112180 364244 112181 364308
rect 112115 364243 112181 364244
rect 113038 364173 113098 365470
rect 113222 365470 113300 365530
rect 114326 365470 114388 365530
rect 115416 365530 115476 366106
rect 115552 365530 115612 366106
rect 116776 365530 116836 366106
rect 117864 365530 117924 366106
rect 115416 365470 115490 365530
rect 115552 365470 115674 365530
rect 113222 364173 113282 365470
rect 113035 364172 113101 364173
rect 113035 364108 113036 364172
rect 113100 364108 113101 364172
rect 113035 364107 113101 364108
rect 113219 364172 113285 364173
rect 113219 364108 113220 364172
rect 113284 364108 113285 364172
rect 113219 364107 113285 364108
rect 110827 363084 110893 363085
rect 110827 363020 110828 363084
rect 110892 363020 110893 363084
rect 110827 363019 110893 363020
rect 109234 350378 109266 350614
rect 109502 350378 109586 350614
rect 109822 350378 109854 350614
rect 109234 339308 109854 350378
rect 111794 353294 112414 364000
rect 111794 353058 111826 353294
rect 112062 353058 112146 353294
rect 112382 353058 112414 353294
rect 111794 339308 112414 353058
rect 112954 354274 113574 364000
rect 114326 363085 114386 365470
rect 115430 364309 115490 365470
rect 115427 364308 115493 364309
rect 115427 364244 115428 364308
rect 115492 364244 115493 364308
rect 115427 364243 115493 364244
rect 115614 364173 115674 365470
rect 116718 365470 116836 365530
rect 117822 365470 117924 365530
rect 118272 365530 118332 366106
rect 118952 365530 119012 366106
rect 118272 365470 118434 365530
rect 115611 364172 115677 364173
rect 115611 364108 115612 364172
rect 115676 364108 115677 364172
rect 115611 364107 115677 364108
rect 114323 363084 114389 363085
rect 114323 363020 114324 363084
rect 114388 363020 114389 363084
rect 114323 363019 114389 363020
rect 112954 354038 112986 354274
rect 113222 354038 113306 354274
rect 113542 354038 113574 354274
rect 112954 339308 113574 354038
rect 115514 356954 116134 364000
rect 116718 363085 116778 365470
rect 117822 363221 117882 365470
rect 117819 363220 117885 363221
rect 117819 363156 117820 363220
rect 117884 363156 117885 363220
rect 117819 363155 117885 363156
rect 118374 363085 118434 365470
rect 118926 365470 119012 365530
rect 120176 365530 120236 366106
rect 120584 365530 120644 366106
rect 120176 365470 120274 365530
rect 118926 363357 118986 365470
rect 120214 364037 120274 365470
rect 120582 365470 120644 365530
rect 121264 365530 121324 366106
rect 122624 365530 122684 366106
rect 123032 365530 123092 366106
rect 123712 365530 123772 366106
rect 121264 365470 121378 365530
rect 120211 364036 120277 364037
rect 118923 363356 118989 363357
rect 118923 363292 118924 363356
rect 118988 363292 118989 363356
rect 118923 363291 118989 363292
rect 116715 363084 116781 363085
rect 116715 363020 116716 363084
rect 116780 363020 116781 363084
rect 116715 363019 116781 363020
rect 118371 363084 118437 363085
rect 118371 363020 118372 363084
rect 118436 363020 118437 363084
rect 118371 363019 118437 363020
rect 115514 356718 115546 356954
rect 115782 356718 115866 356954
rect 116102 356718 116134 356954
rect 115514 339308 116134 356718
rect 119234 360614 119854 364000
rect 120211 363972 120212 364036
rect 120276 363972 120277 364036
rect 120211 363971 120277 363972
rect 120582 363221 120642 365470
rect 120579 363220 120645 363221
rect 120579 363156 120580 363220
rect 120644 363156 120645 363220
rect 120579 363155 120645 363156
rect 121318 363085 121378 365470
rect 122606 365470 122684 365530
rect 122974 365470 123092 365530
rect 123710 365470 123772 365530
rect 124800 365530 124860 366106
rect 125480 365530 125540 366106
rect 124800 365470 124874 365530
rect 121794 363294 122414 364000
rect 122606 363901 122666 365470
rect 122974 364173 123034 365470
rect 122971 364172 123037 364173
rect 122971 364108 122972 364172
rect 123036 364108 123037 364172
rect 122971 364107 123037 364108
rect 122603 363900 122669 363901
rect 122603 363836 122604 363900
rect 122668 363836 122669 363900
rect 122603 363835 122669 363836
rect 121315 363084 121381 363085
rect 121315 363020 121316 363084
rect 121380 363020 121381 363084
rect 121315 363019 121381 363020
rect 121794 363058 121826 363294
rect 122062 363058 122146 363294
rect 122382 363058 122414 363294
rect 119234 360378 119266 360614
rect 119502 360378 119586 360614
rect 119822 360378 119854 360614
rect 119234 340614 119854 360378
rect 119234 340378 119266 340614
rect 119502 340378 119586 340614
rect 119822 340378 119854 340614
rect 119234 339308 119854 340378
rect 121794 343294 122414 363058
rect 121794 343058 121826 343294
rect 122062 343058 122146 343294
rect 122382 343058 122414 343294
rect 121794 339308 122414 343058
rect 122954 344274 123574 364000
rect 123710 363493 123770 365470
rect 123707 363492 123773 363493
rect 123707 363428 123708 363492
rect 123772 363428 123773 363492
rect 123707 363427 123773 363428
rect 124814 363221 124874 365470
rect 125366 365470 125540 365530
rect 125888 365530 125948 366106
rect 127112 365530 127172 366106
rect 128064 365530 128124 366106
rect 128472 365530 128532 366106
rect 129560 365530 129620 366106
rect 130512 365530 130572 366106
rect 130648 365530 130708 366106
rect 132008 365530 132068 366106
rect 132960 365530 133020 366106
rect 133096 365530 133156 366106
rect 125888 365470 125978 365530
rect 127112 365470 127266 365530
rect 128064 365470 128186 365530
rect 128472 365470 128554 365530
rect 129560 365470 129658 365530
rect 130512 365470 130578 365530
rect 130648 365470 130762 365530
rect 124811 363220 124877 363221
rect 124811 363156 124812 363220
rect 124876 363156 124877 363220
rect 124811 363155 124877 363156
rect 125366 363085 125426 365470
rect 125918 364173 125978 365470
rect 125915 364172 125981 364173
rect 125915 364108 125916 364172
rect 125980 364108 125981 364172
rect 125915 364107 125981 364108
rect 125363 363084 125429 363085
rect 125363 363020 125364 363084
rect 125428 363020 125429 363084
rect 125363 363019 125429 363020
rect 122954 344038 122986 344274
rect 123222 344038 123306 344274
rect 123542 344038 123574 344274
rect 122954 339308 123574 344038
rect 125514 346954 126134 364000
rect 127206 363765 127266 365470
rect 127203 363764 127269 363765
rect 127203 363700 127204 363764
rect 127268 363700 127269 363764
rect 127203 363699 127269 363700
rect 128126 363085 128186 365470
rect 128494 363085 128554 365470
rect 129598 364173 129658 365470
rect 129595 364172 129661 364173
rect 129595 364108 129596 364172
rect 129660 364108 129661 364172
rect 129595 364107 129661 364108
rect 128123 363084 128189 363085
rect 128123 363020 128124 363084
rect 128188 363020 128189 363084
rect 128123 363019 128189 363020
rect 128491 363084 128557 363085
rect 128491 363020 128492 363084
rect 128556 363020 128557 363084
rect 128491 363019 128557 363020
rect 125514 346718 125546 346954
rect 125782 346718 125866 346954
rect 126102 346718 126134 346954
rect 125514 339308 126134 346718
rect 129234 350614 129854 364000
rect 130518 363085 130578 365470
rect 130702 363221 130762 365470
rect 131990 365470 132068 365530
rect 132910 365470 133020 365530
rect 133094 365470 133156 365530
rect 134184 365530 134244 366106
rect 135272 365530 135332 366106
rect 135816 365530 135876 366106
rect 136496 365530 136556 366106
rect 137856 365530 137916 366106
rect 138264 365530 138324 366106
rect 134184 365470 134258 365530
rect 135272 365470 135362 365530
rect 135816 365470 135914 365530
rect 136496 365470 136650 365530
rect 137856 365470 137938 365530
rect 131990 364173 132050 365470
rect 132910 364309 132970 365470
rect 132907 364308 132973 364309
rect 132907 364244 132908 364308
rect 132972 364244 132973 364308
rect 132907 364243 132973 364244
rect 133094 364173 133154 365470
rect 131987 364172 132053 364173
rect 131987 364108 131988 364172
rect 132052 364108 132053 364172
rect 131987 364107 132053 364108
rect 133091 364172 133157 364173
rect 133091 364108 133092 364172
rect 133156 364108 133157 364172
rect 133091 364107 133157 364108
rect 130699 363220 130765 363221
rect 130699 363156 130700 363220
rect 130764 363156 130765 363220
rect 130699 363155 130765 363156
rect 130515 363084 130581 363085
rect 130515 363020 130516 363084
rect 130580 363020 130581 363084
rect 130515 363019 130581 363020
rect 129234 350378 129266 350614
rect 129502 350378 129586 350614
rect 129822 350378 129854 350614
rect 129234 339308 129854 350378
rect 131794 353294 132414 364000
rect 131794 353058 131826 353294
rect 132062 353058 132146 353294
rect 132382 353058 132414 353294
rect 131794 339308 132414 353058
rect 132954 354274 133574 364000
rect 134198 363085 134258 365470
rect 135302 364309 135362 365470
rect 135299 364308 135365 364309
rect 135299 364244 135300 364308
rect 135364 364244 135365 364308
rect 135299 364243 135365 364244
rect 135854 364173 135914 365470
rect 135851 364172 135917 364173
rect 135851 364108 135852 364172
rect 135916 364108 135917 364172
rect 135851 364107 135917 364108
rect 134195 363084 134261 363085
rect 134195 363020 134196 363084
rect 134260 363020 134261 363084
rect 134195 363019 134261 363020
rect 132954 354038 132986 354274
rect 133222 354038 133306 354274
rect 133542 354038 133574 354274
rect 132954 339308 133574 354038
rect 135514 356954 136134 364000
rect 136590 363901 136650 365470
rect 136587 363900 136653 363901
rect 136587 363836 136588 363900
rect 136652 363836 136653 363900
rect 136587 363835 136653 363836
rect 137878 363085 137938 365470
rect 138246 365470 138324 365530
rect 138944 365530 139004 366106
rect 140032 365530 140092 366106
rect 141120 365530 141180 366106
rect 142344 365530 142404 366106
rect 143432 365530 143492 366106
rect 144792 365530 144852 366106
rect 146016 365530 146076 366106
rect 146968 365530 147028 366106
rect 148328 365530 148388 366106
rect 149416 365530 149476 366106
rect 150504 365530 150564 366106
rect 138944 365470 139042 365530
rect 140032 365470 140146 365530
rect 141120 365470 141250 365530
rect 138246 363493 138306 365470
rect 138243 363492 138309 363493
rect 138243 363428 138244 363492
rect 138308 363428 138309 363492
rect 138243 363427 138309 363428
rect 138982 363085 139042 365470
rect 137875 363084 137941 363085
rect 137875 363020 137876 363084
rect 137940 363020 137941 363084
rect 137875 363019 137941 363020
rect 138979 363084 139045 363085
rect 138979 363020 138980 363084
rect 139044 363020 139045 363084
rect 138979 363019 139045 363020
rect 135514 356718 135546 356954
rect 135782 356718 135866 356954
rect 136102 356718 136134 356954
rect 135514 339308 136134 356718
rect 139234 360614 139854 364000
rect 140086 363085 140146 365470
rect 141190 363085 141250 365470
rect 142294 365470 142404 365530
rect 143398 365470 143492 365530
rect 144686 365470 144852 365530
rect 145974 365470 148426 365530
rect 149416 365470 149530 365530
rect 150504 365470 150634 365530
rect 142294 364173 142354 365470
rect 143398 364309 143458 365470
rect 144686 364309 144746 365470
rect 145974 364309 146034 365470
rect 143395 364308 143461 364309
rect 143395 364244 143396 364308
rect 143460 364244 143461 364308
rect 143395 364243 143461 364244
rect 144683 364308 144749 364309
rect 144683 364244 144684 364308
rect 144748 364244 144749 364308
rect 144683 364243 144749 364244
rect 145971 364308 146037 364309
rect 145971 364244 145972 364308
rect 146036 364244 146037 364308
rect 145971 364243 146037 364244
rect 142291 364172 142357 364173
rect 142291 364108 142292 364172
rect 142356 364108 142357 364172
rect 142291 364107 142357 364108
rect 141794 363294 142414 364000
rect 140083 363084 140149 363085
rect 140083 363020 140084 363084
rect 140148 363020 140149 363084
rect 140083 363019 140149 363020
rect 141187 363084 141253 363085
rect 141187 363020 141188 363084
rect 141252 363020 141253 363084
rect 141187 363019 141253 363020
rect 141794 363058 141826 363294
rect 142062 363058 142146 363294
rect 142382 363058 142414 363294
rect 139234 360378 139266 360614
rect 139502 360378 139586 360614
rect 139822 360378 139854 360614
rect 139234 340614 139854 360378
rect 139234 340378 139266 340614
rect 139502 340378 139586 340614
rect 139822 340378 139854 340614
rect 139234 339308 139854 340378
rect 141794 343294 142414 363058
rect 141794 343058 141826 343294
rect 142062 343058 142146 343294
rect 142382 343058 142414 343294
rect 141794 339308 142414 343058
rect 142954 344274 143574 364000
rect 142954 344038 142986 344274
rect 143222 344038 143306 344274
rect 143542 344038 143574 344274
rect 142954 339308 143574 344038
rect 145514 346954 146134 364000
rect 148366 363085 148426 365470
rect 149470 364173 149530 365470
rect 149467 364172 149533 364173
rect 149467 364108 149468 364172
rect 149532 364108 149533 364172
rect 149467 364107 149533 364108
rect 148363 363084 148429 363085
rect 148363 363020 148364 363084
rect 148428 363020 148429 363084
rect 148363 363019 148429 363020
rect 145514 346718 145546 346954
rect 145782 346718 145866 346954
rect 146102 346718 146134 346954
rect 145514 339308 146134 346718
rect 149234 350614 149854 364000
rect 150574 363629 150634 365470
rect 150571 363628 150637 363629
rect 150571 363564 150572 363628
rect 150636 363564 150637 363628
rect 150571 363563 150637 363564
rect 149234 350378 149266 350614
rect 149502 350378 149586 350614
rect 149822 350378 149854 350614
rect 149234 339308 149854 350378
rect 151794 353294 152414 364000
rect 151794 353058 151826 353294
rect 152062 353058 152146 353294
rect 152382 353058 152414 353294
rect 151794 339308 152414 353058
rect 152954 354274 153574 364000
rect 152954 354038 152986 354274
rect 153222 354038 153306 354274
rect 153542 354038 153574 354274
rect 152954 339308 153574 354038
rect 155514 356954 156134 364000
rect 155514 356718 155546 356954
rect 155782 356718 155866 356954
rect 156102 356718 156134 356954
rect 155514 339308 156134 356718
rect 159234 360614 159854 364000
rect 159234 360378 159266 360614
rect 159502 360378 159586 360614
rect 159822 360378 159854 360614
rect 159234 340614 159854 360378
rect 159234 340378 159266 340614
rect 159502 340378 159586 340614
rect 159822 340378 159854 340614
rect 159234 339308 159854 340378
rect 161794 363294 162414 364000
rect 161794 363058 161826 363294
rect 162062 363058 162146 363294
rect 162382 363058 162414 363294
rect 161794 343294 162414 363058
rect 161794 343058 161826 343294
rect 162062 343058 162146 343294
rect 162382 343058 162414 343294
rect 161794 339308 162414 343058
rect 162954 344274 163574 364000
rect 162954 344038 162986 344274
rect 163222 344038 163306 344274
rect 163542 344038 163574 344274
rect 162954 339308 163574 344038
rect 165514 346954 166134 364000
rect 166950 363901 167010 425579
rect 167134 364173 167194 449923
rect 167131 364172 167197 364173
rect 167131 364108 167132 364172
rect 167196 364108 167197 364172
rect 167131 364107 167197 364108
rect 166947 363900 167013 363901
rect 166947 363836 166948 363900
rect 167012 363836 167013 363900
rect 166947 363835 167013 363836
rect 167134 363357 167194 364107
rect 167131 363356 167197 363357
rect 167131 363292 167132 363356
rect 167196 363292 167197 363356
rect 167131 363291 167197 363292
rect 165514 346718 165546 346954
rect 165782 346718 165866 346954
rect 166102 346718 166134 346954
rect 165514 339308 166134 346718
rect 35206 337590 35780 337650
rect 46798 337590 46932 337650
rect 48086 337590 48156 337650
rect 35720 337280 35780 337590
rect 46872 337280 46932 337590
rect 48096 337280 48156 337590
rect 30272 333294 30620 333456
rect 30272 333058 30328 333294
rect 30564 333058 30620 333294
rect 30272 332896 30620 333058
rect 166000 333294 166348 333456
rect 166000 333058 166056 333294
rect 166292 333058 166348 333294
rect 166000 332896 166348 333058
rect 25514 326718 25546 326954
rect 25782 326718 25866 326954
rect 26102 326718 26134 326954
rect 25514 306954 26134 326718
rect 30952 323294 31300 323456
rect 30952 323058 31008 323294
rect 31244 323058 31300 323294
rect 30952 322896 31300 323058
rect 165320 323294 165668 323456
rect 165320 323058 165376 323294
rect 165612 323058 165668 323294
rect 165320 322896 165668 323058
rect 30272 313294 30620 313456
rect 30272 313058 30328 313294
rect 30564 313058 30620 313294
rect 30272 312896 30620 313058
rect 166000 313294 166348 313456
rect 166000 313058 166056 313294
rect 166292 313058 166348 313294
rect 166000 312896 166348 313058
rect 25514 306718 25546 306954
rect 25782 306718 25866 306954
rect 26102 306718 26134 306954
rect 25514 286954 26134 306718
rect 30952 303294 31300 303456
rect 30952 303058 31008 303294
rect 31244 303058 31300 303294
rect 30952 302896 31300 303058
rect 165320 303294 165668 303456
rect 165320 303058 165376 303294
rect 165612 303058 165668 303294
rect 165320 302896 165668 303058
rect 30272 293294 30620 293456
rect 30272 293058 30328 293294
rect 30564 293058 30620 293294
rect 30272 292896 30620 293058
rect 166000 293294 166348 293456
rect 166000 293058 166056 293294
rect 166292 293058 166348 293294
rect 166000 292896 166348 293058
rect 25514 286718 25546 286954
rect 25782 286718 25866 286954
rect 26102 286718 26134 286954
rect 25514 266954 26134 286718
rect 30952 283294 31300 283456
rect 30952 283058 31008 283294
rect 31244 283058 31300 283294
rect 30952 282896 31300 283058
rect 165320 283294 165668 283456
rect 165320 283058 165376 283294
rect 165612 283058 165668 283294
rect 165320 282896 165668 283058
rect 30272 273294 30620 273456
rect 30272 273058 30328 273294
rect 30564 273058 30620 273294
rect 30272 272896 30620 273058
rect 166000 273294 166348 273456
rect 166000 273058 166056 273294
rect 166292 273058 166348 273294
rect 166000 272896 166348 273058
rect 25514 266718 25546 266954
rect 25782 266718 25866 266954
rect 26102 266718 26134 266954
rect 25514 246954 26134 266718
rect 30952 263294 31300 263456
rect 30952 263058 31008 263294
rect 31244 263058 31300 263294
rect 30952 262896 31300 263058
rect 165320 263294 165668 263456
rect 165320 263058 165376 263294
rect 165612 263058 165668 263294
rect 165320 262896 165668 263058
rect 43200 253330 43260 254106
rect 43336 253605 43396 254106
rect 60608 253741 60668 254106
rect 60605 253740 60671 253741
rect 60605 253676 60606 253740
rect 60670 253676 60671 253740
rect 60605 253675 60671 253676
rect 43333 253604 43399 253605
rect 43333 253540 43334 253604
rect 43398 253540 43399 253604
rect 43333 253539 43399 253540
rect 63192 253330 63252 254106
rect 65640 253741 65700 254106
rect 65637 253740 65703 253741
rect 65637 253676 65638 253740
rect 65702 253676 65703 253740
rect 65637 253675 65703 253676
rect 43118 253270 43260 253330
rect 63174 253270 63252 253330
rect 68088 253330 68148 254106
rect 70672 253741 70732 254106
rect 70669 253740 70735 253741
rect 70669 253676 70670 253740
rect 70734 253676 70735 253740
rect 70669 253675 70735 253676
rect 73120 253330 73180 254106
rect 75568 253741 75628 254106
rect 75565 253740 75631 253741
rect 75565 253676 75566 253740
rect 75630 253676 75631 253740
rect 75565 253675 75631 253676
rect 68088 253270 68202 253330
rect 43118 252381 43178 253270
rect 63174 252517 63234 253270
rect 68142 252517 68202 253270
rect 73110 253270 73180 253330
rect 78016 253330 78076 254106
rect 80600 253330 80660 254106
rect 83048 254010 83108 254106
rect 83046 253950 83108 254010
rect 78016 253270 78138 253330
rect 80600 253270 80714 253330
rect 73110 252517 73170 253270
rect 78078 252517 78138 253270
rect 80654 252517 80714 253270
rect 83046 252517 83106 253950
rect 85632 253330 85692 254106
rect 85622 253270 85692 253330
rect 88080 253330 88140 254106
rect 90664 253330 90724 254106
rect 93112 253330 93172 254106
rect 95560 254010 95620 254106
rect 95558 253950 95620 254010
rect 88080 253270 88258 253330
rect 90664 253270 90834 253330
rect 93112 253270 93226 253330
rect 85622 252517 85682 253270
rect 88198 252517 88258 253270
rect 90774 252517 90834 253270
rect 93166 252517 93226 253270
rect 95558 252517 95618 253950
rect 98280 253741 98340 254106
rect 98277 253740 98343 253741
rect 98277 253676 98278 253740
rect 98342 253676 98343 253740
rect 98277 253675 98343 253676
rect 100592 253330 100652 254106
rect 100526 253270 100652 253330
rect 103040 253330 103100 254106
rect 105624 253738 105684 254106
rect 107392 253738 107452 254106
rect 108072 253738 108132 254106
rect 108480 253738 108540 254106
rect 109568 253738 109628 254106
rect 110520 253738 110580 254106
rect 105624 253678 105738 253738
rect 103040 253270 103162 253330
rect 100526 252517 100586 253270
rect 103102 252517 103162 253270
rect 105678 252517 105738 253678
rect 107334 253678 107452 253738
rect 108070 253678 108132 253738
rect 108438 253678 108540 253738
rect 109542 253678 109628 253738
rect 110462 253678 110580 253738
rect 110792 253738 110852 254106
rect 112152 253738 112212 254106
rect 110792 253678 110890 253738
rect 63171 252516 63237 252517
rect 63171 252452 63172 252516
rect 63236 252452 63237 252516
rect 63171 252451 63237 252452
rect 68139 252516 68205 252517
rect 68139 252452 68140 252516
rect 68204 252452 68205 252516
rect 68139 252451 68205 252452
rect 73107 252516 73173 252517
rect 73107 252452 73108 252516
rect 73172 252452 73173 252516
rect 73107 252451 73173 252452
rect 78075 252516 78141 252517
rect 78075 252452 78076 252516
rect 78140 252452 78141 252516
rect 78075 252451 78141 252452
rect 80651 252516 80717 252517
rect 80651 252452 80652 252516
rect 80716 252452 80717 252516
rect 80651 252451 80717 252452
rect 83043 252516 83109 252517
rect 83043 252452 83044 252516
rect 83108 252452 83109 252516
rect 83043 252451 83109 252452
rect 85619 252516 85685 252517
rect 85619 252452 85620 252516
rect 85684 252452 85685 252516
rect 85619 252451 85685 252452
rect 88195 252516 88261 252517
rect 88195 252452 88196 252516
rect 88260 252452 88261 252516
rect 88195 252451 88261 252452
rect 90771 252516 90837 252517
rect 90771 252452 90772 252516
rect 90836 252452 90837 252516
rect 90771 252451 90837 252452
rect 93163 252516 93229 252517
rect 93163 252452 93164 252516
rect 93228 252452 93229 252516
rect 93163 252451 93229 252452
rect 95555 252516 95621 252517
rect 95555 252452 95556 252516
rect 95620 252452 95621 252516
rect 95555 252451 95621 252452
rect 100523 252516 100589 252517
rect 100523 252452 100524 252516
rect 100588 252452 100589 252516
rect 100523 252451 100589 252452
rect 103099 252516 103165 252517
rect 103099 252452 103100 252516
rect 103164 252452 103165 252516
rect 103099 252451 103165 252452
rect 105675 252516 105741 252517
rect 105675 252452 105676 252516
rect 105740 252452 105741 252516
rect 105675 252451 105741 252452
rect 43115 252380 43181 252381
rect 43115 252316 43116 252380
rect 43180 252316 43181 252380
rect 43115 252315 43181 252316
rect 25514 246718 25546 246954
rect 25782 246718 25866 246954
rect 26102 246718 26134 246954
rect 25514 226954 26134 246718
rect 29234 250614 29854 252000
rect 29234 250378 29266 250614
rect 29502 250378 29586 250614
rect 29822 250378 29854 250614
rect 29234 230614 29854 250378
rect 29234 230378 29266 230614
rect 29502 230378 29586 230614
rect 29822 230378 29854 230614
rect 29234 227308 29854 230378
rect 31794 233294 32414 252000
rect 31794 233058 31826 233294
rect 32062 233058 32146 233294
rect 32382 233058 32414 233294
rect 31794 227308 32414 233058
rect 32954 234274 33574 252000
rect 32954 234038 32986 234274
rect 33222 234038 33306 234274
rect 33542 234038 33574 234274
rect 32954 227308 33574 234038
rect 35514 236954 36134 252000
rect 35514 236718 35546 236954
rect 35782 236718 35866 236954
rect 36102 236718 36134 236954
rect 35203 227764 35269 227765
rect 35203 227700 35204 227764
rect 35268 227700 35269 227764
rect 35203 227699 35269 227700
rect 25514 226718 25546 226954
rect 25782 226718 25866 226954
rect 26102 226718 26134 226954
rect 25514 206954 26134 226718
rect 35206 225450 35266 227699
rect 35514 227308 36134 236718
rect 39234 240614 39854 252000
rect 39234 240378 39266 240614
rect 39502 240378 39586 240614
rect 39822 240378 39854 240614
rect 39234 227308 39854 240378
rect 41794 243294 42414 252000
rect 41794 243058 41826 243294
rect 42062 243058 42146 243294
rect 42382 243058 42414 243294
rect 41794 227308 42414 243058
rect 42954 244274 43574 252000
rect 42954 244038 42986 244274
rect 43222 244038 43306 244274
rect 43542 244038 43574 244274
rect 42954 227308 43574 244038
rect 45514 246954 46134 252000
rect 45514 246718 45546 246954
rect 45782 246718 45866 246954
rect 46102 246718 46134 246954
rect 45514 227308 46134 246718
rect 49234 250614 49854 252000
rect 49234 250378 49266 250614
rect 49502 250378 49586 250614
rect 49822 250378 49854 250614
rect 49234 230614 49854 250378
rect 49234 230378 49266 230614
rect 49502 230378 49586 230614
rect 49822 230378 49854 230614
rect 46795 227764 46861 227765
rect 46795 227700 46796 227764
rect 46860 227700 46861 227764
rect 46795 227699 46861 227700
rect 48083 227764 48149 227765
rect 48083 227700 48084 227764
rect 48148 227700 48149 227764
rect 48083 227699 48149 227700
rect 46798 225450 46858 227699
rect 48086 225450 48146 227699
rect 49234 227308 49854 230378
rect 51794 233294 52414 252000
rect 51794 233058 51826 233294
rect 52062 233058 52146 233294
rect 52382 233058 52414 233294
rect 51794 227308 52414 233058
rect 52954 234274 53574 252000
rect 52954 234038 52986 234274
rect 53222 234038 53306 234274
rect 53542 234038 53574 234274
rect 52954 227308 53574 234038
rect 55514 236954 56134 252000
rect 55514 236718 55546 236954
rect 55782 236718 55866 236954
rect 56102 236718 56134 236954
rect 55514 227308 56134 236718
rect 59234 240614 59854 252000
rect 59234 240378 59266 240614
rect 59502 240378 59586 240614
rect 59822 240378 59854 240614
rect 59234 227308 59854 240378
rect 61794 243294 62414 252000
rect 61794 243058 61826 243294
rect 62062 243058 62146 243294
rect 62382 243058 62414 243294
rect 61794 227308 62414 243058
rect 62954 244274 63574 252000
rect 62954 244038 62986 244274
rect 63222 244038 63306 244274
rect 63542 244038 63574 244274
rect 62954 227308 63574 244038
rect 65514 246954 66134 252000
rect 65514 246718 65546 246954
rect 65782 246718 65866 246954
rect 66102 246718 66134 246954
rect 65514 227308 66134 246718
rect 69234 250614 69854 252000
rect 69234 250378 69266 250614
rect 69502 250378 69586 250614
rect 69822 250378 69854 250614
rect 69234 230614 69854 250378
rect 69234 230378 69266 230614
rect 69502 230378 69586 230614
rect 69822 230378 69854 230614
rect 69234 227308 69854 230378
rect 71794 233294 72414 252000
rect 71794 233058 71826 233294
rect 72062 233058 72146 233294
rect 72382 233058 72414 233294
rect 71794 227308 72414 233058
rect 72954 234274 73574 252000
rect 72954 234038 72986 234274
rect 73222 234038 73306 234274
rect 73542 234038 73574 234274
rect 72954 227308 73574 234038
rect 75514 236954 76134 252000
rect 75514 236718 75546 236954
rect 75782 236718 75866 236954
rect 76102 236718 76134 236954
rect 75514 227308 76134 236718
rect 79234 240614 79854 252000
rect 79234 240378 79266 240614
rect 79502 240378 79586 240614
rect 79822 240378 79854 240614
rect 79234 227308 79854 240378
rect 81794 243294 82414 252000
rect 81794 243058 81826 243294
rect 82062 243058 82146 243294
rect 82382 243058 82414 243294
rect 81794 227308 82414 243058
rect 82954 244274 83574 252000
rect 82954 244038 82986 244274
rect 83222 244038 83306 244274
rect 83542 244038 83574 244274
rect 82954 227308 83574 244038
rect 85514 246954 86134 252000
rect 85514 246718 85546 246954
rect 85782 246718 85866 246954
rect 86102 246718 86134 246954
rect 85514 227308 86134 246718
rect 89234 250614 89854 252000
rect 89234 250378 89266 250614
rect 89502 250378 89586 250614
rect 89822 250378 89854 250614
rect 89234 230614 89854 250378
rect 89234 230378 89266 230614
rect 89502 230378 89586 230614
rect 89822 230378 89854 230614
rect 89234 227308 89854 230378
rect 91794 233294 92414 252000
rect 91794 233058 91826 233294
rect 92062 233058 92146 233294
rect 92382 233058 92414 233294
rect 91794 227308 92414 233058
rect 92954 234274 93574 252000
rect 92954 234038 92986 234274
rect 93222 234038 93306 234274
rect 93542 234038 93574 234274
rect 92954 227308 93574 234038
rect 95514 236954 96134 252000
rect 95514 236718 95546 236954
rect 95782 236718 95866 236954
rect 96102 236718 96134 236954
rect 95514 227308 96134 236718
rect 99234 240614 99854 252000
rect 99234 240378 99266 240614
rect 99502 240378 99586 240614
rect 99822 240378 99854 240614
rect 99234 227308 99854 240378
rect 101794 243294 102414 252000
rect 101794 243058 101826 243294
rect 102062 243058 102146 243294
rect 102382 243058 102414 243294
rect 101794 227308 102414 243058
rect 102954 244274 103574 252000
rect 102954 244038 102986 244274
rect 103222 244038 103306 244274
rect 103542 244038 103574 244274
rect 102954 227308 103574 244038
rect 105514 246954 106134 252000
rect 107334 251293 107394 253678
rect 108070 252517 108130 253678
rect 108067 252516 108133 252517
rect 108067 252452 108068 252516
rect 108132 252452 108133 252516
rect 108067 252451 108133 252452
rect 108438 251293 108498 253678
rect 109542 252381 109602 253678
rect 110462 252517 110522 253678
rect 110459 252516 110525 252517
rect 110459 252452 110460 252516
rect 110524 252452 110525 252516
rect 110459 252451 110525 252452
rect 110830 252381 110890 253678
rect 112118 253678 112212 253738
rect 112968 253738 113028 254106
rect 113240 253738 113300 254106
rect 114328 253738 114388 254106
rect 112968 253678 113098 253738
rect 112118 252381 112178 253678
rect 113038 252517 113098 253678
rect 113222 253678 113300 253738
rect 114326 253678 114388 253738
rect 115416 253738 115476 254106
rect 115552 253741 115612 254106
rect 115552 253740 115677 253741
rect 115416 253678 115490 253738
rect 115552 253678 115612 253740
rect 113035 252516 113101 252517
rect 113035 252452 113036 252516
rect 113100 252452 113101 252516
rect 113035 252451 113101 252452
rect 113222 252381 113282 253678
rect 109539 252380 109605 252381
rect 109539 252316 109540 252380
rect 109604 252316 109605 252380
rect 109539 252315 109605 252316
rect 110827 252380 110893 252381
rect 110827 252316 110828 252380
rect 110892 252316 110893 252380
rect 110827 252315 110893 252316
rect 112115 252380 112181 252381
rect 112115 252316 112116 252380
rect 112180 252316 112181 252380
rect 112115 252315 112181 252316
rect 113219 252380 113285 252381
rect 113219 252316 113220 252380
rect 113284 252316 113285 252380
rect 113219 252315 113285 252316
rect 107331 251292 107397 251293
rect 107331 251228 107332 251292
rect 107396 251228 107397 251292
rect 107331 251227 107397 251228
rect 108435 251292 108501 251293
rect 108435 251228 108436 251292
rect 108500 251228 108501 251292
rect 108435 251227 108501 251228
rect 105514 246718 105546 246954
rect 105782 246718 105866 246954
rect 106102 246718 106134 246954
rect 105514 227308 106134 246718
rect 109234 250614 109854 252000
rect 109234 250378 109266 250614
rect 109502 250378 109586 250614
rect 109822 250378 109854 250614
rect 109234 230614 109854 250378
rect 109234 230378 109266 230614
rect 109502 230378 109586 230614
rect 109822 230378 109854 230614
rect 109234 227308 109854 230378
rect 111794 233294 112414 252000
rect 111794 233058 111826 233294
rect 112062 233058 112146 233294
rect 112382 233058 112414 233294
rect 111794 227308 112414 233058
rect 112954 234274 113574 252000
rect 114326 251973 114386 253678
rect 115430 252517 115490 253678
rect 115611 253676 115612 253678
rect 115676 253676 115677 253740
rect 116776 253738 116836 254106
rect 117864 253738 117924 254106
rect 118272 253741 118332 254106
rect 115611 253675 115677 253676
rect 116718 253678 116836 253738
rect 117822 253678 117924 253738
rect 118269 253740 118335 253741
rect 115427 252516 115493 252517
rect 115427 252452 115428 252516
rect 115492 252452 115493 252516
rect 115427 252451 115493 252452
rect 114323 251972 114389 251973
rect 114323 251908 114324 251972
rect 114388 251908 114389 251972
rect 114323 251907 114389 251908
rect 112954 234038 112986 234274
rect 113222 234038 113306 234274
rect 113542 234038 113574 234274
rect 112954 227308 113574 234038
rect 115514 236954 116134 252000
rect 116718 251293 116778 253678
rect 117822 251293 117882 253678
rect 118269 253676 118270 253740
rect 118334 253676 118335 253740
rect 118952 253738 119012 254106
rect 118269 253675 118335 253676
rect 118926 253678 119012 253738
rect 120176 253738 120236 254106
rect 120584 253738 120644 254106
rect 120176 253678 120274 253738
rect 118926 251293 118986 253678
rect 116715 251292 116781 251293
rect 116715 251228 116716 251292
rect 116780 251228 116781 251292
rect 116715 251227 116781 251228
rect 117819 251292 117885 251293
rect 117819 251228 117820 251292
rect 117884 251228 117885 251292
rect 117819 251227 117885 251228
rect 118923 251292 118989 251293
rect 118923 251228 118924 251292
rect 118988 251228 118989 251292
rect 118923 251227 118989 251228
rect 115514 236718 115546 236954
rect 115782 236718 115866 236954
rect 116102 236718 116134 236954
rect 115514 227308 116134 236718
rect 119234 240614 119854 252000
rect 120214 251701 120274 253678
rect 120582 253678 120644 253738
rect 121264 253738 121324 254106
rect 122624 253738 122684 254106
rect 123032 253741 123092 254106
rect 121264 253678 121378 253738
rect 120582 252517 120642 253678
rect 120579 252516 120645 252517
rect 120579 252452 120580 252516
rect 120644 252452 120645 252516
rect 120579 252451 120645 252452
rect 120211 251700 120277 251701
rect 120211 251636 120212 251700
rect 120276 251636 120277 251700
rect 120211 251635 120277 251636
rect 121318 251293 121378 253678
rect 122606 253678 122684 253738
rect 123029 253740 123095 253741
rect 121315 251292 121381 251293
rect 121315 251228 121316 251292
rect 121380 251228 121381 251292
rect 121315 251227 121381 251228
rect 119234 240378 119266 240614
rect 119502 240378 119586 240614
rect 119822 240378 119854 240614
rect 119234 227308 119854 240378
rect 121794 243294 122414 252000
rect 122606 251293 122666 253678
rect 123029 253676 123030 253740
rect 123094 253676 123095 253740
rect 123712 253738 123772 254106
rect 123029 253675 123095 253676
rect 123710 253678 123772 253738
rect 124800 253738 124860 254106
rect 125480 253741 125540 254106
rect 125477 253740 125543 253741
rect 124800 253678 124874 253738
rect 122603 251292 122669 251293
rect 122603 251228 122604 251292
rect 122668 251228 122669 251292
rect 122603 251227 122669 251228
rect 121794 243058 121826 243294
rect 122062 243058 122146 243294
rect 122382 243058 122414 243294
rect 121794 227308 122414 243058
rect 122954 244274 123574 252000
rect 123710 251293 123770 253678
rect 124814 251293 124874 253678
rect 125477 253676 125478 253740
rect 125542 253676 125543 253740
rect 125888 253738 125948 254106
rect 127112 253738 127172 254106
rect 128064 253741 128124 254106
rect 128061 253740 128127 253741
rect 125888 253678 125978 253738
rect 127112 253678 127266 253738
rect 125477 253675 125543 253676
rect 125918 252381 125978 253678
rect 125915 252380 125981 252381
rect 125915 252316 125916 252380
rect 125980 252316 125981 252380
rect 125915 252315 125981 252316
rect 123707 251292 123773 251293
rect 123707 251228 123708 251292
rect 123772 251228 123773 251292
rect 123707 251227 123773 251228
rect 124811 251292 124877 251293
rect 124811 251228 124812 251292
rect 124876 251228 124877 251292
rect 124811 251227 124877 251228
rect 122954 244038 122986 244274
rect 123222 244038 123306 244274
rect 123542 244038 123574 244274
rect 122954 227308 123574 244038
rect 125514 246954 126134 252000
rect 127206 251293 127266 253678
rect 128061 253676 128062 253740
rect 128126 253676 128127 253740
rect 128472 253738 128532 254106
rect 129560 253738 129620 254106
rect 130512 253738 130572 254106
rect 130648 253738 130708 254106
rect 132008 253738 132068 254106
rect 132960 253738 133020 254106
rect 133096 254010 133156 254106
rect 128472 253678 128554 253738
rect 129560 253678 129658 253738
rect 130512 253678 130578 253738
rect 130648 253678 130762 253738
rect 128061 253675 128127 253676
rect 128494 251293 128554 253678
rect 129598 252381 129658 253678
rect 130518 253605 130578 253678
rect 130515 253604 130581 253605
rect 130515 253540 130516 253604
rect 130580 253540 130581 253604
rect 130515 253539 130581 253540
rect 129595 252380 129661 252381
rect 129595 252316 129596 252380
rect 129660 252316 129661 252380
rect 129595 252315 129661 252316
rect 127203 251292 127269 251293
rect 127203 251228 127204 251292
rect 127268 251228 127269 251292
rect 127203 251227 127269 251228
rect 128491 251292 128557 251293
rect 128491 251228 128492 251292
rect 128556 251228 128557 251292
rect 128491 251227 128557 251228
rect 125514 246718 125546 246954
rect 125782 246718 125866 246954
rect 126102 246718 126134 246954
rect 125514 227308 126134 246718
rect 129234 250614 129854 252000
rect 130702 251293 130762 253678
rect 131990 253678 132068 253738
rect 132910 253678 133020 253738
rect 133094 253950 133156 254010
rect 131990 252381 132050 253678
rect 132910 253469 132970 253678
rect 132907 253468 132973 253469
rect 132907 253404 132908 253468
rect 132972 253404 132973 253468
rect 132907 253403 132973 253404
rect 133094 252381 133154 253950
rect 134184 253738 134244 254106
rect 135272 253738 135332 254106
rect 135816 253738 135876 254106
rect 134184 253678 134258 253738
rect 135272 253678 135362 253738
rect 135816 253678 135914 253738
rect 131987 252380 132053 252381
rect 131987 252316 131988 252380
rect 132052 252316 132053 252380
rect 131987 252315 132053 252316
rect 133091 252380 133157 252381
rect 133091 252316 133092 252380
rect 133156 252316 133157 252380
rect 133091 252315 133157 252316
rect 130699 251292 130765 251293
rect 130699 251228 130700 251292
rect 130764 251228 130765 251292
rect 130699 251227 130765 251228
rect 129234 250378 129266 250614
rect 129502 250378 129586 250614
rect 129822 250378 129854 250614
rect 129234 230614 129854 250378
rect 129234 230378 129266 230614
rect 129502 230378 129586 230614
rect 129822 230378 129854 230614
rect 129234 227308 129854 230378
rect 131794 233294 132414 252000
rect 131794 233058 131826 233294
rect 132062 233058 132146 233294
rect 132382 233058 132414 233294
rect 131794 227308 132414 233058
rect 132954 234274 133574 252000
rect 134198 251293 134258 253678
rect 135302 251701 135362 253678
rect 135854 252517 135914 253678
rect 136496 253605 136556 254106
rect 137856 253738 137916 254106
rect 137856 253678 137938 253738
rect 136493 253604 136559 253605
rect 136493 253540 136494 253604
rect 136558 253540 136559 253604
rect 136493 253539 136559 253540
rect 135851 252516 135917 252517
rect 135851 252452 135852 252516
rect 135916 252452 135917 252516
rect 135851 252451 135917 252452
rect 135299 251700 135365 251701
rect 135299 251636 135300 251700
rect 135364 251636 135365 251700
rect 135299 251635 135365 251636
rect 134195 251292 134261 251293
rect 134195 251228 134196 251292
rect 134260 251228 134261 251292
rect 134195 251227 134261 251228
rect 132954 234038 132986 234274
rect 133222 234038 133306 234274
rect 133542 234038 133574 234274
rect 132954 227308 133574 234038
rect 135514 236954 136134 252000
rect 137878 251293 137938 253678
rect 138264 253330 138324 254106
rect 138246 253270 138324 253330
rect 138944 253330 139004 254106
rect 140032 253330 140092 254106
rect 141120 253330 141180 254106
rect 142344 253330 142404 254106
rect 143432 253330 143492 254106
rect 138944 253270 139042 253330
rect 140032 253270 140146 253330
rect 141120 253270 141250 253330
rect 138246 252381 138306 253270
rect 138243 252380 138309 252381
rect 138243 252316 138244 252380
rect 138308 252316 138309 252380
rect 138243 252315 138309 252316
rect 138982 251293 139042 253270
rect 137875 251292 137941 251293
rect 137875 251228 137876 251292
rect 137940 251228 137941 251292
rect 137875 251227 137941 251228
rect 138979 251292 139045 251293
rect 138979 251228 138980 251292
rect 139044 251228 139045 251292
rect 138979 251227 139045 251228
rect 135514 236718 135546 236954
rect 135782 236718 135866 236954
rect 136102 236718 136134 236954
rect 135514 227308 136134 236718
rect 139234 240614 139854 252000
rect 140086 251293 140146 253270
rect 141190 251973 141250 253270
rect 142294 253270 142404 253330
rect 143398 253270 143492 253330
rect 144792 253330 144852 254106
rect 146016 253330 146076 254106
rect 144792 253270 144930 253330
rect 142294 252381 142354 253270
rect 143398 252517 143458 253270
rect 144870 252517 144930 253270
rect 145974 253270 146076 253330
rect 146968 253330 147028 254106
rect 148328 253330 148388 254106
rect 149416 253330 149476 254106
rect 150504 253330 150564 254106
rect 146968 253270 147138 253330
rect 148328 253270 148426 253330
rect 149416 253270 150082 253330
rect 150504 253270 150634 253330
rect 145974 252517 146034 253270
rect 147078 252517 147138 253270
rect 148366 252517 148426 253270
rect 143395 252516 143461 252517
rect 143395 252452 143396 252516
rect 143460 252452 143461 252516
rect 143395 252451 143461 252452
rect 144867 252516 144933 252517
rect 144867 252452 144868 252516
rect 144932 252452 144933 252516
rect 144867 252451 144933 252452
rect 145971 252516 146037 252517
rect 145971 252452 145972 252516
rect 146036 252452 146037 252516
rect 145971 252451 146037 252452
rect 147075 252516 147141 252517
rect 147075 252452 147076 252516
rect 147140 252452 147141 252516
rect 147075 252451 147141 252452
rect 148363 252516 148429 252517
rect 148363 252452 148364 252516
rect 148428 252452 148429 252516
rect 148363 252451 148429 252452
rect 142291 252380 142357 252381
rect 142291 252316 142292 252380
rect 142356 252316 142357 252380
rect 142291 252315 142357 252316
rect 150022 252109 150082 253270
rect 150574 252517 150634 253270
rect 150571 252516 150637 252517
rect 150571 252452 150572 252516
rect 150636 252452 150637 252516
rect 150571 252451 150637 252452
rect 150019 252108 150085 252109
rect 150019 252044 150020 252108
rect 150084 252044 150085 252108
rect 150019 252043 150085 252044
rect 141187 251972 141253 251973
rect 141187 251908 141188 251972
rect 141252 251908 141253 251972
rect 141187 251907 141253 251908
rect 140083 251292 140149 251293
rect 140083 251228 140084 251292
rect 140148 251228 140149 251292
rect 140083 251227 140149 251228
rect 139234 240378 139266 240614
rect 139502 240378 139586 240614
rect 139822 240378 139854 240614
rect 139234 227308 139854 240378
rect 141794 243294 142414 252000
rect 141794 243058 141826 243294
rect 142062 243058 142146 243294
rect 142382 243058 142414 243294
rect 141794 227308 142414 243058
rect 142954 244274 143574 252000
rect 142954 244038 142986 244274
rect 143222 244038 143306 244274
rect 143542 244038 143574 244274
rect 142954 227308 143574 244038
rect 145514 246954 146134 252000
rect 145514 246718 145546 246954
rect 145782 246718 145866 246954
rect 146102 246718 146134 246954
rect 145514 227308 146134 246718
rect 149234 250614 149854 252000
rect 149234 250378 149266 250614
rect 149502 250378 149586 250614
rect 149822 250378 149854 250614
rect 149234 230614 149854 250378
rect 149234 230378 149266 230614
rect 149502 230378 149586 230614
rect 149822 230378 149854 230614
rect 149234 227308 149854 230378
rect 151794 233294 152414 252000
rect 151794 233058 151826 233294
rect 152062 233058 152146 233294
rect 152382 233058 152414 233294
rect 151794 227308 152414 233058
rect 152954 234274 153574 252000
rect 152954 234038 152986 234274
rect 153222 234038 153306 234274
rect 153542 234038 153574 234274
rect 152954 227308 153574 234038
rect 155514 236954 156134 252000
rect 155514 236718 155546 236954
rect 155782 236718 155866 236954
rect 156102 236718 156134 236954
rect 155514 227308 156134 236718
rect 159234 240614 159854 252000
rect 159234 240378 159266 240614
rect 159502 240378 159586 240614
rect 159822 240378 159854 240614
rect 159234 227308 159854 240378
rect 161794 243294 162414 252000
rect 161794 243058 161826 243294
rect 162062 243058 162146 243294
rect 162382 243058 162414 243294
rect 161794 227308 162414 243058
rect 162954 244274 163574 252000
rect 162954 244038 162986 244274
rect 163222 244038 163306 244274
rect 163542 244038 163574 244274
rect 162954 227308 163574 244038
rect 165514 246954 166134 252000
rect 165514 246718 165546 246954
rect 165782 246718 165866 246954
rect 166102 246718 166134 246954
rect 165514 227308 166134 246718
rect 167502 245717 167562 451827
rect 167686 421021 167746 581571
rect 167683 421020 167749 421021
rect 167683 420956 167684 421020
rect 167748 420956 167749 421020
rect 167683 420955 167749 420956
rect 168422 382397 168482 584835
rect 168603 581772 168669 581773
rect 168603 581708 168604 581772
rect 168668 581708 168669 581772
rect 168603 581707 168669 581708
rect 168606 448629 168666 581707
rect 169234 570614 169854 590378
rect 171794 705798 172414 705830
rect 171794 705562 171826 705798
rect 172062 705562 172146 705798
rect 172382 705562 172414 705798
rect 171794 705478 172414 705562
rect 171794 705242 171826 705478
rect 172062 705242 172146 705478
rect 172382 705242 172414 705478
rect 171794 693294 172414 705242
rect 171794 693058 171826 693294
rect 172062 693058 172146 693294
rect 172382 693058 172414 693294
rect 171794 673294 172414 693058
rect 171794 673058 171826 673294
rect 172062 673058 172146 673294
rect 172382 673058 172414 673294
rect 171794 653294 172414 673058
rect 171794 653058 171826 653294
rect 172062 653058 172146 653294
rect 172382 653058 172414 653294
rect 171794 633294 172414 653058
rect 171794 633058 171826 633294
rect 172062 633058 172146 633294
rect 172382 633058 172414 633294
rect 171794 613294 172414 633058
rect 171794 613058 171826 613294
rect 172062 613058 172146 613294
rect 172382 613058 172414 613294
rect 171794 593294 172414 613058
rect 171794 593058 171826 593294
rect 172062 593058 172146 593294
rect 172382 593058 172414 593294
rect 170075 587620 170141 587621
rect 170075 587556 170076 587620
rect 170140 587556 170141 587620
rect 170075 587555 170141 587556
rect 169234 570378 169266 570614
rect 169502 570378 169586 570614
rect 169822 570378 169854 570614
rect 169234 550614 169854 570378
rect 169234 550378 169266 550614
rect 169502 550378 169586 550614
rect 169822 550378 169854 550614
rect 169234 530614 169854 550378
rect 169234 530378 169266 530614
rect 169502 530378 169586 530614
rect 169822 530378 169854 530614
rect 169234 510614 169854 530378
rect 169234 510378 169266 510614
rect 169502 510378 169586 510614
rect 169822 510378 169854 510614
rect 169234 490614 169854 510378
rect 169234 490378 169266 490614
rect 169502 490378 169586 490614
rect 169822 490378 169854 490614
rect 169234 470614 169854 490378
rect 169234 470378 169266 470614
rect 169502 470378 169586 470614
rect 169822 470378 169854 470614
rect 168971 455836 169037 455837
rect 168971 455772 168972 455836
rect 169036 455772 169037 455836
rect 168971 455771 169037 455772
rect 168603 448628 168669 448629
rect 168603 448564 168604 448628
rect 168668 448564 168669 448628
rect 168603 448563 168669 448564
rect 168603 421020 168669 421021
rect 168603 420956 168604 421020
rect 168668 420956 168669 421020
rect 168603 420955 168669 420956
rect 168419 382396 168485 382397
rect 168419 382332 168420 382396
rect 168484 382332 168485 382396
rect 168419 382331 168485 382332
rect 168235 379540 168301 379541
rect 168235 379476 168236 379540
rect 168300 379476 168301 379540
rect 168235 379475 168301 379476
rect 168051 259588 168117 259589
rect 168051 259524 168052 259588
rect 168116 259524 168117 259588
rect 168051 259523 168117 259524
rect 168054 252245 168114 259523
rect 168051 252244 168117 252245
rect 168051 252180 168052 252244
rect 168116 252180 168117 252244
rect 168051 252179 168117 252180
rect 167499 245716 167565 245717
rect 167499 245652 167500 245716
rect 167564 245652 167565 245716
rect 167499 245651 167565 245652
rect 168238 238645 168298 379475
rect 168606 353293 168666 420955
rect 168603 353292 168669 353293
rect 168603 353228 168604 353292
rect 168668 353228 168669 353292
rect 168603 353227 168669 353228
rect 168606 352613 168666 353227
rect 168603 352612 168669 352613
rect 168603 352548 168604 352612
rect 168668 352548 168669 352612
rect 168603 352547 168669 352548
rect 168235 238644 168301 238645
rect 168235 238580 168236 238644
rect 168300 238580 168301 238644
rect 168235 238579 168301 238580
rect 168974 228989 169034 455771
rect 169234 450614 169854 470378
rect 169234 450378 169266 450614
rect 169502 450378 169586 450614
rect 169822 450378 169854 450614
rect 169234 430614 169854 450378
rect 169234 430378 169266 430614
rect 169502 430378 169586 430614
rect 169822 430378 169854 430614
rect 169234 410614 169854 430378
rect 170078 423605 170138 587555
rect 170259 587348 170325 587349
rect 170259 587284 170260 587348
rect 170324 587284 170325 587348
rect 170259 587283 170325 587284
rect 170262 460950 170322 587283
rect 171794 573294 172414 593058
rect 172954 694274 173574 710042
rect 182954 711558 183574 711590
rect 182954 711322 182986 711558
rect 183222 711322 183306 711558
rect 183542 711322 183574 711558
rect 182954 711238 183574 711322
rect 182954 711002 182986 711238
rect 183222 711002 183306 711238
rect 183542 711002 183574 711238
rect 179234 709638 179854 709670
rect 179234 709402 179266 709638
rect 179502 709402 179586 709638
rect 179822 709402 179854 709638
rect 179234 709318 179854 709402
rect 179234 709082 179266 709318
rect 179502 709082 179586 709318
rect 179822 709082 179854 709318
rect 175514 707718 176134 707750
rect 175514 707482 175546 707718
rect 175782 707482 175866 707718
rect 176102 707482 176134 707718
rect 175514 707398 176134 707482
rect 175514 707162 175546 707398
rect 175782 707162 175866 707398
rect 176102 707162 176134 707398
rect 174675 700500 174741 700501
rect 174675 700436 174676 700500
rect 174740 700436 174741 700500
rect 174675 700435 174741 700436
rect 174491 700364 174557 700365
rect 174491 700300 174492 700364
rect 174556 700300 174557 700364
rect 174491 700299 174557 700300
rect 172954 694038 172986 694274
rect 173222 694038 173306 694274
rect 173542 694038 173574 694274
rect 172954 674274 173574 694038
rect 172954 674038 172986 674274
rect 173222 674038 173306 674274
rect 173542 674038 173574 674274
rect 172954 654274 173574 674038
rect 172954 654038 172986 654274
rect 173222 654038 173306 654274
rect 173542 654038 173574 654274
rect 172954 634274 173574 654038
rect 172954 634038 172986 634274
rect 173222 634038 173306 634274
rect 173542 634038 173574 634274
rect 172954 614274 173574 634038
rect 172954 614038 172986 614274
rect 173222 614038 173306 614274
rect 173542 614038 173574 614274
rect 172954 594274 173574 614038
rect 172954 594038 172986 594274
rect 173222 594038 173306 594274
rect 173542 594038 173574 594274
rect 172651 584492 172717 584493
rect 172651 584428 172652 584492
rect 172716 584428 172717 584492
rect 172651 584427 172717 584428
rect 171794 573058 171826 573294
rect 172062 573058 172146 573294
rect 172382 573058 172414 573294
rect 171794 553294 172414 573058
rect 171794 553058 171826 553294
rect 172062 553058 172146 553294
rect 172382 553058 172414 553294
rect 171794 533294 172414 553058
rect 171794 533058 171826 533294
rect 172062 533058 172146 533294
rect 172382 533058 172414 533294
rect 171794 513294 172414 533058
rect 171794 513058 171826 513294
rect 172062 513058 172146 513294
rect 172382 513058 172414 513294
rect 171794 493294 172414 513058
rect 171794 493058 171826 493294
rect 172062 493058 172146 493294
rect 172382 493058 172414 493294
rect 171794 473294 172414 493058
rect 171794 473058 171826 473294
rect 172062 473058 172146 473294
rect 172382 473058 172414 473294
rect 170262 460890 170506 460950
rect 170446 451213 170506 460890
rect 171794 453294 172414 473058
rect 171794 453058 171826 453294
rect 172062 453058 172146 453294
rect 172382 453058 172414 453294
rect 170443 451212 170509 451213
rect 170443 451148 170444 451212
rect 170508 451148 170509 451212
rect 170443 451147 170509 451148
rect 170075 423604 170141 423605
rect 170075 423540 170076 423604
rect 170140 423540 170141 423604
rect 170075 423539 170141 423540
rect 170259 421156 170325 421157
rect 170259 421092 170260 421156
rect 170324 421092 170325 421156
rect 170259 421091 170325 421092
rect 169234 410378 169266 410614
rect 169502 410378 169586 410614
rect 169822 410378 169854 410614
rect 169234 390614 169854 410378
rect 169234 390378 169266 390614
rect 169502 390378 169586 390614
rect 169822 390378 169854 390614
rect 169234 370614 169854 390378
rect 169234 370378 169266 370614
rect 169502 370378 169586 370614
rect 169822 370378 169854 370614
rect 169234 350614 169854 370378
rect 169234 350378 169266 350614
rect 169502 350378 169586 350614
rect 169822 350378 169854 350614
rect 169234 330614 169854 350378
rect 169234 330378 169266 330614
rect 169502 330378 169586 330614
rect 169822 330378 169854 330614
rect 169234 310614 169854 330378
rect 169234 310378 169266 310614
rect 169502 310378 169586 310614
rect 169822 310378 169854 310614
rect 169234 290614 169854 310378
rect 169234 290378 169266 290614
rect 169502 290378 169586 290614
rect 169822 290378 169854 290614
rect 169234 270614 169854 290378
rect 169234 270378 169266 270614
rect 169502 270378 169586 270614
rect 169822 270378 169854 270614
rect 169234 250614 169854 270378
rect 169234 250378 169266 250614
rect 169502 250378 169586 250614
rect 169822 250378 169854 250614
rect 169234 230614 169854 250378
rect 169234 230378 169266 230614
rect 169502 230378 169586 230614
rect 169822 230378 169854 230614
rect 168971 228988 169037 228989
rect 168971 228924 168972 228988
rect 169036 228924 169037 228988
rect 168971 228923 169037 228924
rect 35206 225390 35780 225450
rect 46798 225390 46932 225450
rect 48086 225390 48156 225450
rect 35720 225202 35780 225390
rect 46872 225202 46932 225390
rect 48096 225202 48156 225390
rect 30952 223294 31300 223456
rect 30952 223058 31008 223294
rect 31244 223058 31300 223294
rect 30952 222896 31300 223058
rect 165320 223294 165668 223456
rect 165320 223058 165376 223294
rect 165612 223058 165668 223294
rect 165320 222896 165668 223058
rect 30272 213294 30620 213456
rect 30272 213058 30328 213294
rect 30564 213058 30620 213294
rect 30272 212896 30620 213058
rect 166000 213294 166348 213456
rect 166000 213058 166056 213294
rect 166292 213058 166348 213294
rect 166000 212896 166348 213058
rect 25514 206718 25546 206954
rect 25782 206718 25866 206954
rect 26102 206718 26134 206954
rect 25514 186954 26134 206718
rect 169234 210614 169854 230378
rect 170262 227085 170322 421091
rect 170446 361725 170506 451147
rect 171794 433294 172414 453058
rect 171794 433058 171826 433294
rect 172062 433058 172146 433294
rect 172382 433058 172414 433294
rect 170627 427684 170693 427685
rect 170627 427620 170628 427684
rect 170692 427620 170693 427684
rect 170627 427619 170693 427620
rect 170630 364037 170690 427619
rect 171547 421292 171613 421293
rect 171547 421228 171548 421292
rect 171612 421228 171613 421292
rect 171547 421227 171613 421228
rect 170627 364036 170693 364037
rect 170627 363972 170628 364036
rect 170692 363972 170693 364036
rect 170627 363971 170693 363972
rect 170443 361724 170509 361725
rect 170443 361660 170444 361724
rect 170508 361660 170509 361724
rect 170443 361659 170509 361660
rect 170259 227084 170325 227085
rect 170259 227020 170260 227084
rect 170324 227020 170325 227084
rect 170259 227019 170325 227020
rect 171550 226949 171610 421227
rect 171794 413294 172414 433058
rect 171794 413058 171826 413294
rect 172062 413058 172146 413294
rect 172382 413058 172414 413294
rect 171794 393294 172414 413058
rect 171794 393058 171826 393294
rect 172062 393058 172146 393294
rect 172382 393058 172414 393294
rect 171794 373294 172414 393058
rect 171794 373058 171826 373294
rect 172062 373058 172146 373294
rect 172382 373058 172414 373294
rect 171794 353294 172414 373058
rect 171794 353058 171826 353294
rect 172062 353058 172146 353294
rect 172382 353058 172414 353294
rect 171794 333294 172414 353058
rect 172654 342957 172714 584427
rect 172954 574274 173574 594038
rect 172954 574038 172986 574274
rect 173222 574038 173306 574274
rect 173542 574038 173574 574274
rect 172954 554274 173574 574038
rect 172954 554038 172986 554274
rect 173222 554038 173306 554274
rect 173542 554038 173574 554274
rect 172954 534274 173574 554038
rect 172954 534038 172986 534274
rect 173222 534038 173306 534274
rect 173542 534038 173574 534274
rect 172954 514274 173574 534038
rect 172954 514038 172986 514274
rect 173222 514038 173306 514274
rect 173542 514038 173574 514274
rect 172954 494274 173574 514038
rect 172954 494038 172986 494274
rect 173222 494038 173306 494274
rect 173542 494038 173574 494274
rect 172954 474274 173574 494038
rect 172954 474038 172986 474274
rect 173222 474038 173306 474274
rect 173542 474038 173574 474274
rect 172954 454274 173574 474038
rect 172954 454038 172986 454274
rect 173222 454038 173306 454274
rect 173542 454038 173574 454274
rect 172954 434274 173574 454038
rect 174494 438157 174554 700299
rect 174678 447949 174738 700435
rect 175514 696954 176134 707162
rect 175514 696718 175546 696954
rect 175782 696718 175866 696954
rect 176102 696718 176134 696954
rect 175514 676954 176134 696718
rect 175514 676718 175546 676954
rect 175782 676718 175866 676954
rect 176102 676718 176134 676954
rect 175514 656954 176134 676718
rect 175514 656718 175546 656954
rect 175782 656718 175866 656954
rect 176102 656718 176134 656954
rect 175514 636954 176134 656718
rect 175514 636718 175546 636954
rect 175782 636718 175866 636954
rect 176102 636718 176134 636954
rect 175514 616954 176134 636718
rect 175514 616718 175546 616954
rect 175782 616718 175866 616954
rect 176102 616718 176134 616954
rect 175514 596954 176134 616718
rect 175514 596718 175546 596954
rect 175782 596718 175866 596954
rect 176102 596718 176134 596954
rect 175514 576954 176134 596718
rect 175514 576718 175546 576954
rect 175782 576718 175866 576954
rect 176102 576718 176134 576954
rect 175514 556954 176134 576718
rect 175514 556718 175546 556954
rect 175782 556718 175866 556954
rect 176102 556718 176134 556954
rect 175514 536954 176134 556718
rect 175514 536718 175546 536954
rect 175782 536718 175866 536954
rect 176102 536718 176134 536954
rect 175514 516954 176134 536718
rect 175514 516718 175546 516954
rect 175782 516718 175866 516954
rect 176102 516718 176134 516954
rect 175514 496954 176134 516718
rect 175514 496718 175546 496954
rect 175782 496718 175866 496954
rect 176102 496718 176134 496954
rect 175514 476954 176134 496718
rect 175514 476718 175546 476954
rect 175782 476718 175866 476954
rect 176102 476718 176134 476954
rect 175514 456954 176134 476718
rect 175514 456718 175546 456954
rect 175782 456718 175866 456954
rect 176102 456718 176134 456954
rect 174675 447948 174741 447949
rect 174675 447884 174676 447948
rect 174740 447884 174741 447948
rect 174675 447883 174741 447884
rect 174491 438156 174557 438157
rect 174491 438092 174492 438156
rect 174556 438092 174557 438156
rect 174491 438091 174557 438092
rect 172954 434038 172986 434274
rect 173222 434038 173306 434274
rect 173542 434038 173574 434274
rect 172954 414274 173574 434038
rect 175514 436954 176134 456718
rect 175514 436718 175546 436954
rect 175782 436718 175866 436954
rect 176102 436718 176134 436954
rect 174675 421020 174741 421021
rect 174675 420956 174676 421020
rect 174740 420956 174741 421020
rect 174675 420955 174741 420956
rect 174491 419660 174557 419661
rect 174491 419596 174492 419660
rect 174556 419596 174557 419660
rect 174491 419595 174557 419596
rect 172954 414038 172986 414274
rect 173222 414038 173306 414274
rect 173542 414038 173574 414274
rect 172954 394274 173574 414038
rect 172954 394038 172986 394274
rect 173222 394038 173306 394274
rect 173542 394038 173574 394274
rect 172954 374274 173574 394038
rect 172954 374038 172986 374274
rect 173222 374038 173306 374274
rect 173542 374038 173574 374274
rect 172954 354274 173574 374038
rect 172954 354038 172986 354274
rect 173222 354038 173306 354274
rect 173542 354038 173574 354274
rect 172651 342956 172717 342957
rect 172651 342892 172652 342956
rect 172716 342892 172717 342956
rect 172651 342891 172717 342892
rect 171794 333058 171826 333294
rect 172062 333058 172146 333294
rect 172382 333058 172414 333294
rect 171794 313294 172414 333058
rect 171794 313058 171826 313294
rect 172062 313058 172146 313294
rect 172382 313058 172414 313294
rect 171794 293294 172414 313058
rect 171794 293058 171826 293294
rect 172062 293058 172146 293294
rect 172382 293058 172414 293294
rect 171794 273294 172414 293058
rect 171794 273058 171826 273294
rect 172062 273058 172146 273294
rect 172382 273058 172414 273294
rect 171794 253294 172414 273058
rect 171794 253058 171826 253294
rect 172062 253058 172146 253294
rect 172382 253058 172414 253294
rect 171794 233294 172414 253058
rect 171794 233058 171826 233294
rect 172062 233058 172146 233294
rect 172382 233058 172414 233294
rect 171547 226948 171613 226949
rect 171547 226884 171548 226948
rect 171612 226884 171613 226948
rect 171547 226883 171613 226884
rect 169234 210378 169266 210614
rect 169502 210378 169586 210614
rect 169822 210378 169854 210614
rect 30952 203294 31300 203456
rect 30952 203058 31008 203294
rect 31244 203058 31300 203294
rect 30952 202896 31300 203058
rect 165320 203294 165668 203456
rect 165320 203058 165376 203294
rect 165612 203058 165668 203294
rect 165320 202896 165668 203058
rect 30272 193294 30620 193456
rect 30272 193058 30328 193294
rect 30564 193058 30620 193294
rect 30272 192896 30620 193058
rect 166000 193294 166348 193456
rect 166000 193058 166056 193294
rect 166292 193058 166348 193294
rect 166000 192896 166348 193058
rect 25514 186718 25546 186954
rect 25782 186718 25866 186954
rect 26102 186718 26134 186954
rect 25514 166954 26134 186718
rect 169234 190614 169854 210378
rect 169234 190378 169266 190614
rect 169502 190378 169586 190614
rect 169822 190378 169854 190614
rect 30952 183294 31300 183456
rect 30952 183058 31008 183294
rect 31244 183058 31300 183294
rect 30952 182896 31300 183058
rect 165320 183294 165668 183456
rect 165320 183058 165376 183294
rect 165612 183058 165668 183294
rect 165320 182896 165668 183058
rect 30272 173294 30620 173456
rect 30272 173058 30328 173294
rect 30564 173058 30620 173294
rect 30272 172896 30620 173058
rect 166000 173294 166348 173456
rect 166000 173058 166056 173294
rect 166292 173058 166348 173294
rect 166000 172896 166348 173058
rect 25514 166718 25546 166954
rect 25782 166718 25866 166954
rect 26102 166718 26134 166954
rect 25514 146954 26134 166718
rect 169234 170614 169854 190378
rect 169234 170378 169266 170614
rect 169502 170378 169586 170614
rect 169822 170378 169854 170614
rect 30952 163294 31300 163456
rect 30952 163058 31008 163294
rect 31244 163058 31300 163294
rect 30952 162896 31300 163058
rect 165320 163294 165668 163456
rect 165320 163058 165376 163294
rect 165612 163058 165668 163294
rect 165320 162896 165668 163058
rect 30272 153294 30620 153456
rect 30272 153058 30328 153294
rect 30564 153058 30620 153294
rect 30272 152896 30620 153058
rect 166000 153294 166348 153456
rect 166000 153058 166056 153294
rect 166292 153058 166348 153294
rect 166000 152896 166348 153058
rect 25514 146718 25546 146954
rect 25782 146718 25866 146954
rect 26102 146718 26134 146954
rect 25514 126954 26134 146718
rect 169234 150614 169854 170378
rect 169234 150378 169266 150614
rect 169502 150378 169586 150614
rect 169822 150378 169854 150614
rect 43200 141810 43260 142106
rect 43118 141750 43260 141810
rect 43336 141810 43396 142106
rect 60608 141810 60668 142106
rect 63192 141810 63252 142106
rect 43336 141750 43730 141810
rect 43118 140181 43178 141750
rect 43115 140180 43181 140181
rect 43115 140116 43116 140180
rect 43180 140116 43181 140180
rect 43115 140115 43181 140116
rect 25514 126718 25546 126954
rect 25782 126718 25866 126954
rect 26102 126718 26134 126954
rect 25514 106954 26134 126718
rect 29234 130614 29854 140000
rect 29234 130378 29266 130614
rect 29502 130378 29586 130614
rect 29822 130378 29854 130614
rect 29234 115308 29854 130378
rect 31794 133294 32414 140000
rect 31794 133058 31826 133294
rect 32062 133058 32146 133294
rect 32382 133058 32414 133294
rect 31794 115308 32414 133058
rect 32954 134274 33574 140000
rect 32954 134038 32986 134274
rect 33222 134038 33306 134274
rect 33542 134038 33574 134274
rect 32954 115308 33574 134038
rect 35514 136954 36134 140000
rect 35514 136718 35546 136954
rect 35782 136718 35866 136954
rect 36102 136718 36134 136954
rect 35203 117196 35269 117197
rect 35203 117132 35204 117196
rect 35268 117132 35269 117196
rect 35203 117131 35269 117132
rect 35206 113930 35266 117131
rect 35514 116954 36134 136718
rect 35514 116718 35546 116954
rect 35782 116718 35866 116954
rect 36102 116718 36134 116954
rect 35514 115308 36134 116718
rect 39234 120614 39854 140000
rect 39234 120378 39266 120614
rect 39502 120378 39586 120614
rect 39822 120378 39854 120614
rect 39234 115308 39854 120378
rect 41794 123294 42414 140000
rect 41794 123058 41826 123294
rect 42062 123058 42146 123294
rect 42382 123058 42414 123294
rect 41794 115308 42414 123058
rect 42954 124274 43574 140000
rect 43670 139365 43730 141750
rect 60598 141750 60668 141810
rect 63174 141750 63252 141810
rect 65640 141810 65700 142106
rect 68088 141810 68148 142106
rect 70672 141810 70732 142106
rect 73120 141810 73180 142106
rect 75568 141810 75628 142106
rect 65640 141750 65810 141810
rect 68088 141750 68202 141810
rect 70672 141750 70778 141810
rect 73120 141750 73722 141810
rect 43667 139364 43733 139365
rect 43667 139300 43668 139364
rect 43732 139300 43733 139364
rect 43667 139299 43733 139300
rect 42954 124038 42986 124274
rect 43222 124038 43306 124274
rect 43542 124038 43574 124274
rect 42954 115308 43574 124038
rect 45514 126954 46134 140000
rect 45514 126718 45546 126954
rect 45782 126718 45866 126954
rect 46102 126718 46134 126954
rect 45514 115308 46134 126718
rect 49234 130614 49854 140000
rect 49234 130378 49266 130614
rect 49502 130378 49586 130614
rect 49822 130378 49854 130614
rect 46795 117060 46861 117061
rect 46795 116996 46796 117060
rect 46860 116996 46861 117060
rect 46795 116995 46861 116996
rect 46798 113930 46858 116995
rect 48083 116788 48149 116789
rect 48083 116724 48084 116788
rect 48148 116724 48149 116788
rect 48083 116723 48149 116724
rect 48086 113930 48146 116723
rect 49234 115308 49854 130378
rect 51794 133294 52414 140000
rect 51794 133058 51826 133294
rect 52062 133058 52146 133294
rect 52382 133058 52414 133294
rect 51794 115308 52414 133058
rect 52954 134274 53574 140000
rect 52954 134038 52986 134274
rect 53222 134038 53306 134274
rect 53542 134038 53574 134274
rect 52954 115308 53574 134038
rect 55514 136954 56134 140000
rect 55514 136718 55546 136954
rect 55782 136718 55866 136954
rect 56102 136718 56134 136954
rect 55514 116954 56134 136718
rect 55514 116718 55546 116954
rect 55782 116718 55866 116954
rect 56102 116718 56134 116954
rect 55514 115308 56134 116718
rect 59234 120614 59854 140000
rect 60598 139365 60658 141750
rect 63174 140181 63234 141750
rect 65750 140181 65810 141750
rect 63171 140180 63237 140181
rect 63171 140116 63172 140180
rect 63236 140116 63237 140180
rect 63171 140115 63237 140116
rect 65747 140180 65813 140181
rect 65747 140116 65748 140180
rect 65812 140116 65813 140180
rect 65747 140115 65813 140116
rect 60595 139364 60661 139365
rect 60595 139300 60596 139364
rect 60660 139300 60661 139364
rect 60595 139299 60661 139300
rect 59234 120378 59266 120614
rect 59502 120378 59586 120614
rect 59822 120378 59854 120614
rect 59234 115308 59854 120378
rect 61794 123294 62414 140000
rect 61794 123058 61826 123294
rect 62062 123058 62146 123294
rect 62382 123058 62414 123294
rect 61794 115308 62414 123058
rect 62954 124274 63574 140000
rect 62954 124038 62986 124274
rect 63222 124038 63306 124274
rect 63542 124038 63574 124274
rect 62954 115308 63574 124038
rect 65514 126954 66134 140000
rect 68142 138685 68202 141750
rect 68139 138684 68205 138685
rect 68139 138620 68140 138684
rect 68204 138620 68205 138684
rect 68139 138619 68205 138620
rect 65514 126718 65546 126954
rect 65782 126718 65866 126954
rect 66102 126718 66134 126954
rect 65514 115308 66134 126718
rect 69234 130614 69854 140000
rect 70718 138141 70778 141750
rect 70715 138140 70781 138141
rect 70715 138076 70716 138140
rect 70780 138076 70781 138140
rect 70715 138075 70781 138076
rect 69234 130378 69266 130614
rect 69502 130378 69586 130614
rect 69822 130378 69854 130614
rect 69234 115308 69854 130378
rect 71794 133294 72414 140000
rect 71794 133058 71826 133294
rect 72062 133058 72146 133294
rect 72382 133058 72414 133294
rect 71794 115308 72414 133058
rect 72954 134274 73574 140000
rect 73662 138141 73722 141750
rect 75318 141750 75628 141810
rect 78016 141810 78076 142106
rect 80600 141810 80660 142106
rect 83048 141810 83108 142106
rect 85632 141810 85692 142106
rect 88080 141810 88140 142106
rect 90664 141810 90724 142106
rect 93112 141810 93172 142106
rect 95560 141810 95620 142106
rect 98280 141810 98340 142106
rect 100592 141810 100652 142106
rect 103040 141810 103100 142106
rect 105624 141810 105684 142106
rect 107392 141810 107452 142106
rect 108072 141810 108132 142106
rect 78016 141750 78138 141810
rect 80600 141750 80714 141810
rect 83048 141750 83842 141810
rect 85632 141750 86418 141810
rect 88080 141750 88258 141810
rect 90664 141750 90834 141810
rect 93112 141750 93778 141810
rect 95560 141750 96354 141810
rect 98280 141750 98378 141810
rect 75318 138141 75378 141750
rect 73659 138140 73725 138141
rect 73659 138076 73660 138140
rect 73724 138076 73725 138140
rect 73659 138075 73725 138076
rect 75315 138140 75381 138141
rect 75315 138076 75316 138140
rect 75380 138076 75381 138140
rect 75315 138075 75381 138076
rect 72954 134038 72986 134274
rect 73222 134038 73306 134274
rect 73542 134038 73574 134274
rect 72954 115308 73574 134038
rect 75514 136954 76134 140000
rect 78078 138141 78138 141750
rect 78075 138140 78141 138141
rect 78075 138076 78076 138140
rect 78140 138076 78141 138140
rect 78075 138075 78141 138076
rect 75514 136718 75546 136954
rect 75782 136718 75866 136954
rect 76102 136718 76134 136954
rect 75514 116954 76134 136718
rect 75514 116718 75546 116954
rect 75782 116718 75866 116954
rect 76102 116718 76134 116954
rect 75514 115308 76134 116718
rect 79234 120614 79854 140000
rect 80654 138141 80714 141750
rect 80651 138140 80717 138141
rect 80651 138076 80652 138140
rect 80716 138076 80717 138140
rect 80651 138075 80717 138076
rect 79234 120378 79266 120614
rect 79502 120378 79586 120614
rect 79822 120378 79854 120614
rect 79234 115308 79854 120378
rect 81794 123294 82414 140000
rect 81794 123058 81826 123294
rect 82062 123058 82146 123294
rect 82382 123058 82414 123294
rect 81794 115308 82414 123058
rect 82954 124274 83574 140000
rect 83782 138141 83842 141750
rect 83779 138140 83845 138141
rect 83779 138076 83780 138140
rect 83844 138076 83845 138140
rect 83779 138075 83845 138076
rect 82954 124038 82986 124274
rect 83222 124038 83306 124274
rect 83542 124038 83574 124274
rect 82954 115308 83574 124038
rect 85514 126954 86134 140000
rect 86358 138141 86418 141750
rect 88198 138141 88258 141750
rect 86355 138140 86421 138141
rect 86355 138076 86356 138140
rect 86420 138076 86421 138140
rect 86355 138075 86421 138076
rect 88195 138140 88261 138141
rect 88195 138076 88196 138140
rect 88260 138076 88261 138140
rect 88195 138075 88261 138076
rect 85514 126718 85546 126954
rect 85782 126718 85866 126954
rect 86102 126718 86134 126954
rect 85514 115308 86134 126718
rect 89234 130614 89854 140000
rect 90774 138141 90834 141750
rect 90771 138140 90837 138141
rect 90771 138076 90772 138140
rect 90836 138076 90837 138140
rect 90771 138075 90837 138076
rect 89234 130378 89266 130614
rect 89502 130378 89586 130614
rect 89822 130378 89854 130614
rect 89234 115308 89854 130378
rect 91794 133294 92414 140000
rect 91794 133058 91826 133294
rect 92062 133058 92146 133294
rect 92382 133058 92414 133294
rect 91794 115308 92414 133058
rect 92954 134274 93574 140000
rect 93718 138141 93778 141750
rect 93715 138140 93781 138141
rect 93715 138076 93716 138140
rect 93780 138076 93781 138140
rect 93715 138075 93781 138076
rect 92954 134038 92986 134274
rect 93222 134038 93306 134274
rect 93542 134038 93574 134274
rect 92954 115308 93574 134038
rect 95514 136954 96134 140000
rect 96294 138141 96354 141750
rect 98318 138141 98378 141750
rect 100526 141750 100652 141810
rect 102734 141750 103100 141810
rect 105310 141750 105684 141810
rect 107334 141750 107452 141810
rect 108070 141750 108132 141810
rect 96291 138140 96357 138141
rect 96291 138076 96292 138140
rect 96356 138076 96357 138140
rect 96291 138075 96357 138076
rect 98315 138140 98381 138141
rect 98315 138076 98316 138140
rect 98380 138076 98381 138140
rect 98315 138075 98381 138076
rect 95514 136718 95546 136954
rect 95782 136718 95866 136954
rect 96102 136718 96134 136954
rect 95514 116954 96134 136718
rect 95514 116718 95546 116954
rect 95782 116718 95866 116954
rect 96102 116718 96134 116954
rect 95514 115308 96134 116718
rect 99234 120614 99854 140000
rect 100526 138141 100586 141750
rect 100523 138140 100589 138141
rect 100523 138076 100524 138140
rect 100588 138076 100589 138140
rect 100523 138075 100589 138076
rect 99234 120378 99266 120614
rect 99502 120378 99586 120614
rect 99822 120378 99854 120614
rect 99234 115308 99854 120378
rect 101794 123294 102414 140000
rect 102734 138141 102794 141750
rect 102731 138140 102797 138141
rect 102731 138076 102732 138140
rect 102796 138076 102797 138140
rect 102731 138075 102797 138076
rect 101794 123058 101826 123294
rect 102062 123058 102146 123294
rect 102382 123058 102414 123294
rect 101794 115308 102414 123058
rect 102954 124274 103574 140000
rect 105310 138141 105370 141750
rect 105307 138140 105373 138141
rect 105307 138076 105308 138140
rect 105372 138076 105373 138140
rect 105307 138075 105373 138076
rect 102954 124038 102986 124274
rect 103222 124038 103306 124274
rect 103542 124038 103574 124274
rect 102954 115308 103574 124038
rect 105514 126954 106134 140000
rect 107334 139365 107394 141750
rect 107331 139364 107397 139365
rect 107331 139300 107332 139364
rect 107396 139300 107397 139364
rect 107331 139299 107397 139300
rect 108070 138141 108130 141750
rect 108480 141677 108540 142106
rect 109568 141810 109628 142106
rect 110520 141810 110580 142106
rect 109542 141750 109628 141810
rect 110462 141750 110580 141810
rect 110792 141810 110852 142106
rect 110792 141750 110890 141810
rect 108477 141676 108543 141677
rect 108477 141612 108478 141676
rect 108542 141612 108543 141676
rect 108477 141611 108543 141612
rect 109542 140725 109602 141750
rect 109539 140724 109605 140725
rect 109539 140660 109540 140724
rect 109604 140660 109605 140724
rect 109539 140659 109605 140660
rect 108067 138140 108133 138141
rect 108067 138076 108068 138140
rect 108132 138076 108133 138140
rect 108067 138075 108133 138076
rect 105514 126718 105546 126954
rect 105782 126718 105866 126954
rect 106102 126718 106134 126954
rect 105514 115308 106134 126718
rect 109234 130614 109854 140000
rect 110462 138141 110522 141750
rect 110830 139365 110890 141750
rect 112152 141677 112212 142106
rect 112968 141810 113028 142106
rect 113240 141810 113300 142106
rect 114328 141810 114388 142106
rect 112670 141750 113028 141810
rect 113222 141750 113300 141810
rect 114326 141750 114388 141810
rect 115416 141810 115476 142106
rect 115552 141810 115612 142106
rect 116776 141810 116836 142106
rect 117864 141810 117924 142106
rect 115416 141750 115490 141810
rect 115552 141750 115674 141810
rect 112149 141676 112215 141677
rect 112149 141612 112150 141676
rect 112214 141612 112215 141676
rect 112149 141611 112215 141612
rect 110827 139364 110893 139365
rect 110827 139300 110828 139364
rect 110892 139300 110893 139364
rect 110827 139299 110893 139300
rect 110459 138140 110525 138141
rect 110459 138076 110460 138140
rect 110524 138076 110525 138140
rect 110459 138075 110525 138076
rect 109234 130378 109266 130614
rect 109502 130378 109586 130614
rect 109822 130378 109854 130614
rect 109234 115308 109854 130378
rect 111794 133294 112414 140000
rect 112670 138141 112730 141750
rect 113222 140725 113282 141750
rect 113219 140724 113285 140725
rect 113219 140660 113220 140724
rect 113284 140660 113285 140724
rect 113219 140659 113285 140660
rect 112667 138140 112733 138141
rect 112667 138076 112668 138140
rect 112732 138076 112733 138140
rect 112667 138075 112733 138076
rect 111794 133058 111826 133294
rect 112062 133058 112146 133294
rect 112382 133058 112414 133294
rect 111794 115308 112414 133058
rect 112954 134274 113574 140000
rect 114326 139365 114386 141750
rect 115430 140181 115490 141750
rect 115614 140181 115674 141750
rect 116718 141750 116836 141810
rect 117822 141750 117924 141810
rect 118272 141810 118332 142106
rect 118952 141810 119012 142106
rect 118272 141750 118434 141810
rect 116718 140725 116778 141750
rect 116715 140724 116781 140725
rect 116715 140660 116716 140724
rect 116780 140660 116781 140724
rect 116715 140659 116781 140660
rect 115427 140180 115493 140181
rect 115427 140116 115428 140180
rect 115492 140116 115493 140180
rect 115427 140115 115493 140116
rect 115611 140180 115677 140181
rect 115611 140116 115612 140180
rect 115676 140116 115677 140180
rect 115611 140115 115677 140116
rect 114323 139364 114389 139365
rect 114323 139300 114324 139364
rect 114388 139300 114389 139364
rect 114323 139299 114389 139300
rect 112954 134038 112986 134274
rect 113222 134038 113306 134274
rect 113542 134038 113574 134274
rect 112954 115308 113574 134038
rect 115514 136954 116134 140000
rect 117822 139365 117882 141750
rect 117819 139364 117885 139365
rect 117819 139300 117820 139364
rect 117884 139300 117885 139364
rect 117819 139299 117885 139300
rect 118374 138141 118434 141750
rect 118926 141750 119012 141810
rect 120176 141810 120236 142106
rect 120584 141810 120644 142106
rect 120176 141750 120274 141810
rect 118926 140725 118986 141750
rect 118923 140724 118989 140725
rect 118923 140660 118924 140724
rect 118988 140660 118989 140724
rect 118923 140659 118989 140660
rect 118371 138140 118437 138141
rect 118371 138076 118372 138140
rect 118436 138076 118437 138140
rect 118371 138075 118437 138076
rect 115514 136718 115546 136954
rect 115782 136718 115866 136954
rect 116102 136718 116134 136954
rect 115514 116954 116134 136718
rect 115514 116718 115546 116954
rect 115782 116718 115866 116954
rect 116102 116718 116134 116954
rect 115514 115308 116134 116718
rect 119234 120614 119854 140000
rect 120214 139365 120274 141750
rect 120582 141750 120644 141810
rect 121264 141810 121324 142106
rect 122624 141810 122684 142106
rect 123032 141813 123092 142106
rect 121264 141750 121378 141810
rect 120211 139364 120277 139365
rect 120211 139300 120212 139364
rect 120276 139300 120277 139364
rect 120211 139299 120277 139300
rect 120582 138141 120642 141750
rect 121318 139365 121378 141750
rect 122606 141750 122684 141810
rect 123029 141812 123095 141813
rect 121315 139364 121381 139365
rect 121315 139300 121316 139364
rect 121380 139300 121381 139364
rect 121315 139299 121381 139300
rect 120579 138140 120645 138141
rect 120579 138076 120580 138140
rect 120644 138076 120645 138140
rect 120579 138075 120645 138076
rect 119234 120378 119266 120614
rect 119502 120378 119586 120614
rect 119822 120378 119854 120614
rect 119234 115308 119854 120378
rect 121794 123294 122414 140000
rect 122606 139365 122666 141750
rect 123029 141748 123030 141812
rect 123094 141748 123095 141812
rect 123029 141747 123095 141748
rect 123712 141677 123772 142106
rect 123709 141676 123775 141677
rect 123709 141612 123710 141676
rect 123774 141612 123775 141676
rect 124800 141674 124860 142106
rect 125480 141810 125540 142106
rect 125366 141750 125540 141810
rect 124800 141614 124874 141674
rect 123709 141611 123775 141612
rect 122603 139364 122669 139365
rect 122603 139300 122604 139364
rect 122668 139300 122669 139364
rect 122603 139299 122669 139300
rect 121794 123058 121826 123294
rect 122062 123058 122146 123294
rect 122382 123058 122414 123294
rect 121794 115308 122414 123058
rect 122954 124274 123574 140000
rect 124814 139365 124874 141614
rect 124811 139364 124877 139365
rect 124811 139300 124812 139364
rect 124876 139300 124877 139364
rect 124811 139299 124877 139300
rect 125366 138141 125426 141750
rect 125888 141674 125948 142106
rect 127112 141810 127172 142106
rect 127112 141750 127266 141810
rect 125888 141614 125978 141674
rect 125918 140725 125978 141614
rect 125915 140724 125981 140725
rect 125915 140660 125916 140724
rect 125980 140660 125981 140724
rect 125915 140659 125981 140660
rect 125363 138140 125429 138141
rect 125363 138076 125364 138140
rect 125428 138076 125429 138140
rect 125363 138075 125429 138076
rect 122954 124038 122986 124274
rect 123222 124038 123306 124274
rect 123542 124038 123574 124274
rect 122954 115308 123574 124038
rect 125514 126954 126134 140000
rect 127206 139365 127266 141750
rect 128064 141674 128124 142106
rect 128472 141677 128532 142106
rect 128469 141676 128535 141677
rect 128064 141614 128186 141674
rect 127203 139364 127269 139365
rect 127203 139300 127204 139364
rect 127268 139300 127269 139364
rect 127203 139299 127269 139300
rect 128126 138141 128186 141614
rect 128469 141612 128470 141676
rect 128534 141612 128535 141676
rect 129560 141674 129620 142106
rect 130512 141674 130572 142106
rect 130648 141674 130708 142106
rect 132008 141674 132068 142106
rect 132960 141674 133020 142106
rect 133096 141813 133156 142106
rect 133093 141812 133159 141813
rect 133093 141748 133094 141812
rect 133158 141748 133159 141812
rect 133093 141747 133159 141748
rect 134184 141677 134244 142106
rect 129560 141614 129658 141674
rect 130512 141614 130578 141674
rect 130648 141614 130762 141674
rect 128469 141611 128535 141612
rect 129598 140181 129658 141614
rect 129595 140180 129661 140181
rect 129595 140116 129596 140180
rect 129660 140116 129661 140180
rect 129595 140115 129661 140116
rect 128123 138140 128189 138141
rect 128123 138076 128124 138140
rect 128188 138076 128189 138140
rect 128123 138075 128189 138076
rect 125514 126718 125546 126954
rect 125782 126718 125866 126954
rect 126102 126718 126134 126954
rect 125514 115308 126134 126718
rect 129234 130614 129854 140000
rect 130518 138141 130578 141614
rect 130702 139365 130762 141614
rect 131990 141614 132068 141674
rect 132726 141614 133020 141674
rect 134181 141676 134247 141677
rect 131990 140725 132050 141614
rect 131987 140724 132053 140725
rect 131987 140660 131988 140724
rect 132052 140660 132053 140724
rect 131987 140659 132053 140660
rect 130699 139364 130765 139365
rect 130699 139300 130700 139364
rect 130764 139300 130765 139364
rect 130699 139299 130765 139300
rect 130515 138140 130581 138141
rect 130515 138076 130516 138140
rect 130580 138076 130581 138140
rect 130515 138075 130581 138076
rect 129234 130378 129266 130614
rect 129502 130378 129586 130614
rect 129822 130378 129854 130614
rect 129234 115308 129854 130378
rect 131794 133294 132414 140000
rect 132726 138141 132786 141614
rect 134181 141612 134182 141676
rect 134246 141612 134247 141676
rect 135272 141674 135332 142106
rect 135816 141674 135876 142106
rect 136496 141677 136556 142106
rect 136493 141676 136559 141677
rect 135272 141614 135362 141674
rect 135816 141614 136282 141674
rect 134181 141611 134247 141612
rect 135302 140725 135362 141614
rect 135299 140724 135365 140725
rect 135299 140660 135300 140724
rect 135364 140660 135365 140724
rect 135299 140659 135365 140660
rect 132723 138140 132789 138141
rect 132723 138076 132724 138140
rect 132788 138076 132789 138140
rect 132723 138075 132789 138076
rect 131794 133058 131826 133294
rect 132062 133058 132146 133294
rect 132382 133058 132414 133294
rect 131794 115308 132414 133058
rect 132954 134274 133574 140000
rect 132954 134038 132986 134274
rect 133222 134038 133306 134274
rect 133542 134038 133574 134274
rect 132954 115308 133574 134038
rect 135514 136954 136134 140000
rect 136222 139093 136282 141614
rect 136493 141612 136494 141676
rect 136558 141612 136559 141676
rect 137856 141674 137916 142106
rect 138264 141674 138324 142106
rect 137856 141614 137938 141674
rect 136493 141611 136559 141612
rect 137878 140725 137938 141614
rect 138246 141614 138324 141674
rect 138944 141674 139004 142106
rect 140032 141677 140092 142106
rect 141120 141810 141180 142106
rect 141120 141750 141250 141810
rect 140029 141676 140095 141677
rect 138944 141614 139042 141674
rect 137875 140724 137941 140725
rect 137875 140660 137876 140724
rect 137940 140660 137941 140724
rect 137875 140659 137941 140660
rect 136219 139092 136285 139093
rect 136219 139028 136220 139092
rect 136284 139028 136285 139092
rect 136219 139027 136285 139028
rect 138246 138141 138306 141614
rect 138982 140725 139042 141614
rect 140029 141612 140030 141676
rect 140094 141612 140095 141676
rect 140029 141611 140095 141612
rect 141190 140725 141250 141750
rect 142344 141677 142404 142106
rect 143432 141810 143492 142106
rect 143398 141750 143492 141810
rect 144792 141810 144852 142106
rect 146016 141810 146076 142106
rect 146968 141810 147028 142106
rect 148328 141810 148388 142106
rect 149416 141810 149476 142106
rect 150504 141810 150564 142106
rect 144792 141750 148426 141810
rect 149416 141750 149530 141810
rect 150504 141750 150634 141810
rect 142341 141676 142407 141677
rect 142341 141612 142342 141676
rect 142406 141612 142407 141676
rect 142341 141611 142407 141612
rect 143398 140725 143458 141750
rect 138979 140724 139045 140725
rect 138979 140660 138980 140724
rect 139044 140660 139045 140724
rect 138979 140659 139045 140660
rect 141187 140724 141253 140725
rect 141187 140660 141188 140724
rect 141252 140660 141253 140724
rect 141187 140659 141253 140660
rect 143395 140724 143461 140725
rect 143395 140660 143396 140724
rect 143460 140660 143461 140724
rect 143395 140659 143461 140660
rect 138243 138140 138309 138141
rect 138243 138076 138244 138140
rect 138308 138076 138309 138140
rect 138243 138075 138309 138076
rect 135514 136718 135546 136954
rect 135782 136718 135866 136954
rect 136102 136718 136134 136954
rect 135514 116954 136134 136718
rect 135514 116718 135546 116954
rect 135782 116718 135866 116954
rect 136102 116718 136134 116954
rect 135514 115308 136134 116718
rect 139234 120614 139854 140000
rect 139234 120378 139266 120614
rect 139502 120378 139586 120614
rect 139822 120378 139854 120614
rect 139234 115308 139854 120378
rect 141794 123294 142414 140000
rect 141794 123058 141826 123294
rect 142062 123058 142146 123294
rect 142382 123058 142414 123294
rect 141794 115308 142414 123058
rect 142954 124274 143574 140000
rect 142954 124038 142986 124274
rect 143222 124038 143306 124274
rect 143542 124038 143574 124274
rect 142954 115308 143574 124038
rect 145514 126954 146134 140000
rect 148366 139365 148426 141750
rect 149470 140725 149530 141750
rect 149467 140724 149533 140725
rect 149467 140660 149468 140724
rect 149532 140660 149533 140724
rect 149467 140659 149533 140660
rect 148363 139364 148429 139365
rect 148363 139300 148364 139364
rect 148428 139300 148429 139364
rect 148363 139299 148429 139300
rect 145514 126718 145546 126954
rect 145782 126718 145866 126954
rect 146102 126718 146134 126954
rect 145514 115308 146134 126718
rect 149234 130614 149854 140000
rect 150574 139365 150634 141750
rect 150571 139364 150637 139365
rect 150571 139300 150572 139364
rect 150636 139300 150637 139364
rect 150571 139299 150637 139300
rect 149234 130378 149266 130614
rect 149502 130378 149586 130614
rect 149822 130378 149854 130614
rect 149234 115308 149854 130378
rect 151794 133294 152414 140000
rect 151794 133058 151826 133294
rect 152062 133058 152146 133294
rect 152382 133058 152414 133294
rect 151794 115308 152414 133058
rect 152954 134274 153574 140000
rect 152954 134038 152986 134274
rect 153222 134038 153306 134274
rect 153542 134038 153574 134274
rect 152954 115308 153574 134038
rect 155514 136954 156134 140000
rect 155514 136718 155546 136954
rect 155782 136718 155866 136954
rect 156102 136718 156134 136954
rect 155514 116954 156134 136718
rect 155514 116718 155546 116954
rect 155782 116718 155866 116954
rect 156102 116718 156134 116954
rect 155514 115308 156134 116718
rect 159234 120614 159854 140000
rect 159234 120378 159266 120614
rect 159502 120378 159586 120614
rect 159822 120378 159854 120614
rect 159234 115308 159854 120378
rect 161794 123294 162414 140000
rect 161794 123058 161826 123294
rect 162062 123058 162146 123294
rect 162382 123058 162414 123294
rect 161794 115308 162414 123058
rect 162954 124274 163574 140000
rect 162954 124038 162986 124274
rect 163222 124038 163306 124274
rect 163542 124038 163574 124274
rect 162954 115308 163574 124038
rect 165514 126954 166134 140000
rect 165514 126718 165546 126954
rect 165782 126718 165866 126954
rect 166102 126718 166134 126954
rect 165514 115308 166134 126718
rect 169234 130614 169854 150378
rect 169234 130378 169266 130614
rect 169502 130378 169586 130614
rect 169822 130378 169854 130614
rect 35206 113870 35780 113930
rect 46798 113870 46932 113930
rect 48086 113870 48156 113930
rect 35720 113220 35780 113870
rect 46872 113220 46932 113870
rect 48096 113220 48156 113870
rect 25514 106718 25546 106954
rect 25782 106718 25866 106954
rect 26102 106718 26134 106954
rect 25514 86954 26134 106718
rect 169234 110614 169854 130378
rect 169234 110378 169266 110614
rect 169502 110378 169586 110614
rect 169822 110378 169854 110614
rect 30952 103294 31300 103456
rect 30952 103058 31008 103294
rect 31244 103058 31300 103294
rect 30952 102896 31300 103058
rect 165320 103294 165668 103456
rect 165320 103058 165376 103294
rect 165612 103058 165668 103294
rect 165320 102896 165668 103058
rect 30272 93294 30620 93456
rect 30272 93058 30328 93294
rect 30564 93058 30620 93294
rect 30272 92896 30620 93058
rect 166000 93294 166348 93456
rect 166000 93058 166056 93294
rect 166292 93058 166348 93294
rect 166000 92896 166348 93058
rect 25514 86718 25546 86954
rect 25782 86718 25866 86954
rect 26102 86718 26134 86954
rect 25514 66954 26134 86718
rect 169234 90614 169854 110378
rect 169234 90378 169266 90614
rect 169502 90378 169586 90614
rect 169822 90378 169854 90614
rect 30952 83294 31300 83456
rect 30952 83058 31008 83294
rect 31244 83058 31300 83294
rect 30952 82896 31300 83058
rect 165320 83294 165668 83456
rect 165320 83058 165376 83294
rect 165612 83058 165668 83294
rect 165320 82896 165668 83058
rect 30272 73294 30620 73456
rect 30272 73058 30328 73294
rect 30564 73058 30620 73294
rect 30272 72896 30620 73058
rect 166000 73294 166348 73456
rect 166000 73058 166056 73294
rect 166292 73058 166348 73294
rect 166000 72896 166348 73058
rect 25514 66718 25546 66954
rect 25782 66718 25866 66954
rect 26102 66718 26134 66954
rect 25514 46954 26134 66718
rect 169234 70614 169854 90378
rect 169234 70378 169266 70614
rect 169502 70378 169586 70614
rect 169822 70378 169854 70614
rect 30952 63294 31300 63456
rect 30952 63058 31008 63294
rect 31244 63058 31300 63294
rect 30952 62896 31300 63058
rect 165320 63294 165668 63456
rect 165320 63058 165376 63294
rect 165612 63058 165668 63294
rect 165320 62896 165668 63058
rect 30272 53294 30620 53456
rect 30272 53058 30328 53294
rect 30564 53058 30620 53294
rect 30272 52896 30620 53058
rect 166000 53294 166348 53456
rect 166000 53058 166056 53294
rect 166292 53058 166348 53294
rect 166000 52896 166348 53058
rect 25514 46718 25546 46954
rect 25782 46718 25866 46954
rect 26102 46718 26134 46954
rect 25514 26954 26134 46718
rect 169234 50614 169854 70378
rect 169234 50378 169266 50614
rect 169502 50378 169586 50614
rect 169822 50378 169854 50614
rect 30952 43294 31300 43456
rect 30952 43058 31008 43294
rect 31244 43058 31300 43294
rect 30952 42896 31300 43058
rect 165320 43294 165668 43456
rect 165320 43058 165376 43294
rect 165612 43058 165668 43294
rect 165320 42896 165668 43058
rect 30272 33294 30620 33456
rect 30272 33058 30328 33294
rect 30564 33058 30620 33294
rect 30272 32896 30620 33058
rect 166000 33294 166348 33456
rect 166000 33058 166056 33294
rect 166292 33058 166348 33294
rect 166000 32896 166348 33058
rect 169234 30614 169854 50378
rect 169234 30378 169266 30614
rect 169502 30378 169586 30614
rect 169822 30378 169854 30614
rect 43200 29610 43260 30106
rect 42750 29550 43260 29610
rect 43336 29610 43396 30106
rect 60608 29610 60668 30106
rect 63192 29610 63252 30106
rect 65640 29610 65700 30106
rect 43336 29550 43730 29610
rect 25514 26718 25546 26954
rect 25782 26718 25866 26954
rect 26102 26718 26134 26954
rect 25514 6954 26134 26718
rect 25514 6718 25546 6954
rect 25782 6718 25866 6954
rect 26102 6718 26134 6954
rect 25514 -2266 26134 6718
rect 25514 -2502 25546 -2266
rect 25782 -2502 25866 -2266
rect 26102 -2502 26134 -2266
rect 25514 -2586 26134 -2502
rect 25514 -2822 25546 -2586
rect 25782 -2822 25866 -2586
rect 26102 -2822 26134 -2586
rect 25514 -3814 26134 -2822
rect 29234 10614 29854 28000
rect 29234 10378 29266 10614
rect 29502 10378 29586 10614
rect 29822 10378 29854 10614
rect 29234 -4186 29854 10378
rect 31794 13294 32414 28000
rect 31794 13058 31826 13294
rect 32062 13058 32146 13294
rect 32382 13058 32414 13294
rect 31794 -1306 32414 13058
rect 31794 -1542 31826 -1306
rect 32062 -1542 32146 -1306
rect 32382 -1542 32414 -1306
rect 31794 -1626 32414 -1542
rect 31794 -1862 31826 -1626
rect 32062 -1862 32146 -1626
rect 32382 -1862 32414 -1626
rect 31794 -1894 32414 -1862
rect 32954 14274 33574 28000
rect 32954 14038 32986 14274
rect 33222 14038 33306 14274
rect 33542 14038 33574 14274
rect 29234 -4422 29266 -4186
rect 29502 -4422 29586 -4186
rect 29822 -4422 29854 -4186
rect 29234 -4506 29854 -4422
rect 29234 -4742 29266 -4506
rect 29502 -4742 29586 -4506
rect 29822 -4742 29854 -4506
rect 29234 -5734 29854 -4742
rect 22954 -7302 22986 -7066
rect 23222 -7302 23306 -7066
rect 23542 -7302 23574 -7066
rect 22954 -7386 23574 -7302
rect 22954 -7622 22986 -7386
rect 23222 -7622 23306 -7386
rect 23542 -7622 23574 -7386
rect 22954 -7654 23574 -7622
rect 32954 -6106 33574 14038
rect 35514 16954 36134 28000
rect 35514 16718 35546 16954
rect 35782 16718 35866 16954
rect 36102 16718 36134 16954
rect 35514 -3226 36134 16718
rect 35514 -3462 35546 -3226
rect 35782 -3462 35866 -3226
rect 36102 -3462 36134 -3226
rect 35514 -3546 36134 -3462
rect 35514 -3782 35546 -3546
rect 35782 -3782 35866 -3546
rect 36102 -3782 36134 -3546
rect 35514 -3814 36134 -3782
rect 39234 20614 39854 28000
rect 39234 20378 39266 20614
rect 39502 20378 39586 20614
rect 39822 20378 39854 20614
rect 39234 -5146 39854 20378
rect 41794 23294 42414 28000
rect 42750 27573 42810 29550
rect 42747 27572 42813 27573
rect 42747 27508 42748 27572
rect 42812 27508 42813 27572
rect 42747 27507 42813 27508
rect 41794 23058 41826 23294
rect 42062 23058 42146 23294
rect 42382 23058 42414 23294
rect 41794 3294 42414 23058
rect 41794 3058 41826 3294
rect 42062 3058 42146 3294
rect 42382 3058 42414 3294
rect 41794 -346 42414 3058
rect 41794 -582 41826 -346
rect 42062 -582 42146 -346
rect 42382 -582 42414 -346
rect 41794 -666 42414 -582
rect 41794 -902 41826 -666
rect 42062 -902 42146 -666
rect 42382 -902 42414 -666
rect 41794 -1894 42414 -902
rect 42954 24274 43574 28000
rect 43670 27573 43730 29550
rect 60598 29550 60668 29610
rect 63174 29550 63252 29610
rect 65566 29550 65700 29610
rect 68088 29610 68148 30106
rect 70672 29610 70732 30106
rect 73120 29610 73180 30106
rect 75568 29613 75628 30106
rect 75565 29612 75631 29613
rect 68088 29550 68202 29610
rect 70672 29550 70778 29610
rect 73120 29550 73722 29610
rect 60598 28933 60658 29550
rect 60595 28932 60661 28933
rect 60595 28868 60596 28932
rect 60660 28868 60661 28932
rect 60595 28867 60661 28868
rect 63174 28253 63234 29550
rect 65566 29010 65626 29550
rect 64646 28950 65626 29010
rect 63171 28252 63237 28253
rect 63171 28188 63172 28252
rect 63236 28188 63237 28252
rect 63171 28187 63237 28188
rect 43667 27572 43733 27573
rect 43667 27508 43668 27572
rect 43732 27508 43733 27572
rect 43667 27507 43733 27508
rect 42954 24038 42986 24274
rect 43222 24038 43306 24274
rect 43542 24038 43574 24274
rect 39234 -5382 39266 -5146
rect 39502 -5382 39586 -5146
rect 39822 -5382 39854 -5146
rect 39234 -5466 39854 -5382
rect 39234 -5702 39266 -5466
rect 39502 -5702 39586 -5466
rect 39822 -5702 39854 -5466
rect 39234 -5734 39854 -5702
rect 32954 -6342 32986 -6106
rect 33222 -6342 33306 -6106
rect 33542 -6342 33574 -6106
rect 32954 -6426 33574 -6342
rect 32954 -6662 32986 -6426
rect 33222 -6662 33306 -6426
rect 33542 -6662 33574 -6426
rect 32954 -7654 33574 -6662
rect 42954 -7066 43574 24038
rect 45514 26954 46134 28000
rect 45514 26718 45546 26954
rect 45782 26718 45866 26954
rect 46102 26718 46134 26954
rect 45514 6954 46134 26718
rect 45514 6718 45546 6954
rect 45782 6718 45866 6954
rect 46102 6718 46134 6954
rect 45514 -2266 46134 6718
rect 45514 -2502 45546 -2266
rect 45782 -2502 45866 -2266
rect 46102 -2502 46134 -2266
rect 45514 -2586 46134 -2502
rect 45514 -2822 45546 -2586
rect 45782 -2822 45866 -2586
rect 46102 -2822 46134 -2586
rect 45514 -3814 46134 -2822
rect 49234 10614 49854 28000
rect 49234 10378 49266 10614
rect 49502 10378 49586 10614
rect 49822 10378 49854 10614
rect 49234 -4186 49854 10378
rect 51794 13294 52414 28000
rect 51794 13058 51826 13294
rect 52062 13058 52146 13294
rect 52382 13058 52414 13294
rect 51794 -1306 52414 13058
rect 51794 -1542 51826 -1306
rect 52062 -1542 52146 -1306
rect 52382 -1542 52414 -1306
rect 51794 -1626 52414 -1542
rect 51794 -1862 51826 -1626
rect 52062 -1862 52146 -1626
rect 52382 -1862 52414 -1626
rect 51794 -1894 52414 -1862
rect 52954 14274 53574 28000
rect 52954 14038 52986 14274
rect 53222 14038 53306 14274
rect 53542 14038 53574 14274
rect 49234 -4422 49266 -4186
rect 49502 -4422 49586 -4186
rect 49822 -4422 49854 -4186
rect 49234 -4506 49854 -4422
rect 49234 -4742 49266 -4506
rect 49502 -4742 49586 -4506
rect 49822 -4742 49854 -4506
rect 49234 -5734 49854 -4742
rect 42954 -7302 42986 -7066
rect 43222 -7302 43306 -7066
rect 43542 -7302 43574 -7066
rect 42954 -7386 43574 -7302
rect 42954 -7622 42986 -7386
rect 43222 -7622 43306 -7386
rect 43542 -7622 43574 -7386
rect 42954 -7654 43574 -7622
rect 52954 -6106 53574 14038
rect 55514 16954 56134 28000
rect 55514 16718 55546 16954
rect 55782 16718 55866 16954
rect 56102 16718 56134 16954
rect 55514 -3226 56134 16718
rect 55514 -3462 55546 -3226
rect 55782 -3462 55866 -3226
rect 56102 -3462 56134 -3226
rect 55514 -3546 56134 -3462
rect 55514 -3782 55546 -3546
rect 55782 -3782 55866 -3546
rect 56102 -3782 56134 -3546
rect 55514 -3814 56134 -3782
rect 59234 20614 59854 28000
rect 59234 20378 59266 20614
rect 59502 20378 59586 20614
rect 59822 20378 59854 20614
rect 59234 -5146 59854 20378
rect 61794 23294 62414 28000
rect 61794 23058 61826 23294
rect 62062 23058 62146 23294
rect 62382 23058 62414 23294
rect 61794 3294 62414 23058
rect 61794 3058 61826 3294
rect 62062 3058 62146 3294
rect 62382 3058 62414 3294
rect 61794 -346 62414 3058
rect 61794 -582 61826 -346
rect 62062 -582 62146 -346
rect 62382 -582 62414 -346
rect 61794 -666 62414 -582
rect 61794 -902 61826 -666
rect 62062 -902 62146 -666
rect 62382 -902 62414 -666
rect 61794 -1894 62414 -902
rect 62954 24274 63574 28000
rect 64646 27570 64706 28950
rect 68142 28933 68202 29550
rect 68139 28932 68205 28933
rect 68139 28868 68140 28932
rect 68204 28868 68205 28932
rect 68139 28867 68205 28868
rect 64827 27572 64893 27573
rect 64827 27570 64828 27572
rect 64646 27510 64828 27570
rect 64827 27508 64828 27510
rect 64892 27508 64893 27572
rect 64827 27507 64893 27508
rect 62954 24038 62986 24274
rect 63222 24038 63306 24274
rect 63542 24038 63574 24274
rect 59234 -5382 59266 -5146
rect 59502 -5382 59586 -5146
rect 59822 -5382 59854 -5146
rect 59234 -5466 59854 -5382
rect 59234 -5702 59266 -5466
rect 59502 -5702 59586 -5466
rect 59822 -5702 59854 -5466
rect 59234 -5734 59854 -5702
rect 52954 -6342 52986 -6106
rect 53222 -6342 53306 -6106
rect 53542 -6342 53574 -6106
rect 52954 -6426 53574 -6342
rect 52954 -6662 52986 -6426
rect 53222 -6662 53306 -6426
rect 53542 -6662 53574 -6426
rect 52954 -7654 53574 -6662
rect 62954 -7066 63574 24038
rect 65514 26954 66134 28000
rect 65514 26718 65546 26954
rect 65782 26718 65866 26954
rect 66102 26718 66134 26954
rect 65514 6954 66134 26718
rect 65514 6718 65546 6954
rect 65782 6718 65866 6954
rect 66102 6718 66134 6954
rect 65514 -2266 66134 6718
rect 65514 -2502 65546 -2266
rect 65782 -2502 65866 -2266
rect 66102 -2502 66134 -2266
rect 65514 -2586 66134 -2502
rect 65514 -2822 65546 -2586
rect 65782 -2822 65866 -2586
rect 66102 -2822 66134 -2586
rect 65514 -3814 66134 -2822
rect 69234 10614 69854 28000
rect 70718 27573 70778 29550
rect 70715 27572 70781 27573
rect 70715 27508 70716 27572
rect 70780 27508 70781 27572
rect 70715 27507 70781 27508
rect 69234 10378 69266 10614
rect 69502 10378 69586 10614
rect 69822 10378 69854 10614
rect 69234 -4186 69854 10378
rect 71794 13294 72414 28000
rect 71794 13058 71826 13294
rect 72062 13058 72146 13294
rect 72382 13058 72414 13294
rect 71794 -1306 72414 13058
rect 71794 -1542 71826 -1306
rect 72062 -1542 72146 -1306
rect 72382 -1542 72414 -1306
rect 71794 -1626 72414 -1542
rect 71794 -1862 71826 -1626
rect 72062 -1862 72146 -1626
rect 72382 -1862 72414 -1626
rect 71794 -1894 72414 -1862
rect 72954 14274 73574 28000
rect 73662 27573 73722 29550
rect 75565 29548 75566 29612
rect 75630 29548 75631 29612
rect 78016 29610 78076 30106
rect 80600 29610 80660 30106
rect 83048 29610 83108 30106
rect 78016 29550 78138 29610
rect 80600 29550 80714 29610
rect 75565 29547 75631 29548
rect 78078 28933 78138 29550
rect 80654 28933 80714 29550
rect 83046 29550 83108 29610
rect 85632 29610 85692 30106
rect 88080 29613 88140 30106
rect 90664 29613 90724 30106
rect 88077 29612 88143 29613
rect 85632 29550 86418 29610
rect 83046 28933 83106 29550
rect 78075 28932 78141 28933
rect 78075 28868 78076 28932
rect 78140 28868 78141 28932
rect 78075 28867 78141 28868
rect 80651 28932 80717 28933
rect 80651 28868 80652 28932
rect 80716 28868 80717 28932
rect 80651 28867 80717 28868
rect 83043 28932 83109 28933
rect 83043 28868 83044 28932
rect 83108 28868 83109 28932
rect 83043 28867 83109 28868
rect 73659 27572 73725 27573
rect 73659 27508 73660 27572
rect 73724 27508 73725 27572
rect 73659 27507 73725 27508
rect 72954 14038 72986 14274
rect 73222 14038 73306 14274
rect 73542 14038 73574 14274
rect 69234 -4422 69266 -4186
rect 69502 -4422 69586 -4186
rect 69822 -4422 69854 -4186
rect 69234 -4506 69854 -4422
rect 69234 -4742 69266 -4506
rect 69502 -4742 69586 -4506
rect 69822 -4742 69854 -4506
rect 69234 -5734 69854 -4742
rect 62954 -7302 62986 -7066
rect 63222 -7302 63306 -7066
rect 63542 -7302 63574 -7066
rect 62954 -7386 63574 -7302
rect 62954 -7622 62986 -7386
rect 63222 -7622 63306 -7386
rect 63542 -7622 63574 -7386
rect 62954 -7654 63574 -7622
rect 72954 -6106 73574 14038
rect 75514 16954 76134 28000
rect 75514 16718 75546 16954
rect 75782 16718 75866 16954
rect 76102 16718 76134 16954
rect 75514 -3226 76134 16718
rect 75514 -3462 75546 -3226
rect 75782 -3462 75866 -3226
rect 76102 -3462 76134 -3226
rect 75514 -3546 76134 -3462
rect 75514 -3782 75546 -3546
rect 75782 -3782 75866 -3546
rect 76102 -3782 76134 -3546
rect 75514 -3814 76134 -3782
rect 79234 20614 79854 28000
rect 79234 20378 79266 20614
rect 79502 20378 79586 20614
rect 79822 20378 79854 20614
rect 79234 -5146 79854 20378
rect 81794 23294 82414 28000
rect 81794 23058 81826 23294
rect 82062 23058 82146 23294
rect 82382 23058 82414 23294
rect 81794 3294 82414 23058
rect 81794 3058 81826 3294
rect 82062 3058 82146 3294
rect 82382 3058 82414 3294
rect 81794 -346 82414 3058
rect 81794 -582 81826 -346
rect 82062 -582 82146 -346
rect 82382 -582 82414 -346
rect 81794 -666 82414 -582
rect 81794 -902 81826 -666
rect 82062 -902 82146 -666
rect 82382 -902 82414 -666
rect 81794 -1894 82414 -902
rect 82954 24274 83574 28000
rect 82954 24038 82986 24274
rect 83222 24038 83306 24274
rect 83542 24038 83574 24274
rect 79234 -5382 79266 -5146
rect 79502 -5382 79586 -5146
rect 79822 -5382 79854 -5146
rect 79234 -5466 79854 -5382
rect 79234 -5702 79266 -5466
rect 79502 -5702 79586 -5466
rect 79822 -5702 79854 -5466
rect 79234 -5734 79854 -5702
rect 72954 -6342 72986 -6106
rect 73222 -6342 73306 -6106
rect 73542 -6342 73574 -6106
rect 72954 -6426 73574 -6342
rect 72954 -6662 72986 -6426
rect 73222 -6662 73306 -6426
rect 73542 -6662 73574 -6426
rect 72954 -7654 73574 -6662
rect 82954 -7066 83574 24038
rect 85514 26954 86134 28000
rect 86358 27573 86418 29550
rect 88077 29548 88078 29612
rect 88142 29548 88143 29612
rect 88077 29547 88143 29548
rect 90661 29612 90727 29613
rect 90661 29548 90662 29612
rect 90726 29548 90727 29612
rect 93112 29610 93172 30106
rect 95560 29610 95620 30106
rect 90661 29547 90727 29548
rect 92798 29550 93172 29610
rect 95374 29550 95620 29610
rect 98280 29610 98340 30106
rect 100592 29610 100652 30106
rect 98280 29550 98378 29610
rect 86355 27572 86421 27573
rect 86355 27508 86356 27572
rect 86420 27508 86421 27572
rect 86355 27507 86421 27508
rect 85514 26718 85546 26954
rect 85782 26718 85866 26954
rect 86102 26718 86134 26954
rect 85514 6954 86134 26718
rect 85514 6718 85546 6954
rect 85782 6718 85866 6954
rect 86102 6718 86134 6954
rect 85514 -2266 86134 6718
rect 85514 -2502 85546 -2266
rect 85782 -2502 85866 -2266
rect 86102 -2502 86134 -2266
rect 85514 -2586 86134 -2502
rect 85514 -2822 85546 -2586
rect 85782 -2822 85866 -2586
rect 86102 -2822 86134 -2586
rect 85514 -3814 86134 -2822
rect 89234 10614 89854 28000
rect 89234 10378 89266 10614
rect 89502 10378 89586 10614
rect 89822 10378 89854 10614
rect 89234 -4186 89854 10378
rect 91794 13294 92414 28000
rect 92798 27573 92858 29550
rect 92795 27572 92861 27573
rect 92795 27508 92796 27572
rect 92860 27508 92861 27572
rect 92795 27507 92861 27508
rect 91794 13058 91826 13294
rect 92062 13058 92146 13294
rect 92382 13058 92414 13294
rect 91794 -1306 92414 13058
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 92954 14274 93574 28000
rect 95187 27572 95253 27573
rect 95187 27508 95188 27572
rect 95252 27570 95253 27572
rect 95374 27570 95434 29550
rect 95252 27510 95434 27570
rect 95252 27508 95253 27510
rect 95187 27507 95253 27508
rect 92954 14038 92986 14274
rect 93222 14038 93306 14274
rect 93542 14038 93574 14274
rect 89234 -4422 89266 -4186
rect 89502 -4422 89586 -4186
rect 89822 -4422 89854 -4186
rect 89234 -4506 89854 -4422
rect 89234 -4742 89266 -4506
rect 89502 -4742 89586 -4506
rect 89822 -4742 89854 -4506
rect 89234 -5734 89854 -4742
rect 82954 -7302 82986 -7066
rect 83222 -7302 83306 -7066
rect 83542 -7302 83574 -7066
rect 82954 -7386 83574 -7302
rect 82954 -7622 82986 -7386
rect 83222 -7622 83306 -7386
rect 83542 -7622 83574 -7386
rect 82954 -7654 83574 -7622
rect 92954 -6106 93574 14038
rect 95514 16954 96134 28000
rect 98318 27573 98378 29550
rect 100526 29550 100652 29610
rect 103040 29610 103100 30106
rect 105624 29610 105684 30106
rect 107392 29610 107452 30106
rect 108072 29610 108132 30106
rect 108480 29610 108540 30106
rect 103040 29550 103162 29610
rect 98315 27572 98381 27573
rect 98315 27508 98316 27572
rect 98380 27508 98381 27572
rect 98315 27507 98381 27508
rect 95514 16718 95546 16954
rect 95782 16718 95866 16954
rect 96102 16718 96134 16954
rect 95514 -3226 96134 16718
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 20614 99854 28000
rect 100526 27573 100586 29550
rect 103102 28933 103162 29550
rect 105310 29550 105684 29610
rect 107334 29550 107452 29610
rect 108070 29550 108132 29610
rect 108438 29550 108540 29610
rect 109568 29610 109628 30106
rect 110520 29610 110580 30106
rect 109568 29550 110154 29610
rect 103099 28932 103165 28933
rect 103099 28868 103100 28932
rect 103164 28868 103165 28932
rect 103099 28867 103165 28868
rect 100523 27572 100589 27573
rect 100523 27508 100524 27572
rect 100588 27508 100589 27572
rect 100523 27507 100589 27508
rect 99234 20378 99266 20614
rect 99502 20378 99586 20614
rect 99822 20378 99854 20614
rect 99234 -5146 99854 20378
rect 101794 23294 102414 28000
rect 101794 23058 101826 23294
rect 102062 23058 102146 23294
rect 102382 23058 102414 23294
rect 101794 3294 102414 23058
rect 101794 3058 101826 3294
rect 102062 3058 102146 3294
rect 102382 3058 102414 3294
rect 101794 -346 102414 3058
rect 101794 -582 101826 -346
rect 102062 -582 102146 -346
rect 102382 -582 102414 -346
rect 101794 -666 102414 -582
rect 101794 -902 101826 -666
rect 102062 -902 102146 -666
rect 102382 -902 102414 -666
rect 101794 -1894 102414 -902
rect 102954 24274 103574 28000
rect 105310 27573 105370 29550
rect 105307 27572 105373 27573
rect 105307 27508 105308 27572
rect 105372 27508 105373 27572
rect 105307 27507 105373 27508
rect 102954 24038 102986 24274
rect 103222 24038 103306 24274
rect 103542 24038 103574 24274
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 92954 -6342 92986 -6106
rect 93222 -6342 93306 -6106
rect 93542 -6342 93574 -6106
rect 92954 -6426 93574 -6342
rect 92954 -6662 92986 -6426
rect 93222 -6662 93306 -6426
rect 93542 -6662 93574 -6426
rect 92954 -7654 93574 -6662
rect 102954 -7066 103574 24038
rect 105514 26954 106134 28000
rect 107334 27573 107394 29550
rect 108070 27573 108130 29550
rect 108438 27573 108498 29550
rect 107331 27572 107397 27573
rect 107331 27508 107332 27572
rect 107396 27508 107397 27572
rect 107331 27507 107397 27508
rect 108067 27572 108133 27573
rect 108067 27508 108068 27572
rect 108132 27508 108133 27572
rect 108067 27507 108133 27508
rect 108435 27572 108501 27573
rect 108435 27508 108436 27572
rect 108500 27508 108501 27572
rect 108435 27507 108501 27508
rect 105514 26718 105546 26954
rect 105782 26718 105866 26954
rect 106102 26718 106134 26954
rect 105514 6954 106134 26718
rect 105514 6718 105546 6954
rect 105782 6718 105866 6954
rect 106102 6718 106134 6954
rect 105514 -2266 106134 6718
rect 105514 -2502 105546 -2266
rect 105782 -2502 105866 -2266
rect 106102 -2502 106134 -2266
rect 105514 -2586 106134 -2502
rect 105514 -2822 105546 -2586
rect 105782 -2822 105866 -2586
rect 106102 -2822 106134 -2586
rect 105514 -3814 106134 -2822
rect 109234 10614 109854 28000
rect 110094 27573 110154 29550
rect 110462 29550 110580 29610
rect 110792 29610 110852 30106
rect 112152 29610 112212 30106
rect 112968 29610 113028 30106
rect 110792 29550 110890 29610
rect 110091 27572 110157 27573
rect 110091 27508 110092 27572
rect 110156 27508 110157 27572
rect 110091 27507 110157 27508
rect 110462 27437 110522 29550
rect 110830 27573 110890 29550
rect 112118 29550 112212 29610
rect 112670 29550 113028 29610
rect 113240 29610 113300 30106
rect 114328 29610 114388 30106
rect 115416 29610 115476 30106
rect 113240 29550 113834 29610
rect 112118 28253 112178 29550
rect 112115 28252 112181 28253
rect 112115 28188 112116 28252
rect 112180 28188 112181 28252
rect 112115 28187 112181 28188
rect 110827 27572 110893 27573
rect 110827 27508 110828 27572
rect 110892 27508 110893 27572
rect 110827 27507 110893 27508
rect 110459 27436 110525 27437
rect 110459 27372 110460 27436
rect 110524 27372 110525 27436
rect 110459 27371 110525 27372
rect 109234 10378 109266 10614
rect 109502 10378 109586 10614
rect 109822 10378 109854 10614
rect 109234 -4186 109854 10378
rect 111794 13294 112414 28000
rect 112670 27573 112730 29550
rect 112667 27572 112733 27573
rect 112667 27508 112668 27572
rect 112732 27508 112733 27572
rect 112667 27507 112733 27508
rect 111794 13058 111826 13294
rect 112062 13058 112146 13294
rect 112382 13058 112414 13294
rect 111794 -1306 112414 13058
rect 111794 -1542 111826 -1306
rect 112062 -1542 112146 -1306
rect 112382 -1542 112414 -1306
rect 111794 -1626 112414 -1542
rect 111794 -1862 111826 -1626
rect 112062 -1862 112146 -1626
rect 112382 -1862 112414 -1626
rect 111794 -1894 112414 -1862
rect 112954 14274 113574 28000
rect 113774 27165 113834 29550
rect 114326 29550 114388 29610
rect 115246 29550 115476 29610
rect 115552 29610 115612 30106
rect 116776 29610 116836 30106
rect 117864 29610 117924 30106
rect 115552 29550 115674 29610
rect 113771 27164 113837 27165
rect 113771 27100 113772 27164
rect 113836 27100 113837 27164
rect 113771 27099 113837 27100
rect 114326 27029 114386 29550
rect 114323 27028 114389 27029
rect 114323 26964 114324 27028
rect 114388 26964 114389 27028
rect 114323 26963 114389 26964
rect 115246 26349 115306 29550
rect 115614 28253 115674 29550
rect 116718 29550 116836 29610
rect 117822 29550 117924 29610
rect 118272 29610 118332 30106
rect 118952 29610 119012 30106
rect 118272 29550 118434 29610
rect 115611 28252 115677 28253
rect 115611 28188 115612 28252
rect 115676 28188 115677 28252
rect 115611 28187 115677 28188
rect 115243 26348 115309 26349
rect 115243 26284 115244 26348
rect 115308 26284 115309 26348
rect 115243 26283 115309 26284
rect 112954 14038 112986 14274
rect 113222 14038 113306 14274
rect 113542 14038 113574 14274
rect 109234 -4422 109266 -4186
rect 109502 -4422 109586 -4186
rect 109822 -4422 109854 -4186
rect 109234 -4506 109854 -4422
rect 109234 -4742 109266 -4506
rect 109502 -4742 109586 -4506
rect 109822 -4742 109854 -4506
rect 109234 -5734 109854 -4742
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 112954 -6106 113574 14038
rect 115514 16954 116134 28000
rect 116718 27573 116778 29550
rect 117822 27573 117882 29550
rect 118374 27573 118434 29550
rect 118926 29550 119012 29610
rect 120176 29610 120236 30106
rect 120584 29610 120644 30106
rect 120176 29550 120274 29610
rect 116715 27572 116781 27573
rect 116715 27508 116716 27572
rect 116780 27508 116781 27572
rect 116715 27507 116781 27508
rect 117819 27572 117885 27573
rect 117819 27508 117820 27572
rect 117884 27508 117885 27572
rect 117819 27507 117885 27508
rect 118371 27572 118437 27573
rect 118371 27508 118372 27572
rect 118436 27508 118437 27572
rect 118371 27507 118437 27508
rect 118926 26349 118986 29550
rect 118923 26348 118989 26349
rect 118923 26284 118924 26348
rect 118988 26284 118989 26348
rect 118923 26283 118989 26284
rect 115514 16718 115546 16954
rect 115782 16718 115866 16954
rect 116102 16718 116134 16954
rect 115514 -3226 116134 16718
rect 115514 -3462 115546 -3226
rect 115782 -3462 115866 -3226
rect 116102 -3462 116134 -3226
rect 115514 -3546 116134 -3462
rect 115514 -3782 115546 -3546
rect 115782 -3782 115866 -3546
rect 116102 -3782 116134 -3546
rect 115514 -3814 116134 -3782
rect 119234 20614 119854 28000
rect 120214 27573 120274 29550
rect 120582 29550 120644 29610
rect 121264 29610 121324 30106
rect 122624 29610 122684 30106
rect 121264 29550 121378 29610
rect 120211 27572 120277 27573
rect 120211 27508 120212 27572
rect 120276 27508 120277 27572
rect 120211 27507 120277 27508
rect 120582 27301 120642 29550
rect 121318 27437 121378 29550
rect 122606 29550 122684 29610
rect 123032 29610 123092 30106
rect 123712 29613 123772 30106
rect 123709 29612 123775 29613
rect 123032 29550 123218 29610
rect 121315 27436 121381 27437
rect 121315 27372 121316 27436
rect 121380 27372 121381 27436
rect 121315 27371 121381 27372
rect 120579 27300 120645 27301
rect 120579 27236 120580 27300
rect 120644 27236 120645 27300
rect 120579 27235 120645 27236
rect 119234 20378 119266 20614
rect 119502 20378 119586 20614
rect 119822 20378 119854 20614
rect 119234 -5146 119854 20378
rect 121794 23294 122414 28000
rect 122606 26893 122666 29550
rect 123158 28930 123218 29550
rect 123709 29548 123710 29612
rect 123774 29548 123775 29612
rect 124800 29610 124860 30106
rect 125480 29885 125540 30106
rect 125477 29884 125543 29885
rect 125477 29820 125478 29884
rect 125542 29820 125543 29884
rect 125477 29819 125543 29820
rect 125888 29610 125948 30106
rect 127112 29610 127172 30106
rect 128064 29610 128124 30106
rect 128472 29610 128532 30106
rect 129560 29610 129620 30106
rect 130512 29613 130572 30106
rect 130509 29612 130575 29613
rect 124800 29550 124874 29610
rect 125888 29550 126346 29610
rect 127112 29550 127266 29610
rect 128064 29550 128186 29610
rect 128472 29550 128554 29610
rect 129560 29550 129658 29610
rect 123709 29547 123775 29548
rect 123158 28870 123770 28930
rect 122603 26892 122669 26893
rect 122603 26828 122604 26892
rect 122668 26828 122669 26892
rect 122603 26827 122669 26828
rect 121794 23058 121826 23294
rect 122062 23058 122146 23294
rect 122382 23058 122414 23294
rect 121794 3294 122414 23058
rect 121794 3058 121826 3294
rect 122062 3058 122146 3294
rect 122382 3058 122414 3294
rect 121794 -346 122414 3058
rect 121794 -582 121826 -346
rect 122062 -582 122146 -346
rect 122382 -582 122414 -346
rect 121794 -666 122414 -582
rect 121794 -902 121826 -666
rect 122062 -902 122146 -666
rect 122382 -902 122414 -666
rect 121794 -1894 122414 -902
rect 122954 24274 123574 28000
rect 123710 27165 123770 28870
rect 123707 27164 123773 27165
rect 123707 27100 123708 27164
rect 123772 27100 123773 27164
rect 123707 27099 123773 27100
rect 124814 27029 124874 29550
rect 124811 27028 124877 27029
rect 124811 26964 124812 27028
rect 124876 26964 124877 27028
rect 124811 26963 124877 26964
rect 122954 24038 122986 24274
rect 123222 24038 123306 24274
rect 123542 24038 123574 24274
rect 119234 -5382 119266 -5146
rect 119502 -5382 119586 -5146
rect 119822 -5382 119854 -5146
rect 119234 -5466 119854 -5382
rect 119234 -5702 119266 -5466
rect 119502 -5702 119586 -5466
rect 119822 -5702 119854 -5466
rect 119234 -5734 119854 -5702
rect 112954 -6342 112986 -6106
rect 113222 -6342 113306 -6106
rect 113542 -6342 113574 -6106
rect 112954 -6426 113574 -6342
rect 112954 -6662 112986 -6426
rect 113222 -6662 113306 -6426
rect 113542 -6662 113574 -6426
rect 112954 -7654 113574 -6662
rect 122954 -7066 123574 24038
rect 125514 26954 126134 28000
rect 126286 27573 126346 29550
rect 126283 27572 126349 27573
rect 126283 27508 126284 27572
rect 126348 27508 126349 27572
rect 126283 27507 126349 27508
rect 127206 27165 127266 29550
rect 128126 27573 128186 29550
rect 128494 28933 128554 29550
rect 128491 28932 128557 28933
rect 128491 28868 128492 28932
rect 128556 28868 128557 28932
rect 128491 28867 128557 28868
rect 129598 28253 129658 29550
rect 130509 29548 130510 29612
rect 130574 29548 130575 29612
rect 130648 29610 130708 30106
rect 132008 29610 132068 30106
rect 132960 29610 133020 30106
rect 133096 29610 133156 30106
rect 130648 29550 130762 29610
rect 130509 29547 130575 29548
rect 129595 28252 129661 28253
rect 129595 28188 129596 28252
rect 129660 28188 129661 28252
rect 129595 28187 129661 28188
rect 128123 27572 128189 27573
rect 128123 27508 128124 27572
rect 128188 27508 128189 27572
rect 128123 27507 128189 27508
rect 127203 27164 127269 27165
rect 127203 27100 127204 27164
rect 127268 27100 127269 27164
rect 127203 27099 127269 27100
rect 125514 26718 125546 26954
rect 125782 26718 125866 26954
rect 126102 26718 126134 26954
rect 125514 6954 126134 26718
rect 125514 6718 125546 6954
rect 125782 6718 125866 6954
rect 126102 6718 126134 6954
rect 125514 -2266 126134 6718
rect 125514 -2502 125546 -2266
rect 125782 -2502 125866 -2266
rect 126102 -2502 126134 -2266
rect 125514 -2586 126134 -2502
rect 125514 -2822 125546 -2586
rect 125782 -2822 125866 -2586
rect 126102 -2822 126134 -2586
rect 125514 -3814 126134 -2822
rect 129234 10614 129854 28000
rect 130702 26757 130762 29550
rect 131990 29550 132068 29610
rect 132726 29550 133020 29610
rect 133094 29550 133156 29610
rect 134184 29610 134244 30106
rect 135272 29610 135332 30106
rect 135816 29610 135876 30106
rect 136496 29610 136556 30106
rect 134184 29550 134258 29610
rect 135272 29550 135362 29610
rect 135816 29550 135914 29610
rect 131990 28253 132050 29550
rect 131987 28252 132053 28253
rect 131987 28188 131988 28252
rect 132052 28188 132053 28252
rect 131987 28187 132053 28188
rect 130699 26756 130765 26757
rect 130699 26692 130700 26756
rect 130764 26692 130765 26756
rect 130699 26691 130765 26692
rect 129234 10378 129266 10614
rect 129502 10378 129586 10614
rect 129822 10378 129854 10614
rect 129234 -4186 129854 10378
rect 131794 13294 132414 28000
rect 132726 27573 132786 29550
rect 133094 28797 133154 29550
rect 134198 28933 134258 29550
rect 134195 28932 134261 28933
rect 134195 28868 134196 28932
rect 134260 28868 134261 28932
rect 134195 28867 134261 28868
rect 133091 28796 133157 28797
rect 133091 28732 133092 28796
rect 133156 28732 133157 28796
rect 133091 28731 133157 28732
rect 135302 28661 135362 29550
rect 135854 28933 135914 29550
rect 136406 29550 136556 29610
rect 137856 29610 137916 30106
rect 138264 29610 138324 30106
rect 138944 29613 139004 30106
rect 137856 29550 137938 29610
rect 135851 28932 135917 28933
rect 135851 28868 135852 28932
rect 135916 28868 135917 28932
rect 135851 28867 135917 28868
rect 135299 28660 135365 28661
rect 135299 28596 135300 28660
rect 135364 28596 135365 28660
rect 135299 28595 135365 28596
rect 132723 27572 132789 27573
rect 132723 27508 132724 27572
rect 132788 27508 132789 27572
rect 132723 27507 132789 27508
rect 131794 13058 131826 13294
rect 132062 13058 132146 13294
rect 132382 13058 132414 13294
rect 131794 -1306 132414 13058
rect 131794 -1542 131826 -1306
rect 132062 -1542 132146 -1306
rect 132382 -1542 132414 -1306
rect 131794 -1626 132414 -1542
rect 131794 -1862 131826 -1626
rect 132062 -1862 132146 -1626
rect 132382 -1862 132414 -1626
rect 131794 -1894 132414 -1862
rect 132954 14274 133574 28000
rect 132954 14038 132986 14274
rect 133222 14038 133306 14274
rect 133542 14038 133574 14274
rect 129234 -4422 129266 -4186
rect 129502 -4422 129586 -4186
rect 129822 -4422 129854 -4186
rect 129234 -4506 129854 -4422
rect 129234 -4742 129266 -4506
rect 129502 -4742 129586 -4506
rect 129822 -4742 129854 -4506
rect 129234 -5734 129854 -4742
rect 122954 -7302 122986 -7066
rect 123222 -7302 123306 -7066
rect 123542 -7302 123574 -7066
rect 122954 -7386 123574 -7302
rect 122954 -7622 122986 -7386
rect 123222 -7622 123306 -7386
rect 123542 -7622 123574 -7386
rect 122954 -7654 123574 -7622
rect 132954 -6106 133574 14038
rect 135514 16954 136134 28000
rect 136406 27573 136466 29550
rect 137878 27573 137938 29550
rect 138246 29550 138324 29610
rect 138941 29612 139007 29613
rect 138246 28933 138306 29550
rect 138941 29548 138942 29612
rect 139006 29548 139007 29612
rect 140032 29610 140092 30106
rect 141120 29610 141180 30106
rect 142344 29610 142404 30106
rect 143432 29610 143492 30106
rect 140032 29550 140146 29610
rect 141120 29550 141250 29610
rect 142344 29550 142722 29610
rect 138941 29547 139007 29548
rect 138243 28932 138309 28933
rect 138243 28868 138244 28932
rect 138308 28868 138309 28932
rect 138243 28867 138309 28868
rect 136403 27572 136469 27573
rect 136403 27508 136404 27572
rect 136468 27508 136469 27572
rect 136403 27507 136469 27508
rect 137875 27572 137941 27573
rect 137875 27508 137876 27572
rect 137940 27508 137941 27572
rect 137875 27507 137941 27508
rect 135514 16718 135546 16954
rect 135782 16718 135866 16954
rect 136102 16718 136134 16954
rect 135514 -3226 136134 16718
rect 135514 -3462 135546 -3226
rect 135782 -3462 135866 -3226
rect 136102 -3462 136134 -3226
rect 135514 -3546 136134 -3462
rect 135514 -3782 135546 -3546
rect 135782 -3782 135866 -3546
rect 136102 -3782 136134 -3546
rect 135514 -3814 136134 -3782
rect 139234 20614 139854 28000
rect 140086 27573 140146 29550
rect 141190 27573 141250 29550
rect 140083 27572 140149 27573
rect 140083 27508 140084 27572
rect 140148 27508 140149 27572
rect 140083 27507 140149 27508
rect 141187 27572 141253 27573
rect 141187 27508 141188 27572
rect 141252 27508 141253 27572
rect 141187 27507 141253 27508
rect 139234 20378 139266 20614
rect 139502 20378 139586 20614
rect 139822 20378 139854 20614
rect 139234 -5146 139854 20378
rect 141794 23294 142414 28000
rect 142662 26621 142722 29550
rect 143398 29550 143492 29610
rect 144792 29610 144852 30106
rect 146016 29610 146076 30106
rect 146968 29610 147028 30106
rect 148328 29610 148388 30106
rect 149416 29610 149476 30106
rect 150504 29610 150564 30106
rect 144792 29550 147138 29610
rect 148328 29550 148426 29610
rect 149416 29550 150082 29610
rect 150504 29550 150634 29610
rect 143398 28253 143458 29550
rect 143395 28252 143461 28253
rect 143395 28188 143396 28252
rect 143460 28188 143461 28252
rect 143395 28187 143461 28188
rect 142659 26620 142725 26621
rect 142659 26556 142660 26620
rect 142724 26556 142725 26620
rect 142659 26555 142725 26556
rect 141794 23058 141826 23294
rect 142062 23058 142146 23294
rect 142382 23058 142414 23294
rect 141794 3294 142414 23058
rect 141794 3058 141826 3294
rect 142062 3058 142146 3294
rect 142382 3058 142414 3294
rect 141794 -346 142414 3058
rect 141794 -582 141826 -346
rect 142062 -582 142146 -346
rect 142382 -582 142414 -346
rect 141794 -666 142414 -582
rect 141794 -902 141826 -666
rect 142062 -902 142146 -666
rect 142382 -902 142414 -666
rect 141794 -1894 142414 -902
rect 142954 24274 143574 28000
rect 142954 24038 142986 24274
rect 143222 24038 143306 24274
rect 143542 24038 143574 24274
rect 139234 -5382 139266 -5146
rect 139502 -5382 139586 -5146
rect 139822 -5382 139854 -5146
rect 139234 -5466 139854 -5382
rect 139234 -5702 139266 -5466
rect 139502 -5702 139586 -5466
rect 139822 -5702 139854 -5466
rect 139234 -5734 139854 -5702
rect 132954 -6342 132986 -6106
rect 133222 -6342 133306 -6106
rect 133542 -6342 133574 -6106
rect 132954 -6426 133574 -6342
rect 132954 -6662 132986 -6426
rect 133222 -6662 133306 -6426
rect 133542 -6662 133574 -6426
rect 132954 -7654 133574 -6662
rect 142954 -7066 143574 24038
rect 145514 26954 146134 28000
rect 147078 27573 147138 29550
rect 148366 27573 148426 29550
rect 147075 27572 147141 27573
rect 147075 27508 147076 27572
rect 147140 27508 147141 27572
rect 147075 27507 147141 27508
rect 148363 27572 148429 27573
rect 148363 27508 148364 27572
rect 148428 27508 148429 27572
rect 148363 27507 148429 27508
rect 145514 26718 145546 26954
rect 145782 26718 145866 26954
rect 146102 26718 146134 26954
rect 145514 6954 146134 26718
rect 145514 6718 145546 6954
rect 145782 6718 145866 6954
rect 146102 6718 146134 6954
rect 145514 -2266 146134 6718
rect 145514 -2502 145546 -2266
rect 145782 -2502 145866 -2266
rect 146102 -2502 146134 -2266
rect 145514 -2586 146134 -2502
rect 145514 -2822 145546 -2586
rect 145782 -2822 145866 -2586
rect 146102 -2822 146134 -2586
rect 145514 -3814 146134 -2822
rect 149234 10614 149854 28000
rect 150022 27573 150082 29550
rect 150574 27573 150634 29550
rect 150019 27572 150085 27573
rect 150019 27508 150020 27572
rect 150084 27508 150085 27572
rect 150019 27507 150085 27508
rect 150571 27572 150637 27573
rect 150571 27508 150572 27572
rect 150636 27508 150637 27572
rect 150571 27507 150637 27508
rect 149234 10378 149266 10614
rect 149502 10378 149586 10614
rect 149822 10378 149854 10614
rect 149234 -4186 149854 10378
rect 151794 13294 152414 28000
rect 151794 13058 151826 13294
rect 152062 13058 152146 13294
rect 152382 13058 152414 13294
rect 151794 -1306 152414 13058
rect 151794 -1542 151826 -1306
rect 152062 -1542 152146 -1306
rect 152382 -1542 152414 -1306
rect 151794 -1626 152414 -1542
rect 151794 -1862 151826 -1626
rect 152062 -1862 152146 -1626
rect 152382 -1862 152414 -1626
rect 151794 -1894 152414 -1862
rect 152954 14274 153574 28000
rect 152954 14038 152986 14274
rect 153222 14038 153306 14274
rect 153542 14038 153574 14274
rect 149234 -4422 149266 -4186
rect 149502 -4422 149586 -4186
rect 149822 -4422 149854 -4186
rect 149234 -4506 149854 -4422
rect 149234 -4742 149266 -4506
rect 149502 -4742 149586 -4506
rect 149822 -4742 149854 -4506
rect 149234 -5734 149854 -4742
rect 142954 -7302 142986 -7066
rect 143222 -7302 143306 -7066
rect 143542 -7302 143574 -7066
rect 142954 -7386 143574 -7302
rect 142954 -7622 142986 -7386
rect 143222 -7622 143306 -7386
rect 143542 -7622 143574 -7386
rect 142954 -7654 143574 -7622
rect 152954 -6106 153574 14038
rect 155514 16954 156134 28000
rect 155514 16718 155546 16954
rect 155782 16718 155866 16954
rect 156102 16718 156134 16954
rect 155514 -3226 156134 16718
rect 155514 -3462 155546 -3226
rect 155782 -3462 155866 -3226
rect 156102 -3462 156134 -3226
rect 155514 -3546 156134 -3462
rect 155514 -3782 155546 -3546
rect 155782 -3782 155866 -3546
rect 156102 -3782 156134 -3546
rect 155514 -3814 156134 -3782
rect 159234 20614 159854 28000
rect 159234 20378 159266 20614
rect 159502 20378 159586 20614
rect 159822 20378 159854 20614
rect 159234 -5146 159854 20378
rect 161794 23294 162414 28000
rect 161794 23058 161826 23294
rect 162062 23058 162146 23294
rect 162382 23058 162414 23294
rect 161794 3294 162414 23058
rect 161794 3058 161826 3294
rect 162062 3058 162146 3294
rect 162382 3058 162414 3294
rect 161794 -346 162414 3058
rect 161794 -582 161826 -346
rect 162062 -582 162146 -346
rect 162382 -582 162414 -346
rect 161794 -666 162414 -582
rect 161794 -902 161826 -666
rect 162062 -902 162146 -666
rect 162382 -902 162414 -666
rect 161794 -1894 162414 -902
rect 162954 24274 163574 28000
rect 162954 24038 162986 24274
rect 163222 24038 163306 24274
rect 163542 24038 163574 24274
rect 159234 -5382 159266 -5146
rect 159502 -5382 159586 -5146
rect 159822 -5382 159854 -5146
rect 159234 -5466 159854 -5382
rect 159234 -5702 159266 -5466
rect 159502 -5702 159586 -5466
rect 159822 -5702 159854 -5466
rect 159234 -5734 159854 -5702
rect 152954 -6342 152986 -6106
rect 153222 -6342 153306 -6106
rect 153542 -6342 153574 -6106
rect 152954 -6426 153574 -6342
rect 152954 -6662 152986 -6426
rect 153222 -6662 153306 -6426
rect 153542 -6662 153574 -6426
rect 152954 -7654 153574 -6662
rect 162954 -7066 163574 24038
rect 165514 26954 166134 28000
rect 165514 26718 165546 26954
rect 165782 26718 165866 26954
rect 166102 26718 166134 26954
rect 165514 6954 166134 26718
rect 165514 6718 165546 6954
rect 165782 6718 165866 6954
rect 166102 6718 166134 6954
rect 165514 -2266 166134 6718
rect 165514 -2502 165546 -2266
rect 165782 -2502 165866 -2266
rect 166102 -2502 166134 -2266
rect 165514 -2586 166134 -2502
rect 165514 -2822 165546 -2586
rect 165782 -2822 165866 -2586
rect 166102 -2822 166134 -2586
rect 165514 -3814 166134 -2822
rect 169234 10614 169854 30378
rect 169234 10378 169266 10614
rect 169502 10378 169586 10614
rect 169822 10378 169854 10614
rect 169234 -4186 169854 10378
rect 171794 213294 172414 233058
rect 171794 213058 171826 213294
rect 172062 213058 172146 213294
rect 172382 213058 172414 213294
rect 171794 193294 172414 213058
rect 171794 193058 171826 193294
rect 172062 193058 172146 193294
rect 172382 193058 172414 193294
rect 171794 173294 172414 193058
rect 171794 173058 171826 173294
rect 172062 173058 172146 173294
rect 172382 173058 172414 173294
rect 171794 153294 172414 173058
rect 171794 153058 171826 153294
rect 172062 153058 172146 153294
rect 172382 153058 172414 153294
rect 171794 133294 172414 153058
rect 171794 133058 171826 133294
rect 172062 133058 172146 133294
rect 172382 133058 172414 133294
rect 171794 113294 172414 133058
rect 171794 113058 171826 113294
rect 172062 113058 172146 113294
rect 172382 113058 172414 113294
rect 171794 93294 172414 113058
rect 171794 93058 171826 93294
rect 172062 93058 172146 93294
rect 172382 93058 172414 93294
rect 171794 73294 172414 93058
rect 171794 73058 171826 73294
rect 172062 73058 172146 73294
rect 172382 73058 172414 73294
rect 171794 53294 172414 73058
rect 171794 53058 171826 53294
rect 172062 53058 172146 53294
rect 172382 53058 172414 53294
rect 171794 33294 172414 53058
rect 171794 33058 171826 33294
rect 172062 33058 172146 33294
rect 172382 33058 172414 33294
rect 171794 13294 172414 33058
rect 171794 13058 171826 13294
rect 172062 13058 172146 13294
rect 172382 13058 172414 13294
rect 171794 -1306 172414 13058
rect 171794 -1542 171826 -1306
rect 172062 -1542 172146 -1306
rect 172382 -1542 172414 -1306
rect 171794 -1626 172414 -1542
rect 171794 -1862 171826 -1626
rect 172062 -1862 172146 -1626
rect 172382 -1862 172414 -1626
rect 171794 -1894 172414 -1862
rect 172954 334274 173574 354038
rect 172954 334038 172986 334274
rect 173222 334038 173306 334274
rect 173542 334038 173574 334274
rect 172954 314274 173574 334038
rect 172954 314038 172986 314274
rect 173222 314038 173306 314274
rect 173542 314038 173574 314274
rect 172954 294274 173574 314038
rect 172954 294038 172986 294274
rect 173222 294038 173306 294274
rect 173542 294038 173574 294274
rect 172954 274274 173574 294038
rect 172954 274038 172986 274274
rect 173222 274038 173306 274274
rect 173542 274038 173574 274274
rect 172954 254274 173574 274038
rect 172954 254038 172986 254274
rect 173222 254038 173306 254274
rect 173542 254038 173574 254274
rect 172954 234274 173574 254038
rect 172954 234038 172986 234274
rect 173222 234038 173306 234274
rect 173542 234038 173574 234274
rect 172954 214274 173574 234038
rect 172954 214038 172986 214274
rect 173222 214038 173306 214274
rect 173542 214038 173574 214274
rect 172954 194274 173574 214038
rect 172954 194038 172986 194274
rect 173222 194038 173306 194274
rect 173542 194038 173574 194274
rect 172954 174274 173574 194038
rect 172954 174038 172986 174274
rect 173222 174038 173306 174274
rect 173542 174038 173574 174274
rect 172954 154274 173574 174038
rect 172954 154038 172986 154274
rect 173222 154038 173306 154274
rect 173542 154038 173574 154274
rect 172954 134274 173574 154038
rect 172954 134038 172986 134274
rect 173222 134038 173306 134274
rect 173542 134038 173574 134274
rect 172954 114274 173574 134038
rect 172954 114038 172986 114274
rect 173222 114038 173306 114274
rect 173542 114038 173574 114274
rect 172954 94274 173574 114038
rect 172954 94038 172986 94274
rect 173222 94038 173306 94274
rect 173542 94038 173574 94274
rect 172954 74274 173574 94038
rect 172954 74038 172986 74274
rect 173222 74038 173306 74274
rect 173542 74038 173574 74274
rect 172954 54274 173574 74038
rect 172954 54038 172986 54274
rect 173222 54038 173306 54274
rect 173542 54038 173574 54274
rect 172954 34274 173574 54038
rect 172954 34038 172986 34274
rect 173222 34038 173306 34274
rect 173542 34038 173574 34274
rect 172954 14274 173574 34038
rect 172954 14038 172986 14274
rect 173222 14038 173306 14274
rect 173542 14038 173574 14274
rect 169234 -4422 169266 -4186
rect 169502 -4422 169586 -4186
rect 169822 -4422 169854 -4186
rect 169234 -4506 169854 -4422
rect 169234 -4742 169266 -4506
rect 169502 -4742 169586 -4506
rect 169822 -4742 169854 -4506
rect 169234 -5734 169854 -4742
rect 162954 -7302 162986 -7066
rect 163222 -7302 163306 -7066
rect 163542 -7302 163574 -7066
rect 162954 -7386 163574 -7302
rect 162954 -7622 162986 -7386
rect 163222 -7622 163306 -7386
rect 163542 -7622 163574 -7386
rect 162954 -7654 163574 -7622
rect 172954 -6106 173574 14038
rect 174494 5677 174554 419595
rect 174678 340101 174738 420955
rect 175514 416954 176134 436718
rect 175514 416718 175546 416954
rect 175782 416718 175866 416954
rect 176102 416718 176134 416954
rect 175514 396954 176134 416718
rect 175514 396718 175546 396954
rect 175782 396718 175866 396954
rect 176102 396718 176134 396954
rect 175514 376954 176134 396718
rect 175514 376718 175546 376954
rect 175782 376718 175866 376954
rect 176102 376718 176134 376954
rect 175514 356954 176134 376718
rect 175514 356718 175546 356954
rect 175782 356718 175866 356954
rect 176102 356718 176134 356954
rect 174675 340100 174741 340101
rect 174675 340036 174676 340100
rect 174740 340036 174741 340100
rect 174675 340035 174741 340036
rect 175514 336954 176134 356718
rect 175514 336718 175546 336954
rect 175782 336718 175866 336954
rect 176102 336718 176134 336954
rect 175514 316954 176134 336718
rect 175514 316718 175546 316954
rect 175782 316718 175866 316954
rect 176102 316718 176134 316954
rect 175514 296954 176134 316718
rect 175514 296718 175546 296954
rect 175782 296718 175866 296954
rect 176102 296718 176134 296954
rect 175514 276954 176134 296718
rect 175514 276718 175546 276954
rect 175782 276718 175866 276954
rect 176102 276718 176134 276954
rect 175514 256954 176134 276718
rect 175514 256718 175546 256954
rect 175782 256718 175866 256954
rect 176102 256718 176134 256954
rect 175514 236954 176134 256718
rect 175514 236718 175546 236954
rect 175782 236718 175866 236954
rect 176102 236718 176134 236954
rect 175514 216954 176134 236718
rect 175514 216718 175546 216954
rect 175782 216718 175866 216954
rect 176102 216718 176134 216954
rect 175514 196954 176134 216718
rect 175514 196718 175546 196954
rect 175782 196718 175866 196954
rect 176102 196718 176134 196954
rect 175514 176954 176134 196718
rect 175514 176718 175546 176954
rect 175782 176718 175866 176954
rect 176102 176718 176134 176954
rect 175514 156954 176134 176718
rect 175514 156718 175546 156954
rect 175782 156718 175866 156954
rect 176102 156718 176134 156954
rect 175514 136954 176134 156718
rect 175514 136718 175546 136954
rect 175782 136718 175866 136954
rect 176102 136718 176134 136954
rect 175514 116954 176134 136718
rect 175514 116718 175546 116954
rect 175782 116718 175866 116954
rect 176102 116718 176134 116954
rect 175514 96954 176134 116718
rect 175514 96718 175546 96954
rect 175782 96718 175866 96954
rect 176102 96718 176134 96954
rect 175514 76954 176134 96718
rect 175514 76718 175546 76954
rect 175782 76718 175866 76954
rect 176102 76718 176134 76954
rect 175514 56954 176134 76718
rect 175514 56718 175546 56954
rect 175782 56718 175866 56954
rect 176102 56718 176134 56954
rect 175514 36954 176134 56718
rect 175514 36718 175546 36954
rect 175782 36718 175866 36954
rect 176102 36718 176134 36954
rect 175514 16954 176134 36718
rect 175514 16718 175546 16954
rect 175782 16718 175866 16954
rect 176102 16718 176134 16954
rect 174491 5676 174557 5677
rect 174491 5612 174492 5676
rect 174556 5612 174557 5676
rect 174491 5611 174557 5612
rect 175514 -3226 176134 16718
rect 175514 -3462 175546 -3226
rect 175782 -3462 175866 -3226
rect 176102 -3462 176134 -3226
rect 175514 -3546 176134 -3462
rect 175514 -3782 175546 -3546
rect 175782 -3782 175866 -3546
rect 176102 -3782 176134 -3546
rect 175514 -3814 176134 -3782
rect 179234 700614 179854 709082
rect 179234 700378 179266 700614
rect 179502 700378 179586 700614
rect 179822 700378 179854 700614
rect 179234 680614 179854 700378
rect 179234 680378 179266 680614
rect 179502 680378 179586 680614
rect 179822 680378 179854 680614
rect 179234 660614 179854 680378
rect 179234 660378 179266 660614
rect 179502 660378 179586 660614
rect 179822 660378 179854 660614
rect 179234 640614 179854 660378
rect 179234 640378 179266 640614
rect 179502 640378 179586 640614
rect 179822 640378 179854 640614
rect 179234 620614 179854 640378
rect 179234 620378 179266 620614
rect 179502 620378 179586 620614
rect 179822 620378 179854 620614
rect 179234 600614 179854 620378
rect 179234 600378 179266 600614
rect 179502 600378 179586 600614
rect 179822 600378 179854 600614
rect 179234 580614 179854 600378
rect 179234 580378 179266 580614
rect 179502 580378 179586 580614
rect 179822 580378 179854 580614
rect 179234 560614 179854 580378
rect 179234 560378 179266 560614
rect 179502 560378 179586 560614
rect 179822 560378 179854 560614
rect 179234 540614 179854 560378
rect 179234 540378 179266 540614
rect 179502 540378 179586 540614
rect 179822 540378 179854 540614
rect 179234 520614 179854 540378
rect 179234 520378 179266 520614
rect 179502 520378 179586 520614
rect 179822 520378 179854 520614
rect 179234 500614 179854 520378
rect 179234 500378 179266 500614
rect 179502 500378 179586 500614
rect 179822 500378 179854 500614
rect 179234 480614 179854 500378
rect 179234 480378 179266 480614
rect 179502 480378 179586 480614
rect 179822 480378 179854 480614
rect 179234 460614 179854 480378
rect 179234 460378 179266 460614
rect 179502 460378 179586 460614
rect 179822 460378 179854 460614
rect 179234 440614 179854 460378
rect 179234 440378 179266 440614
rect 179502 440378 179586 440614
rect 179822 440378 179854 440614
rect 179234 420614 179854 440378
rect 179234 420378 179266 420614
rect 179502 420378 179586 420614
rect 179822 420378 179854 420614
rect 179234 400614 179854 420378
rect 179234 400378 179266 400614
rect 179502 400378 179586 400614
rect 179822 400378 179854 400614
rect 179234 380614 179854 400378
rect 179234 380378 179266 380614
rect 179502 380378 179586 380614
rect 179822 380378 179854 380614
rect 179234 360614 179854 380378
rect 179234 360378 179266 360614
rect 179502 360378 179586 360614
rect 179822 360378 179854 360614
rect 179234 340614 179854 360378
rect 179234 340378 179266 340614
rect 179502 340378 179586 340614
rect 179822 340378 179854 340614
rect 179234 320614 179854 340378
rect 179234 320378 179266 320614
rect 179502 320378 179586 320614
rect 179822 320378 179854 320614
rect 179234 300614 179854 320378
rect 179234 300378 179266 300614
rect 179502 300378 179586 300614
rect 179822 300378 179854 300614
rect 179234 280614 179854 300378
rect 179234 280378 179266 280614
rect 179502 280378 179586 280614
rect 179822 280378 179854 280614
rect 179234 260614 179854 280378
rect 179234 260378 179266 260614
rect 179502 260378 179586 260614
rect 179822 260378 179854 260614
rect 179234 240614 179854 260378
rect 179234 240378 179266 240614
rect 179502 240378 179586 240614
rect 179822 240378 179854 240614
rect 179234 220614 179854 240378
rect 179234 220378 179266 220614
rect 179502 220378 179586 220614
rect 179822 220378 179854 220614
rect 179234 200614 179854 220378
rect 179234 200378 179266 200614
rect 179502 200378 179586 200614
rect 179822 200378 179854 200614
rect 179234 180614 179854 200378
rect 179234 180378 179266 180614
rect 179502 180378 179586 180614
rect 179822 180378 179854 180614
rect 179234 160614 179854 180378
rect 179234 160378 179266 160614
rect 179502 160378 179586 160614
rect 179822 160378 179854 160614
rect 179234 140614 179854 160378
rect 179234 140378 179266 140614
rect 179502 140378 179586 140614
rect 179822 140378 179854 140614
rect 179234 120614 179854 140378
rect 179234 120378 179266 120614
rect 179502 120378 179586 120614
rect 179822 120378 179854 120614
rect 179234 100614 179854 120378
rect 179234 100378 179266 100614
rect 179502 100378 179586 100614
rect 179822 100378 179854 100614
rect 179234 80614 179854 100378
rect 179234 80378 179266 80614
rect 179502 80378 179586 80614
rect 179822 80378 179854 80614
rect 179234 60614 179854 80378
rect 179234 60378 179266 60614
rect 179502 60378 179586 60614
rect 179822 60378 179854 60614
rect 179234 40614 179854 60378
rect 179234 40378 179266 40614
rect 179502 40378 179586 40614
rect 179822 40378 179854 40614
rect 179234 20614 179854 40378
rect 179234 20378 179266 20614
rect 179502 20378 179586 20614
rect 179822 20378 179854 20614
rect 179234 -5146 179854 20378
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 683294 182414 704282
rect 181794 683058 181826 683294
rect 182062 683058 182146 683294
rect 182382 683058 182414 683294
rect 181794 663294 182414 683058
rect 181794 663058 181826 663294
rect 182062 663058 182146 663294
rect 182382 663058 182414 663294
rect 181794 643294 182414 663058
rect 181794 643058 181826 643294
rect 182062 643058 182146 643294
rect 182382 643058 182414 643294
rect 181794 623294 182414 643058
rect 181794 623058 181826 623294
rect 182062 623058 182146 623294
rect 182382 623058 182414 623294
rect 181794 603294 182414 623058
rect 181794 603058 181826 603294
rect 182062 603058 182146 603294
rect 182382 603058 182414 603294
rect 181794 583294 182414 603058
rect 181794 583058 181826 583294
rect 182062 583058 182146 583294
rect 182382 583058 182414 583294
rect 181794 563294 182414 583058
rect 181794 563058 181826 563294
rect 182062 563058 182146 563294
rect 182382 563058 182414 563294
rect 181794 543294 182414 563058
rect 181794 543058 181826 543294
rect 182062 543058 182146 543294
rect 182382 543058 182414 543294
rect 181794 523294 182414 543058
rect 181794 523058 181826 523294
rect 182062 523058 182146 523294
rect 182382 523058 182414 523294
rect 181794 503294 182414 523058
rect 181794 503058 181826 503294
rect 182062 503058 182146 503294
rect 182382 503058 182414 503294
rect 181794 483294 182414 503058
rect 181794 483058 181826 483294
rect 182062 483058 182146 483294
rect 182382 483058 182414 483294
rect 181794 463294 182414 483058
rect 181794 463058 181826 463294
rect 182062 463058 182146 463294
rect 182382 463058 182414 463294
rect 181794 443294 182414 463058
rect 181794 443058 181826 443294
rect 182062 443058 182146 443294
rect 182382 443058 182414 443294
rect 181794 423294 182414 443058
rect 181794 423058 181826 423294
rect 182062 423058 182146 423294
rect 182382 423058 182414 423294
rect 181794 403294 182414 423058
rect 181794 403058 181826 403294
rect 182062 403058 182146 403294
rect 182382 403058 182414 403294
rect 181794 383294 182414 403058
rect 181794 383058 181826 383294
rect 182062 383058 182146 383294
rect 182382 383058 182414 383294
rect 181794 363294 182414 383058
rect 181794 363058 181826 363294
rect 182062 363058 182146 363294
rect 182382 363058 182414 363294
rect 181794 343294 182414 363058
rect 181794 343058 181826 343294
rect 182062 343058 182146 343294
rect 182382 343058 182414 343294
rect 181794 323294 182414 343058
rect 181794 323058 181826 323294
rect 182062 323058 182146 323294
rect 182382 323058 182414 323294
rect 181794 303294 182414 323058
rect 181794 303058 181826 303294
rect 182062 303058 182146 303294
rect 182382 303058 182414 303294
rect 181794 283294 182414 303058
rect 181794 283058 181826 283294
rect 182062 283058 182146 283294
rect 182382 283058 182414 283294
rect 181794 263294 182414 283058
rect 181794 263058 181826 263294
rect 182062 263058 182146 263294
rect 182382 263058 182414 263294
rect 181794 243294 182414 263058
rect 181794 243058 181826 243294
rect 182062 243058 182146 243294
rect 182382 243058 182414 243294
rect 181794 223294 182414 243058
rect 181794 223058 181826 223294
rect 182062 223058 182146 223294
rect 182382 223058 182414 223294
rect 181794 203294 182414 223058
rect 181794 203058 181826 203294
rect 182062 203058 182146 203294
rect 182382 203058 182414 203294
rect 181794 183294 182414 203058
rect 181794 183058 181826 183294
rect 182062 183058 182146 183294
rect 182382 183058 182414 183294
rect 181794 163294 182414 183058
rect 181794 163058 181826 163294
rect 182062 163058 182146 163294
rect 182382 163058 182414 163294
rect 181794 143294 182414 163058
rect 181794 143058 181826 143294
rect 182062 143058 182146 143294
rect 182382 143058 182414 143294
rect 181794 123294 182414 143058
rect 181794 123058 181826 123294
rect 182062 123058 182146 123294
rect 182382 123058 182414 123294
rect 181794 103294 182414 123058
rect 181794 103058 181826 103294
rect 182062 103058 182146 103294
rect 182382 103058 182414 103294
rect 181794 83294 182414 103058
rect 181794 83058 181826 83294
rect 182062 83058 182146 83294
rect 182382 83058 182414 83294
rect 181794 63294 182414 83058
rect 181794 63058 181826 63294
rect 182062 63058 182146 63294
rect 182382 63058 182414 63294
rect 181794 43294 182414 63058
rect 181794 43058 181826 43294
rect 182062 43058 182146 43294
rect 182382 43058 182414 43294
rect 181794 23294 182414 43058
rect 181794 23058 181826 23294
rect 182062 23058 182146 23294
rect 182382 23058 182414 23294
rect 181794 3294 182414 23058
rect 181794 3058 181826 3294
rect 182062 3058 182146 3294
rect 182382 3058 182414 3294
rect 181794 -346 182414 3058
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 182954 684274 183574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 182954 684038 182986 684274
rect 183222 684038 183306 684274
rect 183542 684038 183574 684274
rect 182954 664274 183574 684038
rect 182954 664038 182986 664274
rect 183222 664038 183306 664274
rect 183542 664038 183574 664274
rect 182954 644274 183574 664038
rect 182954 644038 182986 644274
rect 183222 644038 183306 644274
rect 183542 644038 183574 644274
rect 182954 624274 183574 644038
rect 182954 624038 182986 624274
rect 183222 624038 183306 624274
rect 183542 624038 183574 624274
rect 182954 604274 183574 624038
rect 182954 604038 182986 604274
rect 183222 604038 183306 604274
rect 183542 604038 183574 604274
rect 182954 584274 183574 604038
rect 182954 584038 182986 584274
rect 183222 584038 183306 584274
rect 183542 584038 183574 584274
rect 182954 564274 183574 584038
rect 182954 564038 182986 564274
rect 183222 564038 183306 564274
rect 183542 564038 183574 564274
rect 182954 544274 183574 564038
rect 182954 544038 182986 544274
rect 183222 544038 183306 544274
rect 183542 544038 183574 544274
rect 182954 524274 183574 544038
rect 182954 524038 182986 524274
rect 183222 524038 183306 524274
rect 183542 524038 183574 524274
rect 182954 504274 183574 524038
rect 182954 504038 182986 504274
rect 183222 504038 183306 504274
rect 183542 504038 183574 504274
rect 182954 484274 183574 504038
rect 182954 484038 182986 484274
rect 183222 484038 183306 484274
rect 183542 484038 183574 484274
rect 182954 464274 183574 484038
rect 182954 464038 182986 464274
rect 183222 464038 183306 464274
rect 183542 464038 183574 464274
rect 182954 444274 183574 464038
rect 182954 444038 182986 444274
rect 183222 444038 183306 444274
rect 183542 444038 183574 444274
rect 182954 424274 183574 444038
rect 182954 424038 182986 424274
rect 183222 424038 183306 424274
rect 183542 424038 183574 424274
rect 182954 404274 183574 424038
rect 182954 404038 182986 404274
rect 183222 404038 183306 404274
rect 183542 404038 183574 404274
rect 182954 384274 183574 404038
rect 182954 384038 182986 384274
rect 183222 384038 183306 384274
rect 183542 384038 183574 384274
rect 182954 364274 183574 384038
rect 182954 364038 182986 364274
rect 183222 364038 183306 364274
rect 183542 364038 183574 364274
rect 182954 344274 183574 364038
rect 182954 344038 182986 344274
rect 183222 344038 183306 344274
rect 183542 344038 183574 344274
rect 182954 324274 183574 344038
rect 182954 324038 182986 324274
rect 183222 324038 183306 324274
rect 183542 324038 183574 324274
rect 182954 304274 183574 324038
rect 182954 304038 182986 304274
rect 183222 304038 183306 304274
rect 183542 304038 183574 304274
rect 182954 284274 183574 304038
rect 182954 284038 182986 284274
rect 183222 284038 183306 284274
rect 183542 284038 183574 284274
rect 182954 264274 183574 284038
rect 182954 264038 182986 264274
rect 183222 264038 183306 264274
rect 183542 264038 183574 264274
rect 182954 244274 183574 264038
rect 182954 244038 182986 244274
rect 183222 244038 183306 244274
rect 183542 244038 183574 244274
rect 182954 224274 183574 244038
rect 182954 224038 182986 224274
rect 183222 224038 183306 224274
rect 183542 224038 183574 224274
rect 182954 204274 183574 224038
rect 182954 204038 182986 204274
rect 183222 204038 183306 204274
rect 183542 204038 183574 204274
rect 182954 184274 183574 204038
rect 182954 184038 182986 184274
rect 183222 184038 183306 184274
rect 183542 184038 183574 184274
rect 182954 164274 183574 184038
rect 182954 164038 182986 164274
rect 183222 164038 183306 164274
rect 183542 164038 183574 164274
rect 182954 144274 183574 164038
rect 182954 144038 182986 144274
rect 183222 144038 183306 144274
rect 183542 144038 183574 144274
rect 182954 124274 183574 144038
rect 182954 124038 182986 124274
rect 183222 124038 183306 124274
rect 183542 124038 183574 124274
rect 182954 104274 183574 124038
rect 182954 104038 182986 104274
rect 183222 104038 183306 104274
rect 183542 104038 183574 104274
rect 182954 84274 183574 104038
rect 182954 84038 182986 84274
rect 183222 84038 183306 84274
rect 183542 84038 183574 84274
rect 182954 64274 183574 84038
rect 182954 64038 182986 64274
rect 183222 64038 183306 64274
rect 183542 64038 183574 64274
rect 182954 44274 183574 64038
rect 182954 44038 182986 44274
rect 183222 44038 183306 44274
rect 183542 44038 183574 44274
rect 182954 24274 183574 44038
rect 182954 24038 182986 24274
rect 183222 24038 183306 24274
rect 183542 24038 183574 24274
rect 179234 -5382 179266 -5146
rect 179502 -5382 179586 -5146
rect 179822 -5382 179854 -5146
rect 179234 -5466 179854 -5382
rect 179234 -5702 179266 -5466
rect 179502 -5702 179586 -5466
rect 179822 -5702 179854 -5466
rect 179234 -5734 179854 -5702
rect 172954 -6342 172986 -6106
rect 173222 -6342 173306 -6106
rect 173542 -6342 173574 -6106
rect 172954 -6426 173574 -6342
rect 172954 -6662 172986 -6426
rect 173222 -6662 173306 -6426
rect 173542 -6662 173574 -6426
rect 172954 -7654 173574 -6662
rect 182954 -7066 183574 24038
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 185514 686954 186134 706202
rect 185514 686718 185546 686954
rect 185782 686718 185866 686954
rect 186102 686718 186134 686954
rect 185514 666954 186134 686718
rect 185514 666718 185546 666954
rect 185782 666718 185866 666954
rect 186102 666718 186134 666954
rect 185514 646954 186134 666718
rect 185514 646718 185546 646954
rect 185782 646718 185866 646954
rect 186102 646718 186134 646954
rect 185514 626954 186134 646718
rect 185514 626718 185546 626954
rect 185782 626718 185866 626954
rect 186102 626718 186134 626954
rect 185514 606954 186134 626718
rect 185514 606718 185546 606954
rect 185782 606718 185866 606954
rect 186102 606718 186134 606954
rect 185514 586954 186134 606718
rect 185514 586718 185546 586954
rect 185782 586718 185866 586954
rect 186102 586718 186134 586954
rect 185514 566954 186134 586718
rect 185514 566718 185546 566954
rect 185782 566718 185866 566954
rect 186102 566718 186134 566954
rect 185514 546954 186134 566718
rect 185514 546718 185546 546954
rect 185782 546718 185866 546954
rect 186102 546718 186134 546954
rect 185514 526954 186134 546718
rect 185514 526718 185546 526954
rect 185782 526718 185866 526954
rect 186102 526718 186134 526954
rect 185514 506954 186134 526718
rect 185514 506718 185546 506954
rect 185782 506718 185866 506954
rect 186102 506718 186134 506954
rect 185514 486954 186134 506718
rect 185514 486718 185546 486954
rect 185782 486718 185866 486954
rect 186102 486718 186134 486954
rect 185514 466954 186134 486718
rect 185514 466718 185546 466954
rect 185782 466718 185866 466954
rect 186102 466718 186134 466954
rect 185514 446954 186134 466718
rect 185514 446718 185546 446954
rect 185782 446718 185866 446954
rect 186102 446718 186134 446954
rect 185514 426954 186134 446718
rect 185514 426718 185546 426954
rect 185782 426718 185866 426954
rect 186102 426718 186134 426954
rect 185514 406954 186134 426718
rect 185514 406718 185546 406954
rect 185782 406718 185866 406954
rect 186102 406718 186134 406954
rect 185514 386954 186134 406718
rect 185514 386718 185546 386954
rect 185782 386718 185866 386954
rect 186102 386718 186134 386954
rect 185514 366954 186134 386718
rect 185514 366718 185546 366954
rect 185782 366718 185866 366954
rect 186102 366718 186134 366954
rect 185514 346954 186134 366718
rect 185514 346718 185546 346954
rect 185782 346718 185866 346954
rect 186102 346718 186134 346954
rect 185514 326954 186134 346718
rect 185514 326718 185546 326954
rect 185782 326718 185866 326954
rect 186102 326718 186134 326954
rect 185514 306954 186134 326718
rect 185514 306718 185546 306954
rect 185782 306718 185866 306954
rect 186102 306718 186134 306954
rect 185514 286954 186134 306718
rect 185514 286718 185546 286954
rect 185782 286718 185866 286954
rect 186102 286718 186134 286954
rect 185514 266954 186134 286718
rect 185514 266718 185546 266954
rect 185782 266718 185866 266954
rect 186102 266718 186134 266954
rect 185514 246954 186134 266718
rect 185514 246718 185546 246954
rect 185782 246718 185866 246954
rect 186102 246718 186134 246954
rect 185514 226954 186134 246718
rect 185514 226718 185546 226954
rect 185782 226718 185866 226954
rect 186102 226718 186134 226954
rect 185514 206954 186134 226718
rect 185514 206718 185546 206954
rect 185782 206718 185866 206954
rect 186102 206718 186134 206954
rect 185514 186954 186134 206718
rect 185514 186718 185546 186954
rect 185782 186718 185866 186954
rect 186102 186718 186134 186954
rect 185514 166954 186134 186718
rect 185514 166718 185546 166954
rect 185782 166718 185866 166954
rect 186102 166718 186134 166954
rect 185514 146954 186134 166718
rect 185514 146718 185546 146954
rect 185782 146718 185866 146954
rect 186102 146718 186134 146954
rect 185514 126954 186134 146718
rect 185514 126718 185546 126954
rect 185782 126718 185866 126954
rect 186102 126718 186134 126954
rect 185514 106954 186134 126718
rect 185514 106718 185546 106954
rect 185782 106718 185866 106954
rect 186102 106718 186134 106954
rect 185514 86954 186134 106718
rect 185514 86718 185546 86954
rect 185782 86718 185866 86954
rect 186102 86718 186134 86954
rect 185514 66954 186134 86718
rect 185514 66718 185546 66954
rect 185782 66718 185866 66954
rect 186102 66718 186134 66954
rect 185514 46954 186134 66718
rect 185514 46718 185546 46954
rect 185782 46718 185866 46954
rect 186102 46718 186134 46954
rect 185514 26954 186134 46718
rect 185514 26718 185546 26954
rect 185782 26718 185866 26954
rect 186102 26718 186134 26954
rect 185514 6954 186134 26718
rect 185514 6718 185546 6954
rect 185782 6718 185866 6954
rect 186102 6718 186134 6954
rect 185514 -2266 186134 6718
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 690614 189854 708122
rect 189234 690378 189266 690614
rect 189502 690378 189586 690614
rect 189822 690378 189854 690614
rect 189234 670614 189854 690378
rect 189234 670378 189266 670614
rect 189502 670378 189586 670614
rect 189822 670378 189854 670614
rect 189234 650614 189854 670378
rect 189234 650378 189266 650614
rect 189502 650378 189586 650614
rect 189822 650378 189854 650614
rect 189234 630614 189854 650378
rect 189234 630378 189266 630614
rect 189502 630378 189586 630614
rect 189822 630378 189854 630614
rect 189234 610614 189854 630378
rect 189234 610378 189266 610614
rect 189502 610378 189586 610614
rect 189822 610378 189854 610614
rect 189234 590614 189854 610378
rect 189234 590378 189266 590614
rect 189502 590378 189586 590614
rect 189822 590378 189854 590614
rect 189234 570614 189854 590378
rect 189234 570378 189266 570614
rect 189502 570378 189586 570614
rect 189822 570378 189854 570614
rect 189234 550614 189854 570378
rect 189234 550378 189266 550614
rect 189502 550378 189586 550614
rect 189822 550378 189854 550614
rect 189234 530614 189854 550378
rect 189234 530378 189266 530614
rect 189502 530378 189586 530614
rect 189822 530378 189854 530614
rect 189234 510614 189854 530378
rect 189234 510378 189266 510614
rect 189502 510378 189586 510614
rect 189822 510378 189854 510614
rect 189234 490614 189854 510378
rect 189234 490378 189266 490614
rect 189502 490378 189586 490614
rect 189822 490378 189854 490614
rect 189234 470614 189854 490378
rect 189234 470378 189266 470614
rect 189502 470378 189586 470614
rect 189822 470378 189854 470614
rect 189234 450614 189854 470378
rect 189234 450378 189266 450614
rect 189502 450378 189586 450614
rect 189822 450378 189854 450614
rect 189234 430614 189854 450378
rect 189234 430378 189266 430614
rect 189502 430378 189586 430614
rect 189822 430378 189854 430614
rect 189234 410614 189854 430378
rect 189234 410378 189266 410614
rect 189502 410378 189586 410614
rect 189822 410378 189854 410614
rect 189234 390614 189854 410378
rect 189234 390378 189266 390614
rect 189502 390378 189586 390614
rect 189822 390378 189854 390614
rect 189234 370614 189854 390378
rect 189234 370378 189266 370614
rect 189502 370378 189586 370614
rect 189822 370378 189854 370614
rect 189234 350614 189854 370378
rect 189234 350378 189266 350614
rect 189502 350378 189586 350614
rect 189822 350378 189854 350614
rect 189234 330614 189854 350378
rect 189234 330378 189266 330614
rect 189502 330378 189586 330614
rect 189822 330378 189854 330614
rect 189234 310614 189854 330378
rect 189234 310378 189266 310614
rect 189502 310378 189586 310614
rect 189822 310378 189854 310614
rect 189234 290614 189854 310378
rect 189234 290378 189266 290614
rect 189502 290378 189586 290614
rect 189822 290378 189854 290614
rect 189234 270614 189854 290378
rect 189234 270378 189266 270614
rect 189502 270378 189586 270614
rect 189822 270378 189854 270614
rect 189234 250614 189854 270378
rect 189234 250378 189266 250614
rect 189502 250378 189586 250614
rect 189822 250378 189854 250614
rect 189234 230614 189854 250378
rect 189234 230378 189266 230614
rect 189502 230378 189586 230614
rect 189822 230378 189854 230614
rect 189234 210614 189854 230378
rect 189234 210378 189266 210614
rect 189502 210378 189586 210614
rect 189822 210378 189854 210614
rect 189234 190614 189854 210378
rect 189234 190378 189266 190614
rect 189502 190378 189586 190614
rect 189822 190378 189854 190614
rect 189234 170614 189854 190378
rect 189234 170378 189266 170614
rect 189502 170378 189586 170614
rect 189822 170378 189854 170614
rect 189234 150614 189854 170378
rect 189234 150378 189266 150614
rect 189502 150378 189586 150614
rect 189822 150378 189854 150614
rect 189234 130614 189854 150378
rect 189234 130378 189266 130614
rect 189502 130378 189586 130614
rect 189822 130378 189854 130614
rect 189234 110614 189854 130378
rect 189234 110378 189266 110614
rect 189502 110378 189586 110614
rect 189822 110378 189854 110614
rect 189234 90614 189854 110378
rect 189234 90378 189266 90614
rect 189502 90378 189586 90614
rect 189822 90378 189854 90614
rect 189234 70614 189854 90378
rect 189234 70378 189266 70614
rect 189502 70378 189586 70614
rect 189822 70378 189854 70614
rect 189234 50614 189854 70378
rect 189234 50378 189266 50614
rect 189502 50378 189586 50614
rect 189822 50378 189854 50614
rect 189234 30614 189854 50378
rect 189234 30378 189266 30614
rect 189502 30378 189586 30614
rect 189822 30378 189854 30614
rect 189234 10614 189854 30378
rect 189234 10378 189266 10614
rect 189502 10378 189586 10614
rect 189822 10378 189854 10614
rect 189234 -4186 189854 10378
rect 191794 705798 192414 705830
rect 191794 705562 191826 705798
rect 192062 705562 192146 705798
rect 192382 705562 192414 705798
rect 191794 705478 192414 705562
rect 191794 705242 191826 705478
rect 192062 705242 192146 705478
rect 192382 705242 192414 705478
rect 191794 693294 192414 705242
rect 191794 693058 191826 693294
rect 192062 693058 192146 693294
rect 192382 693058 192414 693294
rect 191794 673294 192414 693058
rect 191794 673058 191826 673294
rect 192062 673058 192146 673294
rect 192382 673058 192414 673294
rect 191794 653294 192414 673058
rect 191794 653058 191826 653294
rect 192062 653058 192146 653294
rect 192382 653058 192414 653294
rect 191794 633294 192414 653058
rect 191794 633058 191826 633294
rect 192062 633058 192146 633294
rect 192382 633058 192414 633294
rect 191794 613294 192414 633058
rect 191794 613058 191826 613294
rect 192062 613058 192146 613294
rect 192382 613058 192414 613294
rect 191794 593294 192414 613058
rect 191794 593058 191826 593294
rect 192062 593058 192146 593294
rect 192382 593058 192414 593294
rect 191794 573294 192414 593058
rect 191794 573058 191826 573294
rect 192062 573058 192146 573294
rect 192382 573058 192414 573294
rect 191794 553294 192414 573058
rect 191794 553058 191826 553294
rect 192062 553058 192146 553294
rect 192382 553058 192414 553294
rect 191794 533294 192414 553058
rect 191794 533058 191826 533294
rect 192062 533058 192146 533294
rect 192382 533058 192414 533294
rect 191794 513294 192414 533058
rect 191794 513058 191826 513294
rect 192062 513058 192146 513294
rect 192382 513058 192414 513294
rect 191794 493294 192414 513058
rect 191794 493058 191826 493294
rect 192062 493058 192146 493294
rect 192382 493058 192414 493294
rect 191794 473294 192414 493058
rect 191794 473058 191826 473294
rect 192062 473058 192146 473294
rect 192382 473058 192414 473294
rect 191794 453294 192414 473058
rect 191794 453058 191826 453294
rect 192062 453058 192146 453294
rect 192382 453058 192414 453294
rect 191794 433294 192414 453058
rect 191794 433058 191826 433294
rect 192062 433058 192146 433294
rect 192382 433058 192414 433294
rect 191794 413294 192414 433058
rect 191794 413058 191826 413294
rect 192062 413058 192146 413294
rect 192382 413058 192414 413294
rect 191794 393294 192414 413058
rect 191794 393058 191826 393294
rect 192062 393058 192146 393294
rect 192382 393058 192414 393294
rect 191794 373294 192414 393058
rect 191794 373058 191826 373294
rect 192062 373058 192146 373294
rect 192382 373058 192414 373294
rect 191794 353294 192414 373058
rect 191794 353058 191826 353294
rect 192062 353058 192146 353294
rect 192382 353058 192414 353294
rect 191794 333294 192414 353058
rect 191794 333058 191826 333294
rect 192062 333058 192146 333294
rect 192382 333058 192414 333294
rect 191794 313294 192414 333058
rect 191794 313058 191826 313294
rect 192062 313058 192146 313294
rect 192382 313058 192414 313294
rect 191794 293294 192414 313058
rect 191794 293058 191826 293294
rect 192062 293058 192146 293294
rect 192382 293058 192414 293294
rect 191794 273294 192414 293058
rect 191794 273058 191826 273294
rect 192062 273058 192146 273294
rect 192382 273058 192414 273294
rect 191794 253294 192414 273058
rect 191794 253058 191826 253294
rect 192062 253058 192146 253294
rect 192382 253058 192414 253294
rect 191794 233294 192414 253058
rect 191794 233058 191826 233294
rect 192062 233058 192146 233294
rect 192382 233058 192414 233294
rect 191794 213294 192414 233058
rect 191794 213058 191826 213294
rect 192062 213058 192146 213294
rect 192382 213058 192414 213294
rect 191794 193294 192414 213058
rect 191794 193058 191826 193294
rect 192062 193058 192146 193294
rect 192382 193058 192414 193294
rect 191794 173294 192414 193058
rect 191794 173058 191826 173294
rect 192062 173058 192146 173294
rect 192382 173058 192414 173294
rect 191794 153294 192414 173058
rect 191794 153058 191826 153294
rect 192062 153058 192146 153294
rect 192382 153058 192414 153294
rect 191794 133294 192414 153058
rect 191794 133058 191826 133294
rect 192062 133058 192146 133294
rect 192382 133058 192414 133294
rect 191794 113294 192414 133058
rect 191794 113058 191826 113294
rect 192062 113058 192146 113294
rect 192382 113058 192414 113294
rect 191794 93294 192414 113058
rect 191794 93058 191826 93294
rect 192062 93058 192146 93294
rect 192382 93058 192414 93294
rect 191794 73294 192414 93058
rect 191794 73058 191826 73294
rect 192062 73058 192146 73294
rect 192382 73058 192414 73294
rect 191794 53294 192414 73058
rect 191794 53058 191826 53294
rect 192062 53058 192146 53294
rect 192382 53058 192414 53294
rect 191794 33294 192414 53058
rect 191794 33058 191826 33294
rect 192062 33058 192146 33294
rect 192382 33058 192414 33294
rect 191794 13294 192414 33058
rect 191794 13058 191826 13294
rect 192062 13058 192146 13294
rect 192382 13058 192414 13294
rect 191794 -1306 192414 13058
rect 191794 -1542 191826 -1306
rect 192062 -1542 192146 -1306
rect 192382 -1542 192414 -1306
rect 191794 -1626 192414 -1542
rect 191794 -1862 191826 -1626
rect 192062 -1862 192146 -1626
rect 192382 -1862 192414 -1626
rect 191794 -1894 192414 -1862
rect 192954 694274 193574 710042
rect 202954 711558 203574 711590
rect 202954 711322 202986 711558
rect 203222 711322 203306 711558
rect 203542 711322 203574 711558
rect 202954 711238 203574 711322
rect 202954 711002 202986 711238
rect 203222 711002 203306 711238
rect 203542 711002 203574 711238
rect 199234 709638 199854 709670
rect 199234 709402 199266 709638
rect 199502 709402 199586 709638
rect 199822 709402 199854 709638
rect 199234 709318 199854 709402
rect 199234 709082 199266 709318
rect 199502 709082 199586 709318
rect 199822 709082 199854 709318
rect 192954 694038 192986 694274
rect 193222 694038 193306 694274
rect 193542 694038 193574 694274
rect 192954 674274 193574 694038
rect 192954 674038 192986 674274
rect 193222 674038 193306 674274
rect 193542 674038 193574 674274
rect 192954 654274 193574 674038
rect 192954 654038 192986 654274
rect 193222 654038 193306 654274
rect 193542 654038 193574 654274
rect 192954 634274 193574 654038
rect 192954 634038 192986 634274
rect 193222 634038 193306 634274
rect 193542 634038 193574 634274
rect 192954 614274 193574 634038
rect 192954 614038 192986 614274
rect 193222 614038 193306 614274
rect 193542 614038 193574 614274
rect 192954 594274 193574 614038
rect 192954 594038 192986 594274
rect 193222 594038 193306 594274
rect 193542 594038 193574 594274
rect 192954 574274 193574 594038
rect 192954 574038 192986 574274
rect 193222 574038 193306 574274
rect 193542 574038 193574 574274
rect 192954 554274 193574 574038
rect 192954 554038 192986 554274
rect 193222 554038 193306 554274
rect 193542 554038 193574 554274
rect 192954 534274 193574 554038
rect 192954 534038 192986 534274
rect 193222 534038 193306 534274
rect 193542 534038 193574 534274
rect 192954 514274 193574 534038
rect 192954 514038 192986 514274
rect 193222 514038 193306 514274
rect 193542 514038 193574 514274
rect 192954 494274 193574 514038
rect 192954 494038 192986 494274
rect 193222 494038 193306 494274
rect 193542 494038 193574 494274
rect 192954 474274 193574 494038
rect 192954 474038 192986 474274
rect 193222 474038 193306 474274
rect 193542 474038 193574 474274
rect 192954 454274 193574 474038
rect 192954 454038 192986 454274
rect 193222 454038 193306 454274
rect 193542 454038 193574 454274
rect 192954 434274 193574 454038
rect 192954 434038 192986 434274
rect 193222 434038 193306 434274
rect 193542 434038 193574 434274
rect 192954 414274 193574 434038
rect 192954 414038 192986 414274
rect 193222 414038 193306 414274
rect 193542 414038 193574 414274
rect 192954 394274 193574 414038
rect 192954 394038 192986 394274
rect 193222 394038 193306 394274
rect 193542 394038 193574 394274
rect 192954 374274 193574 394038
rect 192954 374038 192986 374274
rect 193222 374038 193306 374274
rect 193542 374038 193574 374274
rect 192954 354274 193574 374038
rect 192954 354038 192986 354274
rect 193222 354038 193306 354274
rect 193542 354038 193574 354274
rect 192954 334274 193574 354038
rect 192954 334038 192986 334274
rect 193222 334038 193306 334274
rect 193542 334038 193574 334274
rect 192954 314274 193574 334038
rect 192954 314038 192986 314274
rect 193222 314038 193306 314274
rect 193542 314038 193574 314274
rect 192954 294274 193574 314038
rect 192954 294038 192986 294274
rect 193222 294038 193306 294274
rect 193542 294038 193574 294274
rect 192954 274274 193574 294038
rect 192954 274038 192986 274274
rect 193222 274038 193306 274274
rect 193542 274038 193574 274274
rect 192954 254274 193574 274038
rect 192954 254038 192986 254274
rect 193222 254038 193306 254274
rect 193542 254038 193574 254274
rect 192954 234274 193574 254038
rect 192954 234038 192986 234274
rect 193222 234038 193306 234274
rect 193542 234038 193574 234274
rect 192954 214274 193574 234038
rect 192954 214038 192986 214274
rect 193222 214038 193306 214274
rect 193542 214038 193574 214274
rect 192954 194274 193574 214038
rect 192954 194038 192986 194274
rect 193222 194038 193306 194274
rect 193542 194038 193574 194274
rect 192954 174274 193574 194038
rect 192954 174038 192986 174274
rect 193222 174038 193306 174274
rect 193542 174038 193574 174274
rect 192954 154274 193574 174038
rect 192954 154038 192986 154274
rect 193222 154038 193306 154274
rect 193542 154038 193574 154274
rect 192954 134274 193574 154038
rect 192954 134038 192986 134274
rect 193222 134038 193306 134274
rect 193542 134038 193574 134274
rect 192954 114274 193574 134038
rect 192954 114038 192986 114274
rect 193222 114038 193306 114274
rect 193542 114038 193574 114274
rect 192954 94274 193574 114038
rect 192954 94038 192986 94274
rect 193222 94038 193306 94274
rect 193542 94038 193574 94274
rect 192954 74274 193574 94038
rect 192954 74038 192986 74274
rect 193222 74038 193306 74274
rect 193542 74038 193574 74274
rect 192954 54274 193574 74038
rect 192954 54038 192986 54274
rect 193222 54038 193306 54274
rect 193542 54038 193574 54274
rect 192954 34274 193574 54038
rect 192954 34038 192986 34274
rect 193222 34038 193306 34274
rect 193542 34038 193574 34274
rect 192954 14274 193574 34038
rect 192954 14038 192986 14274
rect 193222 14038 193306 14274
rect 193542 14038 193574 14274
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 182954 -7302 182986 -7066
rect 183222 -7302 183306 -7066
rect 183542 -7302 183574 -7066
rect 182954 -7386 183574 -7302
rect 182954 -7622 182986 -7386
rect 183222 -7622 183306 -7386
rect 183542 -7622 183574 -7386
rect 182954 -7654 183574 -7622
rect 192954 -6106 193574 14038
rect 195514 707718 196134 707750
rect 195514 707482 195546 707718
rect 195782 707482 195866 707718
rect 196102 707482 196134 707718
rect 195514 707398 196134 707482
rect 195514 707162 195546 707398
rect 195782 707162 195866 707398
rect 196102 707162 196134 707398
rect 195514 696954 196134 707162
rect 196571 700636 196637 700637
rect 196571 700572 196572 700636
rect 196636 700572 196637 700636
rect 196571 700571 196637 700572
rect 199234 700614 199854 709082
rect 195514 696718 195546 696954
rect 195782 696718 195866 696954
rect 196102 696718 196134 696954
rect 195514 676954 196134 696718
rect 195514 676718 195546 676954
rect 195782 676718 195866 676954
rect 196102 676718 196134 676954
rect 195514 656954 196134 676718
rect 195514 656718 195546 656954
rect 195782 656718 195866 656954
rect 196102 656718 196134 656954
rect 195514 636954 196134 656718
rect 195514 636718 195546 636954
rect 195782 636718 195866 636954
rect 196102 636718 196134 636954
rect 195514 616954 196134 636718
rect 195514 616718 195546 616954
rect 195782 616718 195866 616954
rect 196102 616718 196134 616954
rect 195514 596954 196134 616718
rect 195514 596718 195546 596954
rect 195782 596718 195866 596954
rect 196102 596718 196134 596954
rect 195514 576954 196134 596718
rect 195514 576718 195546 576954
rect 195782 576718 195866 576954
rect 196102 576718 196134 576954
rect 195514 556954 196134 576718
rect 195514 556718 195546 556954
rect 195782 556718 195866 556954
rect 196102 556718 196134 556954
rect 195514 536954 196134 556718
rect 195514 536718 195546 536954
rect 195782 536718 195866 536954
rect 196102 536718 196134 536954
rect 195514 516954 196134 536718
rect 195514 516718 195546 516954
rect 195782 516718 195866 516954
rect 196102 516718 196134 516954
rect 195514 496954 196134 516718
rect 195514 496718 195546 496954
rect 195782 496718 195866 496954
rect 196102 496718 196134 496954
rect 195514 476954 196134 496718
rect 195514 476718 195546 476954
rect 195782 476718 195866 476954
rect 196102 476718 196134 476954
rect 195514 456954 196134 476718
rect 196387 475420 196453 475421
rect 196387 475356 196388 475420
rect 196452 475356 196453 475420
rect 196387 475355 196453 475356
rect 195514 456718 195546 456954
rect 195782 456718 195866 456954
rect 196102 456718 196134 456954
rect 195514 436954 196134 456718
rect 196390 453253 196450 475355
rect 196387 453252 196453 453253
rect 196387 453188 196388 453252
rect 196452 453188 196453 453252
rect 196387 453187 196453 453188
rect 195514 436718 195546 436954
rect 195782 436718 195866 436954
rect 196102 436718 196134 436954
rect 195514 416954 196134 436718
rect 196574 432581 196634 700571
rect 199234 700378 199266 700614
rect 199502 700378 199586 700614
rect 199822 700378 199854 700614
rect 199234 680614 199854 700378
rect 199234 680378 199266 680614
rect 199502 680378 199586 680614
rect 199822 680378 199854 680614
rect 199234 660614 199854 680378
rect 199234 660378 199266 660614
rect 199502 660378 199586 660614
rect 199822 660378 199854 660614
rect 199234 640614 199854 660378
rect 199234 640378 199266 640614
rect 199502 640378 199586 640614
rect 199822 640378 199854 640614
rect 199234 620614 199854 640378
rect 199234 620378 199266 620614
rect 199502 620378 199586 620614
rect 199822 620378 199854 620614
rect 199234 600614 199854 620378
rect 199234 600378 199266 600614
rect 199502 600378 199586 600614
rect 199822 600378 199854 600614
rect 199234 580614 199854 600378
rect 199234 580378 199266 580614
rect 199502 580378 199586 580614
rect 199822 580378 199854 580614
rect 199234 560614 199854 580378
rect 199234 560378 199266 560614
rect 199502 560378 199586 560614
rect 199822 560378 199854 560614
rect 199234 540614 199854 560378
rect 199234 540378 199266 540614
rect 199502 540378 199586 540614
rect 199822 540378 199854 540614
rect 198595 539748 198661 539749
rect 198595 539684 198596 539748
rect 198660 539684 198661 539748
rect 198595 539683 198661 539684
rect 198043 475148 198109 475149
rect 198043 475084 198044 475148
rect 198108 475084 198109 475148
rect 198043 475083 198109 475084
rect 197859 474876 197925 474877
rect 197859 474812 197860 474876
rect 197924 474812 197925 474876
rect 197859 474811 197925 474812
rect 197307 455564 197373 455565
rect 197307 455500 197308 455564
rect 197372 455500 197373 455564
rect 197307 455499 197373 455500
rect 197310 452165 197370 455499
rect 197862 452709 197922 474811
rect 198046 452845 198106 475083
rect 198043 452844 198109 452845
rect 198043 452780 198044 452844
rect 198108 452780 198109 452844
rect 198043 452779 198109 452780
rect 197859 452708 197925 452709
rect 197859 452644 197860 452708
rect 197924 452644 197925 452708
rect 197859 452643 197925 452644
rect 197307 452164 197373 452165
rect 197307 452100 197308 452164
rect 197372 452100 197373 452164
rect 197307 452099 197373 452100
rect 196571 432580 196637 432581
rect 196571 432516 196572 432580
rect 196636 432516 196637 432580
rect 196571 432515 196637 432516
rect 195514 416718 195546 416954
rect 195782 416718 195866 416954
rect 196102 416718 196134 416954
rect 195514 396954 196134 416718
rect 195514 396718 195546 396954
rect 195782 396718 195866 396954
rect 196102 396718 196134 396954
rect 195514 376954 196134 396718
rect 195514 376718 195546 376954
rect 195782 376718 195866 376954
rect 196102 376718 196134 376954
rect 195514 356954 196134 376718
rect 195514 356718 195546 356954
rect 195782 356718 195866 356954
rect 196102 356718 196134 356954
rect 195514 336954 196134 356718
rect 195514 336718 195546 336954
rect 195782 336718 195866 336954
rect 196102 336718 196134 336954
rect 195514 316954 196134 336718
rect 195514 316718 195546 316954
rect 195782 316718 195866 316954
rect 196102 316718 196134 316954
rect 195514 296954 196134 316718
rect 195514 296718 195546 296954
rect 195782 296718 195866 296954
rect 196102 296718 196134 296954
rect 195514 276954 196134 296718
rect 195514 276718 195546 276954
rect 195782 276718 195866 276954
rect 196102 276718 196134 276954
rect 195514 256954 196134 276718
rect 195514 256718 195546 256954
rect 195782 256718 195866 256954
rect 196102 256718 196134 256954
rect 195514 236954 196134 256718
rect 198598 250477 198658 539683
rect 199234 539308 199854 540378
rect 201794 704838 202414 705830
rect 201794 704602 201826 704838
rect 202062 704602 202146 704838
rect 202382 704602 202414 704838
rect 201794 704518 202414 704602
rect 201794 704282 201826 704518
rect 202062 704282 202146 704518
rect 202382 704282 202414 704518
rect 201794 683294 202414 704282
rect 201794 683058 201826 683294
rect 202062 683058 202146 683294
rect 202382 683058 202414 683294
rect 201794 663294 202414 683058
rect 201794 663058 201826 663294
rect 202062 663058 202146 663294
rect 202382 663058 202414 663294
rect 201794 643294 202414 663058
rect 201794 643058 201826 643294
rect 202062 643058 202146 643294
rect 202382 643058 202414 643294
rect 201794 623294 202414 643058
rect 201794 623058 201826 623294
rect 202062 623058 202146 623294
rect 202382 623058 202414 623294
rect 201794 603294 202414 623058
rect 201794 603058 201826 603294
rect 202062 603058 202146 603294
rect 202382 603058 202414 603294
rect 201794 583294 202414 603058
rect 201794 583058 201826 583294
rect 202062 583058 202146 583294
rect 202382 583058 202414 583294
rect 201794 563294 202414 583058
rect 201794 563058 201826 563294
rect 202062 563058 202146 563294
rect 202382 563058 202414 563294
rect 201794 543294 202414 563058
rect 201794 543058 201826 543294
rect 202062 543058 202146 543294
rect 202382 543058 202414 543294
rect 201794 539308 202414 543058
rect 202954 684274 203574 711002
rect 212954 710598 213574 711590
rect 212954 710362 212986 710598
rect 213222 710362 213306 710598
rect 213542 710362 213574 710598
rect 212954 710278 213574 710362
rect 212954 710042 212986 710278
rect 213222 710042 213306 710278
rect 213542 710042 213574 710278
rect 209234 708678 209854 709670
rect 209234 708442 209266 708678
rect 209502 708442 209586 708678
rect 209822 708442 209854 708678
rect 209234 708358 209854 708442
rect 209234 708122 209266 708358
rect 209502 708122 209586 708358
rect 209822 708122 209854 708358
rect 202954 684038 202986 684274
rect 203222 684038 203306 684274
rect 203542 684038 203574 684274
rect 202954 664274 203574 684038
rect 202954 664038 202986 664274
rect 203222 664038 203306 664274
rect 203542 664038 203574 664274
rect 202954 644274 203574 664038
rect 202954 644038 202986 644274
rect 203222 644038 203306 644274
rect 203542 644038 203574 644274
rect 202954 624274 203574 644038
rect 202954 624038 202986 624274
rect 203222 624038 203306 624274
rect 203542 624038 203574 624274
rect 202954 604274 203574 624038
rect 202954 604038 202986 604274
rect 203222 604038 203306 604274
rect 203542 604038 203574 604274
rect 202954 584274 203574 604038
rect 202954 584038 202986 584274
rect 203222 584038 203306 584274
rect 203542 584038 203574 584274
rect 202954 564274 203574 584038
rect 202954 564038 202986 564274
rect 203222 564038 203306 564274
rect 203542 564038 203574 564274
rect 202954 544274 203574 564038
rect 202954 544038 202986 544274
rect 203222 544038 203306 544274
rect 203542 544038 203574 544274
rect 202954 539308 203574 544038
rect 205514 706758 206134 707750
rect 205514 706522 205546 706758
rect 205782 706522 205866 706758
rect 206102 706522 206134 706758
rect 205514 706438 206134 706522
rect 205514 706202 205546 706438
rect 205782 706202 205866 706438
rect 206102 706202 206134 706438
rect 205514 686954 206134 706202
rect 205514 686718 205546 686954
rect 205782 686718 205866 686954
rect 206102 686718 206134 686954
rect 205514 666954 206134 686718
rect 205514 666718 205546 666954
rect 205782 666718 205866 666954
rect 206102 666718 206134 666954
rect 205514 646954 206134 666718
rect 205514 646718 205546 646954
rect 205782 646718 205866 646954
rect 206102 646718 206134 646954
rect 205514 626954 206134 646718
rect 205514 626718 205546 626954
rect 205782 626718 205866 626954
rect 206102 626718 206134 626954
rect 205514 606954 206134 626718
rect 205514 606718 205546 606954
rect 205782 606718 205866 606954
rect 206102 606718 206134 606954
rect 205514 586954 206134 606718
rect 205514 586718 205546 586954
rect 205782 586718 205866 586954
rect 206102 586718 206134 586954
rect 205514 566954 206134 586718
rect 205514 566718 205546 566954
rect 205782 566718 205866 566954
rect 206102 566718 206134 566954
rect 205514 546954 206134 566718
rect 205514 546718 205546 546954
rect 205782 546718 205866 546954
rect 206102 546718 206134 546954
rect 205514 539308 206134 546718
rect 209234 690614 209854 708122
rect 209234 690378 209266 690614
rect 209502 690378 209586 690614
rect 209822 690378 209854 690614
rect 209234 670614 209854 690378
rect 209234 670378 209266 670614
rect 209502 670378 209586 670614
rect 209822 670378 209854 670614
rect 209234 650614 209854 670378
rect 209234 650378 209266 650614
rect 209502 650378 209586 650614
rect 209822 650378 209854 650614
rect 209234 630614 209854 650378
rect 209234 630378 209266 630614
rect 209502 630378 209586 630614
rect 209822 630378 209854 630614
rect 209234 610614 209854 630378
rect 209234 610378 209266 610614
rect 209502 610378 209586 610614
rect 209822 610378 209854 610614
rect 209234 590614 209854 610378
rect 209234 590378 209266 590614
rect 209502 590378 209586 590614
rect 209822 590378 209854 590614
rect 209234 570614 209854 590378
rect 209234 570378 209266 570614
rect 209502 570378 209586 570614
rect 209822 570378 209854 570614
rect 209234 550614 209854 570378
rect 209234 550378 209266 550614
rect 209502 550378 209586 550614
rect 209822 550378 209854 550614
rect 209234 539308 209854 550378
rect 211794 705798 212414 705830
rect 211794 705562 211826 705798
rect 212062 705562 212146 705798
rect 212382 705562 212414 705798
rect 211794 705478 212414 705562
rect 211794 705242 211826 705478
rect 212062 705242 212146 705478
rect 212382 705242 212414 705478
rect 211794 693294 212414 705242
rect 211794 693058 211826 693294
rect 212062 693058 212146 693294
rect 212382 693058 212414 693294
rect 211794 673294 212414 693058
rect 211794 673058 211826 673294
rect 212062 673058 212146 673294
rect 212382 673058 212414 673294
rect 211794 653294 212414 673058
rect 211794 653058 211826 653294
rect 212062 653058 212146 653294
rect 212382 653058 212414 653294
rect 211794 633294 212414 653058
rect 211794 633058 211826 633294
rect 212062 633058 212146 633294
rect 212382 633058 212414 633294
rect 211794 613294 212414 633058
rect 211794 613058 211826 613294
rect 212062 613058 212146 613294
rect 212382 613058 212414 613294
rect 211794 593294 212414 613058
rect 211794 593058 211826 593294
rect 212062 593058 212146 593294
rect 212382 593058 212414 593294
rect 211794 573294 212414 593058
rect 211794 573058 211826 573294
rect 212062 573058 212146 573294
rect 212382 573058 212414 573294
rect 211794 553294 212414 573058
rect 211794 553058 211826 553294
rect 212062 553058 212146 553294
rect 212382 553058 212414 553294
rect 211794 539308 212414 553058
rect 212954 694274 213574 710042
rect 222954 711558 223574 711590
rect 222954 711322 222986 711558
rect 223222 711322 223306 711558
rect 223542 711322 223574 711558
rect 222954 711238 223574 711322
rect 222954 711002 222986 711238
rect 223222 711002 223306 711238
rect 223542 711002 223574 711238
rect 219234 709638 219854 709670
rect 219234 709402 219266 709638
rect 219502 709402 219586 709638
rect 219822 709402 219854 709638
rect 219234 709318 219854 709402
rect 219234 709082 219266 709318
rect 219502 709082 219586 709318
rect 219822 709082 219854 709318
rect 212954 694038 212986 694274
rect 213222 694038 213306 694274
rect 213542 694038 213574 694274
rect 212954 674274 213574 694038
rect 212954 674038 212986 674274
rect 213222 674038 213306 674274
rect 213542 674038 213574 674274
rect 212954 654274 213574 674038
rect 212954 654038 212986 654274
rect 213222 654038 213306 654274
rect 213542 654038 213574 654274
rect 212954 634274 213574 654038
rect 212954 634038 212986 634274
rect 213222 634038 213306 634274
rect 213542 634038 213574 634274
rect 212954 614274 213574 634038
rect 212954 614038 212986 614274
rect 213222 614038 213306 614274
rect 213542 614038 213574 614274
rect 212954 594274 213574 614038
rect 212954 594038 212986 594274
rect 213222 594038 213306 594274
rect 213542 594038 213574 594274
rect 212954 574274 213574 594038
rect 212954 574038 212986 574274
rect 213222 574038 213306 574274
rect 213542 574038 213574 574274
rect 212954 554274 213574 574038
rect 212954 554038 212986 554274
rect 213222 554038 213306 554274
rect 213542 554038 213574 554274
rect 212954 539308 213574 554038
rect 215514 707718 216134 707750
rect 215514 707482 215546 707718
rect 215782 707482 215866 707718
rect 216102 707482 216134 707718
rect 215514 707398 216134 707482
rect 215514 707162 215546 707398
rect 215782 707162 215866 707398
rect 216102 707162 216134 707398
rect 215514 696954 216134 707162
rect 215514 696718 215546 696954
rect 215782 696718 215866 696954
rect 216102 696718 216134 696954
rect 215514 676954 216134 696718
rect 215514 676718 215546 676954
rect 215782 676718 215866 676954
rect 216102 676718 216134 676954
rect 215514 656954 216134 676718
rect 215514 656718 215546 656954
rect 215782 656718 215866 656954
rect 216102 656718 216134 656954
rect 215514 636954 216134 656718
rect 215514 636718 215546 636954
rect 215782 636718 215866 636954
rect 216102 636718 216134 636954
rect 215514 616954 216134 636718
rect 215514 616718 215546 616954
rect 215782 616718 215866 616954
rect 216102 616718 216134 616954
rect 215514 596954 216134 616718
rect 215514 596718 215546 596954
rect 215782 596718 215866 596954
rect 216102 596718 216134 596954
rect 215514 576954 216134 596718
rect 215514 576718 215546 576954
rect 215782 576718 215866 576954
rect 216102 576718 216134 576954
rect 215514 556954 216134 576718
rect 215514 556718 215546 556954
rect 215782 556718 215866 556954
rect 216102 556718 216134 556954
rect 215514 539308 216134 556718
rect 219234 700614 219854 709082
rect 219234 700378 219266 700614
rect 219502 700378 219586 700614
rect 219822 700378 219854 700614
rect 219234 680614 219854 700378
rect 219234 680378 219266 680614
rect 219502 680378 219586 680614
rect 219822 680378 219854 680614
rect 219234 660614 219854 680378
rect 219234 660378 219266 660614
rect 219502 660378 219586 660614
rect 219822 660378 219854 660614
rect 219234 640614 219854 660378
rect 219234 640378 219266 640614
rect 219502 640378 219586 640614
rect 219822 640378 219854 640614
rect 219234 620614 219854 640378
rect 219234 620378 219266 620614
rect 219502 620378 219586 620614
rect 219822 620378 219854 620614
rect 219234 600614 219854 620378
rect 219234 600378 219266 600614
rect 219502 600378 219586 600614
rect 219822 600378 219854 600614
rect 219234 580614 219854 600378
rect 219234 580378 219266 580614
rect 219502 580378 219586 580614
rect 219822 580378 219854 580614
rect 219234 560614 219854 580378
rect 219234 560378 219266 560614
rect 219502 560378 219586 560614
rect 219822 560378 219854 560614
rect 219234 540614 219854 560378
rect 219234 540378 219266 540614
rect 219502 540378 219586 540614
rect 219822 540378 219854 540614
rect 216811 539748 216877 539749
rect 216811 539684 216812 539748
rect 216876 539684 216877 539748
rect 216811 539683 216877 539684
rect 205771 539204 205837 539205
rect 205771 539140 205772 539204
rect 205836 539140 205837 539204
rect 205771 539139 205837 539140
rect 205774 537570 205834 539139
rect 205720 537510 205834 537570
rect 216814 537570 216874 539683
rect 218099 539612 218165 539613
rect 218099 539548 218100 539612
rect 218164 539548 218165 539612
rect 218099 539547 218165 539548
rect 218102 537570 218162 539547
rect 219234 539308 219854 540378
rect 221794 704838 222414 705830
rect 221794 704602 221826 704838
rect 222062 704602 222146 704838
rect 222382 704602 222414 704838
rect 221794 704518 222414 704602
rect 221794 704282 221826 704518
rect 222062 704282 222146 704518
rect 222382 704282 222414 704518
rect 221794 683294 222414 704282
rect 221794 683058 221826 683294
rect 222062 683058 222146 683294
rect 222382 683058 222414 683294
rect 221794 663294 222414 683058
rect 221794 663058 221826 663294
rect 222062 663058 222146 663294
rect 222382 663058 222414 663294
rect 221794 643294 222414 663058
rect 221794 643058 221826 643294
rect 222062 643058 222146 643294
rect 222382 643058 222414 643294
rect 221794 623294 222414 643058
rect 221794 623058 221826 623294
rect 222062 623058 222146 623294
rect 222382 623058 222414 623294
rect 221794 603294 222414 623058
rect 221794 603058 221826 603294
rect 222062 603058 222146 603294
rect 222382 603058 222414 603294
rect 221794 583294 222414 603058
rect 221794 583058 221826 583294
rect 222062 583058 222146 583294
rect 222382 583058 222414 583294
rect 221794 563294 222414 583058
rect 221794 563058 221826 563294
rect 222062 563058 222146 563294
rect 222382 563058 222414 563294
rect 221794 543294 222414 563058
rect 221794 543058 221826 543294
rect 222062 543058 222146 543294
rect 222382 543058 222414 543294
rect 221794 539308 222414 543058
rect 222954 684274 223574 711002
rect 232954 710598 233574 711590
rect 232954 710362 232986 710598
rect 233222 710362 233306 710598
rect 233542 710362 233574 710598
rect 232954 710278 233574 710362
rect 232954 710042 232986 710278
rect 233222 710042 233306 710278
rect 233542 710042 233574 710278
rect 229234 708678 229854 709670
rect 229234 708442 229266 708678
rect 229502 708442 229586 708678
rect 229822 708442 229854 708678
rect 229234 708358 229854 708442
rect 229234 708122 229266 708358
rect 229502 708122 229586 708358
rect 229822 708122 229854 708358
rect 222954 684038 222986 684274
rect 223222 684038 223306 684274
rect 223542 684038 223574 684274
rect 222954 664274 223574 684038
rect 222954 664038 222986 664274
rect 223222 664038 223306 664274
rect 223542 664038 223574 664274
rect 222954 644274 223574 664038
rect 222954 644038 222986 644274
rect 223222 644038 223306 644274
rect 223542 644038 223574 644274
rect 222954 624274 223574 644038
rect 222954 624038 222986 624274
rect 223222 624038 223306 624274
rect 223542 624038 223574 624274
rect 222954 604274 223574 624038
rect 222954 604038 222986 604274
rect 223222 604038 223306 604274
rect 223542 604038 223574 604274
rect 222954 584274 223574 604038
rect 222954 584038 222986 584274
rect 223222 584038 223306 584274
rect 223542 584038 223574 584274
rect 222954 564274 223574 584038
rect 222954 564038 222986 564274
rect 223222 564038 223306 564274
rect 223542 564038 223574 564274
rect 222954 544274 223574 564038
rect 222954 544038 222986 544274
rect 223222 544038 223306 544274
rect 223542 544038 223574 544274
rect 222954 539308 223574 544038
rect 225514 706758 226134 707750
rect 225514 706522 225546 706758
rect 225782 706522 225866 706758
rect 226102 706522 226134 706758
rect 225514 706438 226134 706522
rect 225514 706202 225546 706438
rect 225782 706202 225866 706438
rect 226102 706202 226134 706438
rect 225514 686954 226134 706202
rect 225514 686718 225546 686954
rect 225782 686718 225866 686954
rect 226102 686718 226134 686954
rect 225514 666954 226134 686718
rect 225514 666718 225546 666954
rect 225782 666718 225866 666954
rect 226102 666718 226134 666954
rect 225514 646954 226134 666718
rect 225514 646718 225546 646954
rect 225782 646718 225866 646954
rect 226102 646718 226134 646954
rect 225514 626954 226134 646718
rect 225514 626718 225546 626954
rect 225782 626718 225866 626954
rect 226102 626718 226134 626954
rect 225514 606954 226134 626718
rect 225514 606718 225546 606954
rect 225782 606718 225866 606954
rect 226102 606718 226134 606954
rect 225514 586954 226134 606718
rect 225514 586718 225546 586954
rect 225782 586718 225866 586954
rect 226102 586718 226134 586954
rect 225514 566954 226134 586718
rect 225514 566718 225546 566954
rect 225782 566718 225866 566954
rect 226102 566718 226134 566954
rect 225514 546954 226134 566718
rect 225514 546718 225546 546954
rect 225782 546718 225866 546954
rect 226102 546718 226134 546954
rect 225514 539308 226134 546718
rect 229234 690614 229854 708122
rect 229234 690378 229266 690614
rect 229502 690378 229586 690614
rect 229822 690378 229854 690614
rect 229234 670614 229854 690378
rect 229234 670378 229266 670614
rect 229502 670378 229586 670614
rect 229822 670378 229854 670614
rect 229234 650614 229854 670378
rect 229234 650378 229266 650614
rect 229502 650378 229586 650614
rect 229822 650378 229854 650614
rect 229234 630614 229854 650378
rect 229234 630378 229266 630614
rect 229502 630378 229586 630614
rect 229822 630378 229854 630614
rect 229234 610614 229854 630378
rect 229234 610378 229266 610614
rect 229502 610378 229586 610614
rect 229822 610378 229854 610614
rect 229234 590614 229854 610378
rect 229234 590378 229266 590614
rect 229502 590378 229586 590614
rect 229822 590378 229854 590614
rect 229234 570614 229854 590378
rect 229234 570378 229266 570614
rect 229502 570378 229586 570614
rect 229822 570378 229854 570614
rect 229234 550614 229854 570378
rect 229234 550378 229266 550614
rect 229502 550378 229586 550614
rect 229822 550378 229854 550614
rect 229234 539308 229854 550378
rect 231794 705798 232414 705830
rect 231794 705562 231826 705798
rect 232062 705562 232146 705798
rect 232382 705562 232414 705798
rect 231794 705478 232414 705562
rect 231794 705242 231826 705478
rect 232062 705242 232146 705478
rect 232382 705242 232414 705478
rect 231794 693294 232414 705242
rect 231794 693058 231826 693294
rect 232062 693058 232146 693294
rect 232382 693058 232414 693294
rect 231794 673294 232414 693058
rect 231794 673058 231826 673294
rect 232062 673058 232146 673294
rect 232382 673058 232414 673294
rect 231794 653294 232414 673058
rect 231794 653058 231826 653294
rect 232062 653058 232146 653294
rect 232382 653058 232414 653294
rect 231794 633294 232414 653058
rect 231794 633058 231826 633294
rect 232062 633058 232146 633294
rect 232382 633058 232414 633294
rect 231794 613294 232414 633058
rect 231794 613058 231826 613294
rect 232062 613058 232146 613294
rect 232382 613058 232414 613294
rect 231794 593294 232414 613058
rect 231794 593058 231826 593294
rect 232062 593058 232146 593294
rect 232382 593058 232414 593294
rect 231794 573294 232414 593058
rect 231794 573058 231826 573294
rect 232062 573058 232146 573294
rect 232382 573058 232414 573294
rect 231794 553294 232414 573058
rect 231794 553058 231826 553294
rect 232062 553058 232146 553294
rect 232382 553058 232414 553294
rect 231794 539308 232414 553058
rect 232954 694274 233574 710042
rect 242954 711558 243574 711590
rect 242954 711322 242986 711558
rect 243222 711322 243306 711558
rect 243542 711322 243574 711558
rect 242954 711238 243574 711322
rect 242954 711002 242986 711238
rect 243222 711002 243306 711238
rect 243542 711002 243574 711238
rect 239234 709638 239854 709670
rect 239234 709402 239266 709638
rect 239502 709402 239586 709638
rect 239822 709402 239854 709638
rect 239234 709318 239854 709402
rect 239234 709082 239266 709318
rect 239502 709082 239586 709318
rect 239822 709082 239854 709318
rect 232954 694038 232986 694274
rect 233222 694038 233306 694274
rect 233542 694038 233574 694274
rect 232954 674274 233574 694038
rect 232954 674038 232986 674274
rect 233222 674038 233306 674274
rect 233542 674038 233574 674274
rect 232954 654274 233574 674038
rect 232954 654038 232986 654274
rect 233222 654038 233306 654274
rect 233542 654038 233574 654274
rect 232954 634274 233574 654038
rect 232954 634038 232986 634274
rect 233222 634038 233306 634274
rect 233542 634038 233574 634274
rect 232954 614274 233574 634038
rect 232954 614038 232986 614274
rect 233222 614038 233306 614274
rect 233542 614038 233574 614274
rect 232954 594274 233574 614038
rect 232954 594038 232986 594274
rect 233222 594038 233306 594274
rect 233542 594038 233574 594274
rect 232954 574274 233574 594038
rect 232954 574038 232986 574274
rect 233222 574038 233306 574274
rect 233542 574038 233574 574274
rect 232954 554274 233574 574038
rect 232954 554038 232986 554274
rect 233222 554038 233306 554274
rect 233542 554038 233574 554274
rect 232954 539308 233574 554038
rect 235514 707718 236134 707750
rect 235514 707482 235546 707718
rect 235782 707482 235866 707718
rect 236102 707482 236134 707718
rect 235514 707398 236134 707482
rect 235514 707162 235546 707398
rect 235782 707162 235866 707398
rect 236102 707162 236134 707398
rect 235514 696954 236134 707162
rect 235514 696718 235546 696954
rect 235782 696718 235866 696954
rect 236102 696718 236134 696954
rect 235514 676954 236134 696718
rect 235514 676718 235546 676954
rect 235782 676718 235866 676954
rect 236102 676718 236134 676954
rect 235514 656954 236134 676718
rect 239234 700614 239854 709082
rect 239234 700378 239266 700614
rect 239502 700378 239586 700614
rect 239822 700378 239854 700614
rect 239234 680614 239854 700378
rect 239234 680378 239266 680614
rect 239502 680378 239586 680614
rect 239822 680378 239854 680614
rect 239234 660614 239854 680378
rect 239234 660378 239266 660614
rect 239502 660378 239586 660614
rect 239822 660378 239854 660614
rect 239234 659500 239854 660378
rect 241794 704838 242414 705830
rect 241794 704602 241826 704838
rect 242062 704602 242146 704838
rect 242382 704602 242414 704838
rect 241794 704518 242414 704602
rect 241794 704282 241826 704518
rect 242062 704282 242146 704518
rect 242382 704282 242414 704518
rect 241794 683294 242414 704282
rect 241794 683058 241826 683294
rect 242062 683058 242146 683294
rect 242382 683058 242414 683294
rect 241794 663294 242414 683058
rect 241794 663058 241826 663294
rect 242062 663058 242146 663294
rect 242382 663058 242414 663294
rect 241794 659500 242414 663058
rect 242954 684274 243574 711002
rect 252954 710598 253574 711590
rect 252954 710362 252986 710598
rect 253222 710362 253306 710598
rect 253542 710362 253574 710598
rect 252954 710278 253574 710362
rect 252954 710042 252986 710278
rect 253222 710042 253306 710278
rect 253542 710042 253574 710278
rect 249234 708678 249854 709670
rect 249234 708442 249266 708678
rect 249502 708442 249586 708678
rect 249822 708442 249854 708678
rect 249234 708358 249854 708442
rect 249234 708122 249266 708358
rect 249502 708122 249586 708358
rect 249822 708122 249854 708358
rect 242954 684038 242986 684274
rect 243222 684038 243306 684274
rect 243542 684038 243574 684274
rect 242954 664274 243574 684038
rect 242954 664038 242986 664274
rect 243222 664038 243306 664274
rect 243542 664038 243574 664274
rect 242954 659500 243574 664038
rect 245514 706758 246134 707750
rect 245514 706522 245546 706758
rect 245782 706522 245866 706758
rect 246102 706522 246134 706758
rect 245514 706438 246134 706522
rect 245514 706202 245546 706438
rect 245782 706202 245866 706438
rect 246102 706202 246134 706438
rect 245514 686954 246134 706202
rect 245514 686718 245546 686954
rect 245782 686718 245866 686954
rect 246102 686718 246134 686954
rect 245514 666954 246134 686718
rect 245514 666718 245546 666954
rect 245782 666718 245866 666954
rect 246102 666718 246134 666954
rect 245514 659500 246134 666718
rect 249234 690614 249854 708122
rect 249234 690378 249266 690614
rect 249502 690378 249586 690614
rect 249822 690378 249854 690614
rect 249234 670614 249854 690378
rect 249234 670378 249266 670614
rect 249502 670378 249586 670614
rect 249822 670378 249854 670614
rect 246251 659700 246317 659701
rect 246251 659636 246252 659700
rect 246316 659636 246317 659700
rect 246251 659635 246317 659636
rect 246254 657930 246314 659635
rect 249234 659500 249854 670378
rect 251794 705798 252414 705830
rect 251794 705562 251826 705798
rect 252062 705562 252146 705798
rect 252382 705562 252414 705798
rect 251794 705478 252414 705562
rect 251794 705242 251826 705478
rect 252062 705242 252146 705478
rect 252382 705242 252414 705478
rect 251794 693294 252414 705242
rect 251794 693058 251826 693294
rect 252062 693058 252146 693294
rect 252382 693058 252414 693294
rect 251794 673294 252414 693058
rect 251794 673058 251826 673294
rect 252062 673058 252146 673294
rect 252382 673058 252414 673294
rect 251794 659500 252414 673058
rect 252954 694274 253574 710042
rect 262954 711558 263574 711590
rect 262954 711322 262986 711558
rect 263222 711322 263306 711558
rect 263542 711322 263574 711558
rect 262954 711238 263574 711322
rect 262954 711002 262986 711238
rect 263222 711002 263306 711238
rect 263542 711002 263574 711238
rect 259234 709638 259854 709670
rect 259234 709402 259266 709638
rect 259502 709402 259586 709638
rect 259822 709402 259854 709638
rect 259234 709318 259854 709402
rect 259234 709082 259266 709318
rect 259502 709082 259586 709318
rect 259822 709082 259854 709318
rect 252954 694038 252986 694274
rect 253222 694038 253306 694274
rect 253542 694038 253574 694274
rect 252954 674274 253574 694038
rect 252954 674038 252986 674274
rect 253222 674038 253306 674274
rect 253542 674038 253574 674274
rect 252954 659500 253574 674038
rect 255514 707718 256134 707750
rect 255514 707482 255546 707718
rect 255782 707482 255866 707718
rect 256102 707482 256134 707718
rect 255514 707398 256134 707482
rect 255514 707162 255546 707398
rect 255782 707162 255866 707398
rect 256102 707162 256134 707398
rect 255514 696954 256134 707162
rect 255514 696718 255546 696954
rect 255782 696718 255866 696954
rect 256102 696718 256134 696954
rect 255514 676954 256134 696718
rect 255514 676718 255546 676954
rect 255782 676718 255866 676954
rect 256102 676718 256134 676954
rect 255514 659500 256134 676718
rect 259234 700614 259854 709082
rect 259234 700378 259266 700614
rect 259502 700378 259586 700614
rect 259822 700378 259854 700614
rect 259234 680614 259854 700378
rect 259234 680378 259266 680614
rect 259502 680378 259586 680614
rect 259822 680378 259854 680614
rect 259234 660614 259854 680378
rect 259234 660378 259266 660614
rect 259502 660378 259586 660614
rect 259822 660378 259854 660614
rect 256555 659700 256621 659701
rect 256555 659636 256556 659700
rect 256620 659636 256621 659700
rect 256555 659635 256621 659636
rect 256558 657930 256618 659635
rect 259234 659500 259854 660378
rect 261794 704838 262414 705830
rect 261794 704602 261826 704838
rect 262062 704602 262146 704838
rect 262382 704602 262414 704838
rect 261794 704518 262414 704602
rect 261794 704282 261826 704518
rect 262062 704282 262146 704518
rect 262382 704282 262414 704518
rect 261794 683294 262414 704282
rect 261794 683058 261826 683294
rect 262062 683058 262146 683294
rect 262382 683058 262414 683294
rect 261794 663294 262414 683058
rect 261794 663058 261826 663294
rect 262062 663058 262146 663294
rect 262382 663058 262414 663294
rect 261794 659500 262414 663058
rect 262954 684274 263574 711002
rect 272954 710598 273574 711590
rect 272954 710362 272986 710598
rect 273222 710362 273306 710598
rect 273542 710362 273574 710598
rect 272954 710278 273574 710362
rect 272954 710042 272986 710278
rect 273222 710042 273306 710278
rect 273542 710042 273574 710278
rect 269234 708678 269854 709670
rect 269234 708442 269266 708678
rect 269502 708442 269586 708678
rect 269822 708442 269854 708678
rect 269234 708358 269854 708442
rect 269234 708122 269266 708358
rect 269502 708122 269586 708358
rect 269822 708122 269854 708358
rect 262954 684038 262986 684274
rect 263222 684038 263306 684274
rect 263542 684038 263574 684274
rect 262954 664274 263574 684038
rect 262954 664038 262986 664274
rect 263222 664038 263306 664274
rect 263542 664038 263574 664274
rect 262954 659500 263574 664038
rect 265514 706758 266134 707750
rect 265514 706522 265546 706758
rect 265782 706522 265866 706758
rect 266102 706522 266134 706758
rect 265514 706438 266134 706522
rect 265514 706202 265546 706438
rect 265782 706202 265866 706438
rect 266102 706202 266134 706438
rect 265514 686954 266134 706202
rect 265514 686718 265546 686954
rect 265782 686718 265866 686954
rect 266102 686718 266134 686954
rect 265514 666954 266134 686718
rect 265514 666718 265546 666954
rect 265782 666718 265866 666954
rect 266102 666718 266134 666954
rect 265514 659500 266134 666718
rect 269234 690614 269854 708122
rect 269234 690378 269266 690614
rect 269502 690378 269586 690614
rect 269822 690378 269854 690614
rect 269234 670614 269854 690378
rect 269234 670378 269266 670614
rect 269502 670378 269586 670614
rect 269822 670378 269854 670614
rect 269234 659500 269854 670378
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 693294 272414 705242
rect 271794 693058 271826 693294
rect 272062 693058 272146 693294
rect 272382 693058 272414 693294
rect 271794 673294 272414 693058
rect 271794 673058 271826 673294
rect 272062 673058 272146 673294
rect 272382 673058 272414 673294
rect 271794 659500 272414 673058
rect 272954 694274 273574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 272954 694038 272986 694274
rect 273222 694038 273306 694274
rect 273542 694038 273574 694274
rect 272954 674274 273574 694038
rect 272954 674038 272986 674274
rect 273222 674038 273306 674274
rect 273542 674038 273574 674274
rect 272954 659500 273574 674038
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 275514 696954 276134 707162
rect 275514 696718 275546 696954
rect 275782 696718 275866 696954
rect 276102 696718 276134 696954
rect 275514 676954 276134 696718
rect 275514 676718 275546 676954
rect 275782 676718 275866 676954
rect 276102 676718 276134 676954
rect 275514 659500 276134 676718
rect 279234 700614 279854 709082
rect 279234 700378 279266 700614
rect 279502 700378 279586 700614
rect 279822 700378 279854 700614
rect 279234 680614 279854 700378
rect 279234 680378 279266 680614
rect 279502 680378 279586 680614
rect 279822 680378 279854 680614
rect 279234 660614 279854 680378
rect 279234 660378 279266 660614
rect 279502 660378 279586 660614
rect 279822 660378 279854 660614
rect 279234 659500 279854 660378
rect 281794 704838 282414 705830
rect 281794 704602 281826 704838
rect 282062 704602 282146 704838
rect 282382 704602 282414 704838
rect 281794 704518 282414 704602
rect 281794 704282 281826 704518
rect 282062 704282 282146 704518
rect 282382 704282 282414 704518
rect 281794 683294 282414 704282
rect 281794 683058 281826 683294
rect 282062 683058 282146 683294
rect 282382 683058 282414 683294
rect 281794 663294 282414 683058
rect 281794 663058 281826 663294
rect 282062 663058 282146 663294
rect 282382 663058 282414 663294
rect 281794 659500 282414 663058
rect 282954 684274 283574 711002
rect 292954 710598 293574 711590
rect 292954 710362 292986 710598
rect 293222 710362 293306 710598
rect 293542 710362 293574 710598
rect 292954 710278 293574 710362
rect 292954 710042 292986 710278
rect 293222 710042 293306 710278
rect 293542 710042 293574 710278
rect 289234 708678 289854 709670
rect 289234 708442 289266 708678
rect 289502 708442 289586 708678
rect 289822 708442 289854 708678
rect 289234 708358 289854 708442
rect 289234 708122 289266 708358
rect 289502 708122 289586 708358
rect 289822 708122 289854 708358
rect 282954 684038 282986 684274
rect 283222 684038 283306 684274
rect 283542 684038 283574 684274
rect 282954 664274 283574 684038
rect 282954 664038 282986 664274
rect 283222 664038 283306 664274
rect 283542 664038 283574 664274
rect 282954 659500 283574 664038
rect 285514 706758 286134 707750
rect 285514 706522 285546 706758
rect 285782 706522 285866 706758
rect 286102 706522 286134 706758
rect 285514 706438 286134 706522
rect 285514 706202 285546 706438
rect 285782 706202 285866 706438
rect 286102 706202 286134 706438
rect 285514 686954 286134 706202
rect 285514 686718 285546 686954
rect 285782 686718 285866 686954
rect 286102 686718 286134 686954
rect 285514 666954 286134 686718
rect 285514 666718 285546 666954
rect 285782 666718 285866 666954
rect 286102 666718 286134 666954
rect 285514 659500 286134 666718
rect 289234 690614 289854 708122
rect 289234 690378 289266 690614
rect 289502 690378 289586 690614
rect 289822 690378 289854 690614
rect 289234 670614 289854 690378
rect 289234 670378 289266 670614
rect 289502 670378 289586 670614
rect 289822 670378 289854 670614
rect 289234 659500 289854 670378
rect 291794 705798 292414 705830
rect 291794 705562 291826 705798
rect 292062 705562 292146 705798
rect 292382 705562 292414 705798
rect 291794 705478 292414 705562
rect 291794 705242 291826 705478
rect 292062 705242 292146 705478
rect 292382 705242 292414 705478
rect 291794 693294 292414 705242
rect 291794 693058 291826 693294
rect 292062 693058 292146 693294
rect 292382 693058 292414 693294
rect 291794 673294 292414 693058
rect 291794 673058 291826 673294
rect 292062 673058 292146 673294
rect 292382 673058 292414 673294
rect 291794 659500 292414 673058
rect 292954 694274 293574 710042
rect 302954 711558 303574 711590
rect 302954 711322 302986 711558
rect 303222 711322 303306 711558
rect 303542 711322 303574 711558
rect 302954 711238 303574 711322
rect 302954 711002 302986 711238
rect 303222 711002 303306 711238
rect 303542 711002 303574 711238
rect 299234 709638 299854 709670
rect 299234 709402 299266 709638
rect 299502 709402 299586 709638
rect 299822 709402 299854 709638
rect 299234 709318 299854 709402
rect 299234 709082 299266 709318
rect 299502 709082 299586 709318
rect 299822 709082 299854 709318
rect 292954 694038 292986 694274
rect 293222 694038 293306 694274
rect 293542 694038 293574 694274
rect 292954 674274 293574 694038
rect 292954 674038 292986 674274
rect 293222 674038 293306 674274
rect 293542 674038 293574 674274
rect 292954 659500 293574 674038
rect 295514 707718 296134 707750
rect 295514 707482 295546 707718
rect 295782 707482 295866 707718
rect 296102 707482 296134 707718
rect 295514 707398 296134 707482
rect 295514 707162 295546 707398
rect 295782 707162 295866 707398
rect 296102 707162 296134 707398
rect 295514 696954 296134 707162
rect 295514 696718 295546 696954
rect 295782 696718 295866 696954
rect 296102 696718 296134 696954
rect 295514 676954 296134 696718
rect 295514 676718 295546 676954
rect 295782 676718 295866 676954
rect 296102 676718 296134 676954
rect 295514 659500 296134 676718
rect 299234 700614 299854 709082
rect 299234 700378 299266 700614
rect 299502 700378 299586 700614
rect 299822 700378 299854 700614
rect 299234 680614 299854 700378
rect 299234 680378 299266 680614
rect 299502 680378 299586 680614
rect 299822 680378 299854 680614
rect 299234 660614 299854 680378
rect 299234 660378 299266 660614
rect 299502 660378 299586 660614
rect 299822 660378 299854 660614
rect 299234 659500 299854 660378
rect 301794 704838 302414 705830
rect 301794 704602 301826 704838
rect 302062 704602 302146 704838
rect 302382 704602 302414 704838
rect 301794 704518 302414 704602
rect 301794 704282 301826 704518
rect 302062 704282 302146 704518
rect 302382 704282 302414 704518
rect 301794 683294 302414 704282
rect 301794 683058 301826 683294
rect 302062 683058 302146 683294
rect 302382 683058 302414 683294
rect 301794 663294 302414 683058
rect 301794 663058 301826 663294
rect 302062 663058 302146 663294
rect 302382 663058 302414 663294
rect 301794 659500 302414 663058
rect 302954 684274 303574 711002
rect 312954 710598 313574 711590
rect 312954 710362 312986 710598
rect 313222 710362 313306 710598
rect 313542 710362 313574 710598
rect 312954 710278 313574 710362
rect 312954 710042 312986 710278
rect 313222 710042 313306 710278
rect 313542 710042 313574 710278
rect 309234 708678 309854 709670
rect 309234 708442 309266 708678
rect 309502 708442 309586 708678
rect 309822 708442 309854 708678
rect 309234 708358 309854 708442
rect 309234 708122 309266 708358
rect 309502 708122 309586 708358
rect 309822 708122 309854 708358
rect 302954 684038 302986 684274
rect 303222 684038 303306 684274
rect 303542 684038 303574 684274
rect 302954 664274 303574 684038
rect 302954 664038 302986 664274
rect 303222 664038 303306 664274
rect 303542 664038 303574 664274
rect 302954 659500 303574 664038
rect 305514 706758 306134 707750
rect 305514 706522 305546 706758
rect 305782 706522 305866 706758
rect 306102 706522 306134 706758
rect 305514 706438 306134 706522
rect 305514 706202 305546 706438
rect 305782 706202 305866 706438
rect 306102 706202 306134 706438
rect 305514 686954 306134 706202
rect 305514 686718 305546 686954
rect 305782 686718 305866 686954
rect 306102 686718 306134 686954
rect 305514 666954 306134 686718
rect 305514 666718 305546 666954
rect 305782 666718 305866 666954
rect 306102 666718 306134 666954
rect 305514 659500 306134 666718
rect 309234 690614 309854 708122
rect 309234 690378 309266 690614
rect 309502 690378 309586 690614
rect 309822 690378 309854 690614
rect 309234 670614 309854 690378
rect 309234 670378 309266 670614
rect 309502 670378 309586 670614
rect 309822 670378 309854 670614
rect 309234 659500 309854 670378
rect 311794 705798 312414 705830
rect 311794 705562 311826 705798
rect 312062 705562 312146 705798
rect 312382 705562 312414 705798
rect 311794 705478 312414 705562
rect 311794 705242 311826 705478
rect 312062 705242 312146 705478
rect 312382 705242 312414 705478
rect 311794 693294 312414 705242
rect 311794 693058 311826 693294
rect 312062 693058 312146 693294
rect 312382 693058 312414 693294
rect 311794 673294 312414 693058
rect 311794 673058 311826 673294
rect 312062 673058 312146 673294
rect 312382 673058 312414 673294
rect 311794 659500 312414 673058
rect 312954 694274 313574 710042
rect 322954 711558 323574 711590
rect 322954 711322 322986 711558
rect 323222 711322 323306 711558
rect 323542 711322 323574 711558
rect 322954 711238 323574 711322
rect 322954 711002 322986 711238
rect 323222 711002 323306 711238
rect 323542 711002 323574 711238
rect 319234 709638 319854 709670
rect 319234 709402 319266 709638
rect 319502 709402 319586 709638
rect 319822 709402 319854 709638
rect 319234 709318 319854 709402
rect 319234 709082 319266 709318
rect 319502 709082 319586 709318
rect 319822 709082 319854 709318
rect 312954 694038 312986 694274
rect 313222 694038 313306 694274
rect 313542 694038 313574 694274
rect 312954 674274 313574 694038
rect 312954 674038 312986 674274
rect 313222 674038 313306 674274
rect 313542 674038 313574 674274
rect 312954 659500 313574 674038
rect 315514 707718 316134 707750
rect 315514 707482 315546 707718
rect 315782 707482 315866 707718
rect 316102 707482 316134 707718
rect 315514 707398 316134 707482
rect 315514 707162 315546 707398
rect 315782 707162 315866 707398
rect 316102 707162 316134 707398
rect 315514 696954 316134 707162
rect 315514 696718 315546 696954
rect 315782 696718 315866 696954
rect 316102 696718 316134 696954
rect 315514 676954 316134 696718
rect 315514 676718 315546 676954
rect 315782 676718 315866 676954
rect 316102 676718 316134 676954
rect 315514 659500 316134 676718
rect 319234 700614 319854 709082
rect 319234 700378 319266 700614
rect 319502 700378 319586 700614
rect 319822 700378 319854 700614
rect 319234 680614 319854 700378
rect 319234 680378 319266 680614
rect 319502 680378 319586 680614
rect 319822 680378 319854 680614
rect 319234 660614 319854 680378
rect 319234 660378 319266 660614
rect 319502 660378 319586 660614
rect 319822 660378 319854 660614
rect 319234 659500 319854 660378
rect 321794 704838 322414 705830
rect 321794 704602 321826 704838
rect 322062 704602 322146 704838
rect 322382 704602 322414 704838
rect 321794 704518 322414 704602
rect 321794 704282 321826 704518
rect 322062 704282 322146 704518
rect 322382 704282 322414 704518
rect 321794 683294 322414 704282
rect 321794 683058 321826 683294
rect 322062 683058 322146 683294
rect 322382 683058 322414 683294
rect 321794 663294 322414 683058
rect 321794 663058 321826 663294
rect 322062 663058 322146 663294
rect 322382 663058 322414 663294
rect 321794 659500 322414 663058
rect 322954 684274 323574 711002
rect 332954 710598 333574 711590
rect 332954 710362 332986 710598
rect 333222 710362 333306 710598
rect 333542 710362 333574 710598
rect 332954 710278 333574 710362
rect 332954 710042 332986 710278
rect 333222 710042 333306 710278
rect 333542 710042 333574 710278
rect 329234 708678 329854 709670
rect 329234 708442 329266 708678
rect 329502 708442 329586 708678
rect 329822 708442 329854 708678
rect 329234 708358 329854 708442
rect 329234 708122 329266 708358
rect 329502 708122 329586 708358
rect 329822 708122 329854 708358
rect 322954 684038 322986 684274
rect 323222 684038 323306 684274
rect 323542 684038 323574 684274
rect 322954 664274 323574 684038
rect 322954 664038 322986 664274
rect 323222 664038 323306 664274
rect 323542 664038 323574 664274
rect 322954 659500 323574 664038
rect 325514 706758 326134 707750
rect 325514 706522 325546 706758
rect 325782 706522 325866 706758
rect 326102 706522 326134 706758
rect 325514 706438 326134 706522
rect 325514 706202 325546 706438
rect 325782 706202 325866 706438
rect 326102 706202 326134 706438
rect 325514 686954 326134 706202
rect 325514 686718 325546 686954
rect 325782 686718 325866 686954
rect 326102 686718 326134 686954
rect 325514 666954 326134 686718
rect 325514 666718 325546 666954
rect 325782 666718 325866 666954
rect 326102 666718 326134 666954
rect 325514 659500 326134 666718
rect 329234 690614 329854 708122
rect 329234 690378 329266 690614
rect 329502 690378 329586 690614
rect 329822 690378 329854 690614
rect 329234 670614 329854 690378
rect 329234 670378 329266 670614
rect 329502 670378 329586 670614
rect 329822 670378 329854 670614
rect 329234 659500 329854 670378
rect 331794 705798 332414 705830
rect 331794 705562 331826 705798
rect 332062 705562 332146 705798
rect 332382 705562 332414 705798
rect 331794 705478 332414 705562
rect 331794 705242 331826 705478
rect 332062 705242 332146 705478
rect 332382 705242 332414 705478
rect 331794 693294 332414 705242
rect 331794 693058 331826 693294
rect 332062 693058 332146 693294
rect 332382 693058 332414 693294
rect 331794 673294 332414 693058
rect 331794 673058 331826 673294
rect 332062 673058 332146 673294
rect 332382 673058 332414 673294
rect 331794 659500 332414 673058
rect 332954 694274 333574 710042
rect 342954 711558 343574 711590
rect 342954 711322 342986 711558
rect 343222 711322 343306 711558
rect 343542 711322 343574 711558
rect 342954 711238 343574 711322
rect 342954 711002 342986 711238
rect 343222 711002 343306 711238
rect 343542 711002 343574 711238
rect 339234 709638 339854 709670
rect 339234 709402 339266 709638
rect 339502 709402 339586 709638
rect 339822 709402 339854 709638
rect 339234 709318 339854 709402
rect 339234 709082 339266 709318
rect 339502 709082 339586 709318
rect 339822 709082 339854 709318
rect 332954 694038 332986 694274
rect 333222 694038 333306 694274
rect 333542 694038 333574 694274
rect 332954 674274 333574 694038
rect 332954 674038 332986 674274
rect 333222 674038 333306 674274
rect 333542 674038 333574 674274
rect 332954 659500 333574 674038
rect 335514 707718 336134 707750
rect 335514 707482 335546 707718
rect 335782 707482 335866 707718
rect 336102 707482 336134 707718
rect 335514 707398 336134 707482
rect 335514 707162 335546 707398
rect 335782 707162 335866 707398
rect 336102 707162 336134 707398
rect 335514 696954 336134 707162
rect 335514 696718 335546 696954
rect 335782 696718 335866 696954
rect 336102 696718 336134 696954
rect 335514 676954 336134 696718
rect 335514 676718 335546 676954
rect 335782 676718 335866 676954
rect 336102 676718 336134 676954
rect 335514 659500 336134 676718
rect 339234 700614 339854 709082
rect 339234 700378 339266 700614
rect 339502 700378 339586 700614
rect 339822 700378 339854 700614
rect 339234 680614 339854 700378
rect 339234 680378 339266 680614
rect 339502 680378 339586 680614
rect 339822 680378 339854 680614
rect 339234 660614 339854 680378
rect 339234 660378 339266 660614
rect 339502 660378 339586 660614
rect 339822 660378 339854 660614
rect 245856 657870 246314 657930
rect 256464 657870 256618 657930
rect 245856 657394 245916 657870
rect 256464 657394 256524 657870
rect 235514 656718 235546 656954
rect 235782 656718 235866 656954
rect 236102 656718 236134 656954
rect 235514 636954 236134 656718
rect 240272 653294 240620 653456
rect 240272 653058 240328 653294
rect 240564 653058 240620 653294
rect 240272 652896 240620 653058
rect 335336 653294 335684 653456
rect 335336 653058 335392 653294
rect 335628 653058 335684 653294
rect 335336 652896 335684 653058
rect 240952 643294 241300 643456
rect 240952 643058 241008 643294
rect 241244 643058 241300 643294
rect 240952 642896 241300 643058
rect 334656 643294 335004 643456
rect 334656 643058 334712 643294
rect 334948 643058 335004 643294
rect 334656 642896 335004 643058
rect 235514 636718 235546 636954
rect 235782 636718 235866 636954
rect 236102 636718 236134 636954
rect 235514 616954 236134 636718
rect 339234 640614 339854 660378
rect 341794 704838 342414 705830
rect 341794 704602 341826 704838
rect 342062 704602 342146 704838
rect 342382 704602 342414 704838
rect 341794 704518 342414 704602
rect 341794 704282 341826 704518
rect 342062 704282 342146 704518
rect 342382 704282 342414 704518
rect 341794 683294 342414 704282
rect 341794 683058 341826 683294
rect 342062 683058 342146 683294
rect 342382 683058 342414 683294
rect 341794 663294 342414 683058
rect 341794 663058 341826 663294
rect 342062 663058 342146 663294
rect 342382 663058 342414 663294
rect 340091 659700 340157 659701
rect 340091 659636 340092 659700
rect 340156 659636 340157 659700
rect 340091 659635 340157 659636
rect 339234 640378 339266 640614
rect 339502 640378 339586 640614
rect 339822 640378 339854 640614
rect 240272 633294 240620 633456
rect 240272 633058 240328 633294
rect 240564 633058 240620 633294
rect 240272 632896 240620 633058
rect 335336 633294 335684 633456
rect 335336 633058 335392 633294
rect 335628 633058 335684 633294
rect 335336 632896 335684 633058
rect 240952 623294 241300 623456
rect 240952 623058 241008 623294
rect 241244 623058 241300 623294
rect 240952 622896 241300 623058
rect 334656 623294 335004 623456
rect 334656 623058 334712 623294
rect 334948 623058 335004 623294
rect 334656 622896 335004 623058
rect 235514 616718 235546 616954
rect 235782 616718 235866 616954
rect 236102 616718 236134 616954
rect 235514 596954 236134 616718
rect 339234 620614 339854 640378
rect 339234 620378 339266 620614
rect 339502 620378 339586 620614
rect 339822 620378 339854 620614
rect 240272 613294 240620 613456
rect 240272 613058 240328 613294
rect 240564 613058 240620 613294
rect 240272 612896 240620 613058
rect 335336 613294 335684 613456
rect 335336 613058 335392 613294
rect 335628 613058 335684 613294
rect 335336 612896 335684 613058
rect 338251 612236 338317 612237
rect 338251 612172 338252 612236
rect 338316 612172 338317 612236
rect 338251 612171 338317 612172
rect 338067 611012 338133 611013
rect 338067 610948 338068 611012
rect 338132 610948 338133 611012
rect 338067 610947 338133 610948
rect 240952 603294 241300 603456
rect 240952 603058 241008 603294
rect 241244 603058 241300 603294
rect 240952 602896 241300 603058
rect 334656 603294 335004 603456
rect 334656 603058 334712 603294
rect 334948 603058 335004 603294
rect 334656 602896 335004 603058
rect 235514 596718 235546 596954
rect 235782 596718 235866 596954
rect 236102 596718 236134 596954
rect 235514 576954 236134 596718
rect 240272 593294 240620 593456
rect 240272 593058 240328 593294
rect 240564 593058 240620 593294
rect 240272 592896 240620 593058
rect 335336 593294 335684 593456
rect 335336 593058 335392 593294
rect 335628 593058 335684 593294
rect 335336 592896 335684 593058
rect 240952 583294 241300 583456
rect 240952 583058 241008 583294
rect 241244 583058 241300 583294
rect 240952 582896 241300 583058
rect 334656 583294 335004 583456
rect 334656 583058 334712 583294
rect 334948 583058 335004 583294
rect 334656 582896 335004 583058
rect 252507 577828 252573 577829
rect 252507 577764 252508 577828
rect 252572 577764 252573 577828
rect 252507 577763 252573 577764
rect 235514 576718 235546 576954
rect 235782 576718 235866 576954
rect 236102 576718 236134 576954
rect 235514 556954 236134 576718
rect 235514 556718 235546 556954
rect 235782 556718 235866 556954
rect 236102 556718 236134 556954
rect 235514 539308 236134 556718
rect 239234 560614 239854 576000
rect 239234 560378 239266 560614
rect 239502 560378 239586 560614
rect 239822 560378 239854 560614
rect 239234 540614 239854 560378
rect 239234 540378 239266 540614
rect 239502 540378 239586 540614
rect 239822 540378 239854 540614
rect 239234 539308 239854 540378
rect 241794 563294 242414 576000
rect 241794 563058 241826 563294
rect 242062 563058 242146 563294
rect 242382 563058 242414 563294
rect 241794 543294 242414 563058
rect 241794 543058 241826 543294
rect 242062 543058 242146 543294
rect 242382 543058 242414 543294
rect 241794 539308 242414 543058
rect 242954 564274 243574 576000
rect 242954 564038 242986 564274
rect 243222 564038 243306 564274
rect 243542 564038 243574 564274
rect 242954 544274 243574 564038
rect 242954 544038 242986 544274
rect 243222 544038 243306 544274
rect 243542 544038 243574 544274
rect 242954 539308 243574 544038
rect 245514 566954 246134 576000
rect 245514 566718 245546 566954
rect 245782 566718 245866 566954
rect 246102 566718 246134 566954
rect 245514 546954 246134 566718
rect 245514 546718 245546 546954
rect 245782 546718 245866 546954
rect 246102 546718 246134 546954
rect 245514 539308 246134 546718
rect 249234 570614 249854 576000
rect 249234 570378 249266 570614
rect 249502 570378 249586 570614
rect 249822 570378 249854 570614
rect 249234 550614 249854 570378
rect 249234 550378 249266 550614
rect 249502 550378 249586 550614
rect 249822 550378 249854 550614
rect 249234 539308 249854 550378
rect 251794 573294 252414 576000
rect 252510 574157 252570 577763
rect 252792 577690 252852 578000
rect 252928 577829 252988 578000
rect 252925 577828 252991 577829
rect 252925 577764 252926 577828
rect 252990 577764 252991 577828
rect 252925 577763 252991 577764
rect 253064 577690 253124 578000
rect 252792 577630 252938 577690
rect 252878 576870 252938 577630
rect 252694 576810 252938 576870
rect 253062 577630 253124 577690
rect 253200 577690 253260 578000
rect 269112 577690 269172 578000
rect 253200 577630 253858 577690
rect 252694 574293 252754 576810
rect 253062 576197 253122 577630
rect 253059 576196 253125 576197
rect 253059 576132 253060 576196
rect 253124 576132 253125 576196
rect 253059 576131 253125 576132
rect 252691 574292 252757 574293
rect 252691 574228 252692 574292
rect 252756 574228 252757 574292
rect 252691 574227 252757 574228
rect 252954 574274 253574 576000
rect 253798 574429 253858 577630
rect 269070 577630 269172 577690
rect 270336 577690 270396 578000
rect 271560 577690 271620 578000
rect 272784 577690 272844 578000
rect 270336 577630 270418 577690
rect 253795 574428 253861 574429
rect 253795 574364 253796 574428
rect 253860 574364 253861 574428
rect 253795 574363 253861 574364
rect 252507 574156 252573 574157
rect 252507 574092 252508 574156
rect 252572 574092 252573 574156
rect 252507 574091 252573 574092
rect 251794 573058 251826 573294
rect 252062 573058 252146 573294
rect 252382 573058 252414 573294
rect 251794 553294 252414 573058
rect 251794 553058 251826 553294
rect 252062 553058 252146 553294
rect 252382 553058 252414 553294
rect 251794 539308 252414 553058
rect 252954 574038 252986 574274
rect 253222 574038 253306 574274
rect 253542 574038 253574 574274
rect 252954 554274 253574 574038
rect 252954 554038 252986 554274
rect 253222 554038 253306 554274
rect 253542 554038 253574 554274
rect 252954 539308 253574 554038
rect 255514 556954 256134 576000
rect 255514 556718 255546 556954
rect 255782 556718 255866 556954
rect 256102 556718 256134 556954
rect 255514 539308 256134 556718
rect 259234 560614 259854 576000
rect 259234 560378 259266 560614
rect 259502 560378 259586 560614
rect 259822 560378 259854 560614
rect 259234 540614 259854 560378
rect 259234 540378 259266 540614
rect 259502 540378 259586 540614
rect 259822 540378 259854 540614
rect 259234 539308 259854 540378
rect 261794 563294 262414 576000
rect 261794 563058 261826 563294
rect 262062 563058 262146 563294
rect 262382 563058 262414 563294
rect 261794 543294 262414 563058
rect 261794 543058 261826 543294
rect 262062 543058 262146 543294
rect 262382 543058 262414 543294
rect 261794 539308 262414 543058
rect 262954 564274 263574 576000
rect 262954 564038 262986 564274
rect 263222 564038 263306 564274
rect 263542 564038 263574 564274
rect 262954 544274 263574 564038
rect 262954 544038 262986 544274
rect 263222 544038 263306 544274
rect 263542 544038 263574 544274
rect 262954 539308 263574 544038
rect 265514 566954 266134 576000
rect 269070 574157 269130 577630
rect 269067 574156 269133 574157
rect 269067 574092 269068 574156
rect 269132 574092 269133 574156
rect 269067 574091 269133 574092
rect 265514 566718 265546 566954
rect 265782 566718 265866 566954
rect 266102 566718 266134 566954
rect 265514 546954 266134 566718
rect 265514 546718 265546 546954
rect 265782 546718 265866 546954
rect 266102 546718 266134 546954
rect 265514 539308 266134 546718
rect 269234 570614 269854 576000
rect 270358 574293 270418 577630
rect 271462 577630 271620 577690
rect 272750 577630 272844 577690
rect 274008 577690 274068 578000
rect 275368 577690 275428 578000
rect 274008 577630 274098 577690
rect 270355 574292 270421 574293
rect 270355 574228 270356 574292
rect 270420 574228 270421 574292
rect 270355 574227 270421 574228
rect 271462 574157 271522 577630
rect 271459 574156 271525 574157
rect 271459 574092 271460 574156
rect 271524 574092 271525 574156
rect 271459 574091 271525 574092
rect 269234 570378 269266 570614
rect 269502 570378 269586 570614
rect 269822 570378 269854 570614
rect 269234 550614 269854 570378
rect 269234 550378 269266 550614
rect 269502 550378 269586 550614
rect 269822 550378 269854 550614
rect 269234 539308 269854 550378
rect 271794 573294 272414 576000
rect 272750 574157 272810 577630
rect 272954 574274 273574 576000
rect 274038 574429 274098 577630
rect 275326 577630 275428 577690
rect 276592 577690 276652 578000
rect 278088 577690 278148 578000
rect 276592 577630 276674 577690
rect 274035 574428 274101 574429
rect 274035 574364 274036 574428
rect 274100 574364 274101 574428
rect 274035 574363 274101 574364
rect 275326 574293 275386 577630
rect 272747 574156 272813 574157
rect 272747 574092 272748 574156
rect 272812 574092 272813 574156
rect 272747 574091 272813 574092
rect 271794 573058 271826 573294
rect 272062 573058 272146 573294
rect 272382 573058 272414 573294
rect 271794 553294 272414 573058
rect 271794 553058 271826 553294
rect 272062 553058 272146 553294
rect 272382 553058 272414 553294
rect 271794 539308 272414 553058
rect 272954 574038 272986 574274
rect 273222 574038 273306 574274
rect 273542 574038 273574 574274
rect 275323 574292 275389 574293
rect 275323 574228 275324 574292
rect 275388 574228 275389 574292
rect 275323 574227 275389 574228
rect 272954 554274 273574 574038
rect 272954 554038 272986 554274
rect 273222 554038 273306 554274
rect 273542 554038 273574 554274
rect 272954 539308 273574 554038
rect 275514 556954 276134 576000
rect 276614 574429 276674 577630
rect 278086 577630 278148 577690
rect 278224 577690 278284 578000
rect 279040 577690 279100 578000
rect 279312 577690 279372 578000
rect 278224 577630 278330 577690
rect 276611 574428 276677 574429
rect 276611 574364 276612 574428
rect 276676 574364 276677 574428
rect 276611 574363 276677 574364
rect 278086 574157 278146 577630
rect 278270 574157 278330 577630
rect 278822 577630 279100 577690
rect 279190 577630 279372 577690
rect 280264 577690 280324 578000
rect 280672 577690 280732 578000
rect 280264 577630 280354 577690
rect 278822 574293 278882 577630
rect 279190 576870 279250 577630
rect 280107 577556 280173 577557
rect 280107 577492 280108 577556
rect 280172 577492 280173 577556
rect 280107 577491 280173 577492
rect 279006 576810 279250 576870
rect 278819 574292 278885 574293
rect 278819 574228 278820 574292
rect 278884 574228 278885 574292
rect 278819 574227 278885 574228
rect 279006 574157 279066 576810
rect 278083 574156 278149 574157
rect 278083 574092 278084 574156
rect 278148 574092 278149 574156
rect 278083 574091 278149 574092
rect 278267 574156 278333 574157
rect 278267 574092 278268 574156
rect 278332 574092 278333 574156
rect 278267 574091 278333 574092
rect 279003 574156 279069 574157
rect 279003 574092 279004 574156
rect 279068 574092 279069 574156
rect 279003 574091 279069 574092
rect 275514 556718 275546 556954
rect 275782 556718 275866 556954
rect 276102 556718 276134 556954
rect 275514 539308 276134 556718
rect 279234 560614 279854 576000
rect 280110 575109 280170 577491
rect 280107 575108 280173 575109
rect 280107 575044 280108 575108
rect 280172 575044 280173 575108
rect 280107 575043 280173 575044
rect 280294 574973 280354 577630
rect 280662 577630 280732 577690
rect 280291 574972 280357 574973
rect 280291 574908 280292 574972
rect 280356 574908 280357 574972
rect 280291 574907 280357 574908
rect 280662 574157 280722 577630
rect 281488 577557 281548 578000
rect 281896 577690 281956 578000
rect 282712 577690 282772 578000
rect 281896 577630 282562 577690
rect 281485 577556 281551 577557
rect 281485 577492 281486 577556
rect 281550 577492 281551 577556
rect 281485 577491 281551 577492
rect 280659 574156 280725 574157
rect 280659 574092 280660 574156
rect 280724 574092 280725 574156
rect 280659 574091 280725 574092
rect 279234 560378 279266 560614
rect 279502 560378 279586 560614
rect 279822 560378 279854 560614
rect 279234 540614 279854 560378
rect 279234 540378 279266 540614
rect 279502 540378 279586 540614
rect 279822 540378 279854 540614
rect 279234 539308 279854 540378
rect 281794 563294 282414 576000
rect 282502 574157 282562 577630
rect 282686 577630 282772 577690
rect 282984 577690 283044 578000
rect 284072 577690 284132 578000
rect 284480 577690 284540 578000
rect 284891 577828 284957 577829
rect 284891 577764 284892 577828
rect 284956 577764 284957 577828
rect 284891 577763 284957 577764
rect 282984 577630 283850 577690
rect 284072 577630 284218 577690
rect 284480 577630 284586 577690
rect 282686 574973 282746 577630
rect 282683 574972 282749 574973
rect 282683 574908 282684 574972
rect 282748 574908 282749 574972
rect 282683 574907 282749 574908
rect 282499 574156 282565 574157
rect 282499 574092 282500 574156
rect 282564 574092 282565 574156
rect 282499 574091 282565 574092
rect 281794 563058 281826 563294
rect 282062 563058 282146 563294
rect 282382 563058 282414 563294
rect 281794 543294 282414 563058
rect 281794 543058 281826 543294
rect 282062 543058 282146 543294
rect 282382 543058 282414 543294
rect 281794 539308 282414 543058
rect 282954 564274 283574 576000
rect 283790 574157 283850 577630
rect 284158 575381 284218 577630
rect 284155 575380 284221 575381
rect 284155 575316 284156 575380
rect 284220 575316 284221 575380
rect 284155 575315 284221 575316
rect 284526 574837 284586 577630
rect 284894 575245 284954 577763
rect 285160 577690 285220 578000
rect 285296 577829 285356 578000
rect 285293 577828 285359 577829
rect 285293 577764 285294 577828
rect 285358 577764 285359 577828
rect 285293 577763 285359 577764
rect 286520 577690 286580 578000
rect 286792 577690 286852 578000
rect 285160 577630 285322 577690
rect 286520 577630 286610 577690
rect 285262 575381 285322 577630
rect 285259 575380 285325 575381
rect 285259 575316 285260 575380
rect 285324 575316 285325 575380
rect 285259 575315 285325 575316
rect 284891 575244 284957 575245
rect 284891 575180 284892 575244
rect 284956 575180 284957 575244
rect 284891 575179 284957 575180
rect 284523 574836 284589 574837
rect 284523 574772 284524 574836
rect 284588 574772 284589 574836
rect 284523 574771 284589 574772
rect 283787 574156 283853 574157
rect 283787 574092 283788 574156
rect 283852 574092 283853 574156
rect 283787 574091 283853 574092
rect 282954 564038 282986 564274
rect 283222 564038 283306 564274
rect 283542 564038 283574 564274
rect 282954 544274 283574 564038
rect 282954 544038 282986 544274
rect 283222 544038 283306 544274
rect 283542 544038 283574 544274
rect 282954 539308 283574 544038
rect 285514 566954 286134 576000
rect 286550 575381 286610 577630
rect 286734 577630 286852 577690
rect 287608 577690 287668 578000
rect 288016 577690 288076 578000
rect 288832 577690 288892 578000
rect 289240 577690 289300 578000
rect 287608 577630 287714 577690
rect 288016 577630 288082 577690
rect 288832 577630 289002 577690
rect 286547 575380 286613 575381
rect 286547 575316 286548 575380
rect 286612 575316 286613 575380
rect 286547 575315 286613 575316
rect 286734 574293 286794 577630
rect 287654 575381 287714 577630
rect 287651 575380 287717 575381
rect 287651 575316 287652 575380
rect 287716 575316 287717 575380
rect 287651 575315 287717 575316
rect 288022 574973 288082 577630
rect 288942 576870 289002 577630
rect 288758 576810 289002 576870
rect 289126 577630 289300 577690
rect 289920 577690 289980 578000
rect 290328 577690 290388 578000
rect 291008 577690 291068 578000
rect 291552 577690 291612 578000
rect 289920 577630 290106 577690
rect 288019 574972 288085 574973
rect 288019 574908 288020 574972
rect 288084 574908 288085 574972
rect 288019 574907 288085 574908
rect 288758 574565 288818 576810
rect 289126 576330 289186 577630
rect 288942 576270 289186 576330
rect 288942 574837 289002 576270
rect 288939 574836 289005 574837
rect 288939 574772 288940 574836
rect 289004 574772 289005 574836
rect 288939 574771 289005 574772
rect 288755 574564 288821 574565
rect 288755 574500 288756 574564
rect 288820 574500 288821 574564
rect 288755 574499 288821 574500
rect 286731 574292 286797 574293
rect 286731 574228 286732 574292
rect 286796 574228 286797 574292
rect 286731 574227 286797 574228
rect 285514 566718 285546 566954
rect 285782 566718 285866 566954
rect 286102 566718 286134 566954
rect 285514 546954 286134 566718
rect 285514 546718 285546 546954
rect 285782 546718 285866 546954
rect 286102 546718 286134 546954
rect 285514 539308 286134 546718
rect 289234 570614 289854 576000
rect 290046 574973 290106 577630
rect 290230 577630 290388 577690
rect 290966 577630 291068 577690
rect 291518 577630 291612 577690
rect 292368 577690 292428 578000
rect 292776 577690 292836 578000
rect 293456 577690 293516 578000
rect 294000 577690 294060 578000
rect 292368 577630 292498 577690
rect 292776 577630 292866 577690
rect 293456 577630 293786 577690
rect 290230 575245 290290 577630
rect 290227 575244 290293 575245
rect 290227 575180 290228 575244
rect 290292 575180 290293 575244
rect 290227 575179 290293 575180
rect 290043 574972 290109 574973
rect 290043 574908 290044 574972
rect 290108 574908 290109 574972
rect 290043 574907 290109 574908
rect 290966 574837 291026 577630
rect 291518 575109 291578 577630
rect 292438 576197 292498 577630
rect 292435 576196 292501 576197
rect 292435 576132 292436 576196
rect 292500 576132 292501 576196
rect 292435 576131 292501 576132
rect 291515 575108 291581 575109
rect 291515 575044 291516 575108
rect 291580 575044 291581 575108
rect 291515 575043 291581 575044
rect 290963 574836 291029 574837
rect 290963 574772 290964 574836
rect 291028 574772 291029 574836
rect 290963 574771 291029 574772
rect 289234 570378 289266 570614
rect 289502 570378 289586 570614
rect 289822 570378 289854 570614
rect 289234 550614 289854 570378
rect 289234 550378 289266 550614
rect 289502 550378 289586 550614
rect 289822 550378 289854 550614
rect 289234 539308 289854 550378
rect 291794 573294 292414 576000
rect 292806 574837 292866 577630
rect 292803 574836 292869 574837
rect 292803 574772 292804 574836
rect 292868 574772 292869 574836
rect 292803 574771 292869 574772
rect 291794 573058 291826 573294
rect 292062 573058 292146 573294
rect 292382 573058 292414 573294
rect 291794 553294 292414 573058
rect 291794 553058 291826 553294
rect 292062 553058 292146 553294
rect 292382 553058 292414 553294
rect 291794 539308 292414 553058
rect 292954 574274 293574 576000
rect 293726 574429 293786 577630
rect 293910 577630 294060 577690
rect 294544 577690 294604 578000
rect 295224 577690 295284 578000
rect 294544 577630 294706 577690
rect 293910 575245 293970 577630
rect 293907 575244 293973 575245
rect 293907 575180 293908 575244
rect 293972 575180 293973 575244
rect 293907 575179 293973 575180
rect 294646 574429 294706 577630
rect 295198 577630 295284 577690
rect 295632 577690 295692 578000
rect 296584 577690 296644 578000
rect 295632 577630 296362 577690
rect 295198 575109 295258 577630
rect 295195 575108 295261 575109
rect 295195 575044 295196 575108
rect 295260 575044 295261 575108
rect 295195 575043 295261 575044
rect 293723 574428 293789 574429
rect 293723 574364 293724 574428
rect 293788 574364 293789 574428
rect 293723 574363 293789 574364
rect 294643 574428 294709 574429
rect 294643 574364 294644 574428
rect 294708 574364 294709 574428
rect 294643 574363 294709 574364
rect 292954 574038 292986 574274
rect 293222 574038 293306 574274
rect 293542 574038 293574 574274
rect 292954 554274 293574 574038
rect 292954 554038 292986 554274
rect 293222 554038 293306 554274
rect 293542 554038 293574 554274
rect 292954 539308 293574 554038
rect 295514 556954 296134 576000
rect 296302 574565 296362 577630
rect 296486 577630 296644 577690
rect 296992 577690 297052 578000
rect 296992 577630 297098 577690
rect 296299 574564 296365 574565
rect 296299 574500 296300 574564
rect 296364 574500 296365 574564
rect 296299 574499 296365 574500
rect 296486 574157 296546 577630
rect 297038 575381 297098 577630
rect 298080 577010 298140 578000
rect 298216 577690 298276 578000
rect 299032 577690 299092 578000
rect 299304 577690 299364 578000
rect 300256 577690 300316 578000
rect 298216 577630 298386 577690
rect 298080 576950 298202 577010
rect 297035 575380 297101 575381
rect 297035 575316 297036 575380
rect 297100 575316 297101 575380
rect 297035 575315 297101 575316
rect 298142 574157 298202 576950
rect 298326 574565 298386 577630
rect 298878 577630 299092 577690
rect 299246 577630 299364 577690
rect 300166 577630 300316 577690
rect 300392 577690 300452 578000
rect 301480 577690 301540 578000
rect 301752 577690 301812 578000
rect 302704 577690 302764 578000
rect 300392 577630 300594 577690
rect 298323 574564 298389 574565
rect 298323 574500 298324 574564
rect 298388 574500 298389 574564
rect 298323 574499 298389 574500
rect 298878 574293 298938 577630
rect 299246 576870 299306 577630
rect 299062 576810 299306 576870
rect 299062 574565 299122 576810
rect 299059 574564 299125 574565
rect 299059 574500 299060 574564
rect 299124 574500 299125 574564
rect 299059 574499 299125 574500
rect 298875 574292 298941 574293
rect 298875 574228 298876 574292
rect 298940 574228 298941 574292
rect 298875 574227 298941 574228
rect 296483 574156 296549 574157
rect 296483 574092 296484 574156
rect 296548 574092 296549 574156
rect 296483 574091 296549 574092
rect 298139 574156 298205 574157
rect 298139 574092 298140 574156
rect 298204 574092 298205 574156
rect 298139 574091 298205 574092
rect 295514 556718 295546 556954
rect 295782 556718 295866 556954
rect 296102 556718 296134 556954
rect 295514 539308 296134 556718
rect 299234 560614 299854 576000
rect 300166 574565 300226 577630
rect 300534 575381 300594 577630
rect 301454 577630 301540 577690
rect 301638 577630 301812 577690
rect 302558 577630 302764 577690
rect 302840 577690 302900 578000
rect 303928 577690 303988 578000
rect 302840 577630 302986 577690
rect 300531 575380 300597 575381
rect 300531 575316 300532 575380
rect 300596 575316 300597 575380
rect 300531 575315 300597 575316
rect 300163 574564 300229 574565
rect 300163 574500 300164 574564
rect 300228 574500 300229 574564
rect 300163 574499 300229 574500
rect 301454 574157 301514 577630
rect 301638 575381 301698 577630
rect 301635 575380 301701 575381
rect 301635 575316 301636 575380
rect 301700 575316 301701 575380
rect 301635 575315 301701 575316
rect 301451 574156 301517 574157
rect 301451 574092 301452 574156
rect 301516 574092 301517 574156
rect 301451 574091 301517 574092
rect 299234 560378 299266 560614
rect 299502 560378 299586 560614
rect 299822 560378 299854 560614
rect 299234 540614 299854 560378
rect 299234 540378 299266 540614
rect 299502 540378 299586 540614
rect 299822 540378 299854 540614
rect 299234 539308 299854 540378
rect 301794 563294 302414 576000
rect 302558 574157 302618 577630
rect 302926 576870 302986 577630
rect 302742 576810 302986 576870
rect 303846 577630 303988 577690
rect 304064 577690 304124 578000
rect 305152 577690 305212 578000
rect 305560 577690 305620 578000
rect 306240 577690 306300 578000
rect 306648 577690 306708 578000
rect 307600 577690 307660 578000
rect 308008 577690 308068 578000
rect 308688 577690 308748 578000
rect 304064 577630 304274 577690
rect 302742 575381 302802 576810
rect 302739 575380 302805 575381
rect 302739 575316 302740 575380
rect 302804 575316 302805 575380
rect 302739 575315 302805 575316
rect 302555 574156 302621 574157
rect 302555 574092 302556 574156
rect 302620 574092 302621 574156
rect 302555 574091 302621 574092
rect 301794 563058 301826 563294
rect 302062 563058 302146 563294
rect 302382 563058 302414 563294
rect 301794 543294 302414 563058
rect 301794 543058 301826 543294
rect 302062 543058 302146 543294
rect 302382 543058 302414 543294
rect 301794 539308 302414 543058
rect 302954 564274 303574 576000
rect 303846 574293 303906 577630
rect 304214 575381 304274 577630
rect 305134 577630 305212 577690
rect 305318 577630 305620 577690
rect 306238 577630 306300 577690
rect 306606 577630 306708 577690
rect 307526 577630 307660 577690
rect 307894 577630 308068 577690
rect 308630 577630 308748 577690
rect 309776 577690 309836 578000
rect 310864 577690 310924 578000
rect 309776 577630 310162 577690
rect 305134 575381 305194 577630
rect 304211 575380 304277 575381
rect 304211 575316 304212 575380
rect 304276 575316 304277 575380
rect 304211 575315 304277 575316
rect 305131 575380 305197 575381
rect 305131 575316 305132 575380
rect 305196 575316 305197 575380
rect 305131 575315 305197 575316
rect 303843 574292 303909 574293
rect 303843 574228 303844 574292
rect 303908 574228 303909 574292
rect 303843 574227 303909 574228
rect 305318 574157 305378 577630
rect 305315 574156 305381 574157
rect 305315 574092 305316 574156
rect 305380 574092 305381 574156
rect 305315 574091 305381 574092
rect 302954 564038 302986 564274
rect 303222 564038 303306 564274
rect 303542 564038 303574 564274
rect 302954 544274 303574 564038
rect 302954 544038 302986 544274
rect 303222 544038 303306 544274
rect 303542 544038 303574 544274
rect 302954 539308 303574 544038
rect 305514 566954 306134 576000
rect 306238 575381 306298 577630
rect 306235 575380 306301 575381
rect 306235 575316 306236 575380
rect 306300 575316 306301 575380
rect 306235 575315 306301 575316
rect 306606 574157 306666 577630
rect 307526 575381 307586 577630
rect 307523 575380 307589 575381
rect 307523 575316 307524 575380
rect 307588 575316 307589 575380
rect 307523 575315 307589 575316
rect 307894 574701 307954 577630
rect 308630 574701 308690 577630
rect 307891 574700 307957 574701
rect 307891 574636 307892 574700
rect 307956 574636 307957 574700
rect 307891 574635 307957 574636
rect 308627 574700 308693 574701
rect 308627 574636 308628 574700
rect 308692 574636 308693 574700
rect 308627 574635 308693 574636
rect 306603 574156 306669 574157
rect 306603 574092 306604 574156
rect 306668 574092 306669 574156
rect 306603 574091 306669 574092
rect 305514 566718 305546 566954
rect 305782 566718 305866 566954
rect 306102 566718 306134 566954
rect 305514 546954 306134 566718
rect 305514 546718 305546 546954
rect 305782 546718 305866 546954
rect 306102 546718 306134 546954
rect 305514 539308 306134 546718
rect 309234 570614 309854 576000
rect 310102 574837 310162 577630
rect 310838 577630 310924 577690
rect 312224 577690 312284 578000
rect 313312 577690 313372 578000
rect 314536 577690 314596 578000
rect 312224 577630 312738 577690
rect 313312 577630 313842 577690
rect 310838 574973 310898 577630
rect 310835 574972 310901 574973
rect 310835 574908 310836 574972
rect 310900 574908 310901 574972
rect 310835 574907 310901 574908
rect 310099 574836 310165 574837
rect 310099 574772 310100 574836
rect 310164 574772 310165 574836
rect 310099 574771 310165 574772
rect 309234 570378 309266 570614
rect 309502 570378 309586 570614
rect 309822 570378 309854 570614
rect 309234 550614 309854 570378
rect 309234 550378 309266 550614
rect 309502 550378 309586 550614
rect 309822 550378 309854 550614
rect 309234 539308 309854 550378
rect 311794 573294 312414 576000
rect 312678 575109 312738 577630
rect 312675 575108 312741 575109
rect 312675 575044 312676 575108
rect 312740 575044 312741 575108
rect 312675 575043 312741 575044
rect 311794 573058 311826 573294
rect 312062 573058 312146 573294
rect 312382 573058 312414 573294
rect 311794 553294 312414 573058
rect 311794 553058 311826 553294
rect 312062 553058 312146 553294
rect 312382 553058 312414 553294
rect 311794 539308 312414 553058
rect 312954 574274 313574 576000
rect 313782 574293 313842 577630
rect 314518 577630 314596 577690
rect 315760 577690 315820 578000
rect 316712 577690 316772 578000
rect 318072 577690 318132 578000
rect 319160 577690 319220 578000
rect 315760 577630 318132 577690
rect 318934 577630 319220 577690
rect 320384 577690 320444 578000
rect 330040 577690 330100 578000
rect 320384 577630 320466 577690
rect 330040 577630 330218 577690
rect 314518 575245 314578 577630
rect 318014 576870 318074 577630
rect 318934 576870 318994 577630
rect 318014 576810 318994 576870
rect 314515 575244 314581 575245
rect 314515 575180 314516 575244
rect 314580 575180 314581 575244
rect 314515 575179 314581 575180
rect 312954 574038 312986 574274
rect 313222 574038 313306 574274
rect 313542 574038 313574 574274
rect 313779 574292 313845 574293
rect 313779 574228 313780 574292
rect 313844 574228 313845 574292
rect 313779 574227 313845 574228
rect 312954 554274 313574 574038
rect 312954 554038 312986 554274
rect 313222 554038 313306 554274
rect 313542 554038 313574 554274
rect 312954 539308 313574 554038
rect 315514 556954 316134 576000
rect 318934 574157 318994 576810
rect 318931 574156 318997 574157
rect 318931 574092 318932 574156
rect 318996 574092 318997 574156
rect 318931 574091 318997 574092
rect 315514 556718 315546 556954
rect 315782 556718 315866 556954
rect 316102 556718 316134 556954
rect 315514 539308 316134 556718
rect 319234 560614 319854 576000
rect 320406 575381 320466 577630
rect 320403 575380 320469 575381
rect 320403 575316 320404 575380
rect 320468 575316 320469 575380
rect 320403 575315 320469 575316
rect 319234 560378 319266 560614
rect 319502 560378 319586 560614
rect 319822 560378 319854 560614
rect 319234 540614 319854 560378
rect 319234 540378 319266 540614
rect 319502 540378 319586 540614
rect 319822 540378 319854 540614
rect 319234 539308 319854 540378
rect 321794 563294 322414 576000
rect 321794 563058 321826 563294
rect 322062 563058 322146 563294
rect 322382 563058 322414 563294
rect 321794 543294 322414 563058
rect 321794 543058 321826 543294
rect 322062 543058 322146 543294
rect 322382 543058 322414 543294
rect 321794 539308 322414 543058
rect 322954 564274 323574 576000
rect 322954 564038 322986 564274
rect 323222 564038 323306 564274
rect 323542 564038 323574 564274
rect 322954 544274 323574 564038
rect 322954 544038 322986 544274
rect 323222 544038 323306 544274
rect 323542 544038 323574 544274
rect 322954 539308 323574 544038
rect 325514 566954 326134 576000
rect 325514 566718 325546 566954
rect 325782 566718 325866 566954
rect 326102 566718 326134 566954
rect 325514 546954 326134 566718
rect 325514 546718 325546 546954
rect 325782 546718 325866 546954
rect 326102 546718 326134 546954
rect 325514 539308 326134 546718
rect 329234 570614 329854 576000
rect 330158 575381 330218 577630
rect 330155 575380 330221 575381
rect 330155 575316 330156 575380
rect 330220 575316 330221 575380
rect 330155 575315 330221 575316
rect 329234 570378 329266 570614
rect 329502 570378 329586 570614
rect 329822 570378 329854 570614
rect 329234 550614 329854 570378
rect 329234 550378 329266 550614
rect 329502 550378 329586 550614
rect 329822 550378 329854 550614
rect 329234 539308 329854 550378
rect 331794 573294 332414 576000
rect 331794 573058 331826 573294
rect 332062 573058 332146 573294
rect 332382 573058 332414 573294
rect 331794 553294 332414 573058
rect 331794 553058 331826 553294
rect 332062 553058 332146 553294
rect 332382 553058 332414 553294
rect 331794 539308 332414 553058
rect 332954 574274 333574 576000
rect 332954 574038 332986 574274
rect 333222 574038 333306 574274
rect 333542 574038 333574 574274
rect 332954 554274 333574 574038
rect 332954 554038 332986 554274
rect 333222 554038 333306 554274
rect 333542 554038 333574 554274
rect 332954 539308 333574 554038
rect 335514 556954 336134 576000
rect 336963 575380 337029 575381
rect 336963 575316 336964 575380
rect 337028 575316 337029 575380
rect 336963 575315 337029 575316
rect 336779 574156 336845 574157
rect 336779 574092 336780 574156
rect 336844 574092 336845 574156
rect 336779 574091 336845 574092
rect 335514 556718 335546 556954
rect 335782 556718 335866 556954
rect 336102 556718 336134 556954
rect 335514 539308 336134 556718
rect 216814 537510 216932 537570
rect 205720 537202 205780 537510
rect 216872 537202 216932 537510
rect 218096 537510 218162 537570
rect 218096 537202 218156 537510
rect 200272 533294 200620 533456
rect 200272 533058 200328 533294
rect 200564 533058 200620 533294
rect 200272 532896 200620 533058
rect 336000 533294 336348 533456
rect 336000 533058 336056 533294
rect 336292 533058 336348 533294
rect 336000 532896 336348 533058
rect 200952 523294 201300 523456
rect 200952 523058 201008 523294
rect 201244 523058 201300 523294
rect 200952 522896 201300 523058
rect 335320 523294 335668 523456
rect 335320 523058 335376 523294
rect 335612 523058 335668 523294
rect 335320 522896 335668 523058
rect 200272 513294 200620 513456
rect 200272 513058 200328 513294
rect 200564 513058 200620 513294
rect 200272 512896 200620 513058
rect 336000 513294 336348 513456
rect 336000 513058 336056 513294
rect 336292 513058 336348 513294
rect 336000 512896 336348 513058
rect 200952 503294 201300 503456
rect 200952 503058 201008 503294
rect 201244 503058 201300 503294
rect 200952 502896 201300 503058
rect 335320 503294 335668 503456
rect 335320 503058 335376 503294
rect 335612 503058 335668 503294
rect 335320 502896 335668 503058
rect 200272 493294 200620 493456
rect 200272 493058 200328 493294
rect 200564 493058 200620 493294
rect 200272 492896 200620 493058
rect 336000 493294 336348 493456
rect 336000 493058 336056 493294
rect 336292 493058 336348 493294
rect 336000 492896 336348 493058
rect 200952 483294 201300 483456
rect 200952 483058 201008 483294
rect 201244 483058 201300 483294
rect 200952 482896 201300 483058
rect 335320 483294 335668 483456
rect 335320 483058 335376 483294
rect 335612 483058 335668 483294
rect 335320 482896 335668 483058
rect 199515 475284 199581 475285
rect 199515 475220 199516 475284
rect 199580 475220 199581 475284
rect 199515 475219 199581 475220
rect 199331 475012 199397 475013
rect 199331 474948 199332 475012
rect 199396 474948 199397 475012
rect 199331 474947 199397 474948
rect 198963 455700 199029 455701
rect 198963 455636 198964 455700
rect 199028 455636 199029 455700
rect 198963 455635 199029 455636
rect 198779 454068 198845 454069
rect 198779 454004 198780 454068
rect 198844 454004 198845 454068
rect 198779 454003 198845 454004
rect 198782 452029 198842 454003
rect 198966 452301 199026 455635
rect 199334 452981 199394 474947
rect 199518 453117 199578 475219
rect 200272 473294 200620 473456
rect 200272 473058 200328 473294
rect 200564 473058 200620 473294
rect 200272 472896 200620 473058
rect 336000 473294 336348 473456
rect 336000 473058 336056 473294
rect 336292 473058 336348 473294
rect 336000 472896 336348 473058
rect 200952 463294 201300 463456
rect 200952 463058 201008 463294
rect 201244 463058 201300 463294
rect 200952 462896 201300 463058
rect 335320 463294 335668 463456
rect 335320 463058 335376 463294
rect 335612 463058 335668 463294
rect 335320 462896 335668 463058
rect 213200 453250 213260 454106
rect 213336 453661 213396 454106
rect 213333 453660 213399 453661
rect 213333 453596 213334 453660
rect 213398 453596 213399 453660
rect 213333 453595 213399 453596
rect 230608 453250 230668 454106
rect 233192 453250 233252 454106
rect 235640 453250 235700 454106
rect 213200 453190 213378 453250
rect 230608 453190 230674 453250
rect 199515 453116 199581 453117
rect 199515 453052 199516 453116
rect 199580 453052 199581 453116
rect 199515 453051 199581 453052
rect 199331 452980 199397 452981
rect 199331 452916 199332 452980
rect 199396 452916 199397 452980
rect 199331 452915 199397 452916
rect 213318 452437 213378 453190
rect 230614 452573 230674 453190
rect 233190 453190 233252 453250
rect 235582 453190 235700 453250
rect 238088 453250 238148 454106
rect 240672 453250 240732 454106
rect 243120 453250 243180 454106
rect 245568 453250 245628 454106
rect 238088 453190 238218 453250
rect 240672 453190 240794 453250
rect 243120 453190 243186 453250
rect 233190 452573 233250 453190
rect 235582 452573 235642 453190
rect 238158 452573 238218 453190
rect 240734 452573 240794 453190
rect 243126 452573 243186 453190
rect 245518 453190 245628 453250
rect 248016 453250 248076 454106
rect 250600 453250 250660 454106
rect 253048 453250 253108 454106
rect 255632 454040 255692 454106
rect 255632 453980 255698 454040
rect 248016 453190 248154 453250
rect 250600 453190 250730 453250
rect 253048 453190 253122 453250
rect 245518 452573 245578 453190
rect 230611 452572 230677 452573
rect 230611 452508 230612 452572
rect 230676 452508 230677 452572
rect 230611 452507 230677 452508
rect 233187 452572 233253 452573
rect 233187 452508 233188 452572
rect 233252 452508 233253 452572
rect 233187 452507 233253 452508
rect 235579 452572 235645 452573
rect 235579 452508 235580 452572
rect 235644 452508 235645 452572
rect 235579 452507 235645 452508
rect 238155 452572 238221 452573
rect 238155 452508 238156 452572
rect 238220 452508 238221 452572
rect 238155 452507 238221 452508
rect 240731 452572 240797 452573
rect 240731 452508 240732 452572
rect 240796 452508 240797 452572
rect 240731 452507 240797 452508
rect 243123 452572 243189 452573
rect 243123 452508 243124 452572
rect 243188 452508 243189 452572
rect 243123 452507 243189 452508
rect 245515 452572 245581 452573
rect 245515 452508 245516 452572
rect 245580 452508 245581 452572
rect 245515 452507 245581 452508
rect 213315 452436 213381 452437
rect 213315 452372 213316 452436
rect 213380 452372 213381 452436
rect 213315 452371 213381 452372
rect 198963 452300 199029 452301
rect 198963 452236 198964 452300
rect 199028 452236 199029 452300
rect 198963 452235 199029 452236
rect 198779 452028 198845 452029
rect 198779 451964 198780 452028
rect 198844 451964 198845 452028
rect 198779 451963 198845 451964
rect 199234 440614 199854 452000
rect 199234 440378 199266 440614
rect 199502 440378 199586 440614
rect 199822 440378 199854 440614
rect 198779 422924 198845 422925
rect 198779 422860 198780 422924
rect 198844 422860 198845 422924
rect 198779 422859 198845 422860
rect 198595 250476 198661 250477
rect 198595 250412 198596 250476
rect 198660 250412 198661 250476
rect 198595 250411 198661 250412
rect 198782 248029 198842 422859
rect 199234 421162 199854 440378
rect 201794 443294 202414 452000
rect 201794 443058 201826 443294
rect 202062 443058 202146 443294
rect 202382 443058 202414 443294
rect 201794 423294 202414 443058
rect 201794 423058 201826 423294
rect 202062 423058 202146 423294
rect 202382 423058 202414 423294
rect 201794 421162 202414 423058
rect 202954 444274 203574 452000
rect 202954 444038 202986 444274
rect 203222 444038 203306 444274
rect 203542 444038 203574 444274
rect 202954 424274 203574 444038
rect 202954 424038 202986 424274
rect 203222 424038 203306 424274
rect 203542 424038 203574 424274
rect 202954 421162 203574 424038
rect 205514 446954 206134 452000
rect 205514 446718 205546 446954
rect 205782 446718 205866 446954
rect 206102 446718 206134 446954
rect 205514 426954 206134 446718
rect 205514 426718 205546 426954
rect 205782 426718 205866 426954
rect 206102 426718 206134 426954
rect 205514 421162 206134 426718
rect 209234 450614 209854 452000
rect 209234 450378 209266 450614
rect 209502 450378 209586 450614
rect 209822 450378 209854 450614
rect 209234 430614 209854 450378
rect 209234 430378 209266 430614
rect 209502 430378 209586 430614
rect 209822 430378 209854 430614
rect 209234 421162 209854 430378
rect 211794 433294 212414 452000
rect 211794 433058 211826 433294
rect 212062 433058 212146 433294
rect 212382 433058 212414 433294
rect 211794 421162 212414 433058
rect 212954 434274 213574 452000
rect 212954 434038 212986 434274
rect 213222 434038 213306 434274
rect 213542 434038 213574 434274
rect 212954 421162 213574 434038
rect 215514 436954 216134 452000
rect 215514 436718 215546 436954
rect 215782 436718 215866 436954
rect 216102 436718 216134 436954
rect 215514 421162 216134 436718
rect 219234 440614 219854 452000
rect 219234 440378 219266 440614
rect 219502 440378 219586 440614
rect 219822 440378 219854 440614
rect 219234 421162 219854 440378
rect 221794 443294 222414 452000
rect 221794 443058 221826 443294
rect 222062 443058 222146 443294
rect 222382 443058 222414 443294
rect 221794 423294 222414 443058
rect 221794 423058 221826 423294
rect 222062 423058 222146 423294
rect 222382 423058 222414 423294
rect 221794 421162 222414 423058
rect 222954 444274 223574 452000
rect 222954 444038 222986 444274
rect 223222 444038 223306 444274
rect 223542 444038 223574 444274
rect 222954 424274 223574 444038
rect 222954 424038 222986 424274
rect 223222 424038 223306 424274
rect 223542 424038 223574 424274
rect 222954 421162 223574 424038
rect 225514 446954 226134 452000
rect 225514 446718 225546 446954
rect 225782 446718 225866 446954
rect 226102 446718 226134 446954
rect 225514 426954 226134 446718
rect 225514 426718 225546 426954
rect 225782 426718 225866 426954
rect 226102 426718 226134 426954
rect 225514 421162 226134 426718
rect 229234 450614 229854 452000
rect 229234 450378 229266 450614
rect 229502 450378 229586 450614
rect 229822 450378 229854 450614
rect 229234 430614 229854 450378
rect 229234 430378 229266 430614
rect 229502 430378 229586 430614
rect 229822 430378 229854 430614
rect 229234 421162 229854 430378
rect 231794 433294 232414 452000
rect 231794 433058 231826 433294
rect 232062 433058 232146 433294
rect 232382 433058 232414 433294
rect 231794 421162 232414 433058
rect 232954 434274 233574 452000
rect 232954 434038 232986 434274
rect 233222 434038 233306 434274
rect 233542 434038 233574 434274
rect 232954 421162 233574 434038
rect 235514 436954 236134 452000
rect 235514 436718 235546 436954
rect 235782 436718 235866 436954
rect 236102 436718 236134 436954
rect 235514 421162 236134 436718
rect 239234 440614 239854 452000
rect 239234 440378 239266 440614
rect 239502 440378 239586 440614
rect 239822 440378 239854 440614
rect 239234 421162 239854 440378
rect 241794 443294 242414 452000
rect 241794 443058 241826 443294
rect 242062 443058 242146 443294
rect 242382 443058 242414 443294
rect 241794 423294 242414 443058
rect 241794 423058 241826 423294
rect 242062 423058 242146 423294
rect 242382 423058 242414 423294
rect 241794 421162 242414 423058
rect 242954 444274 243574 452000
rect 242954 444038 242986 444274
rect 243222 444038 243306 444274
rect 243542 444038 243574 444274
rect 242954 424274 243574 444038
rect 242954 424038 242986 424274
rect 243222 424038 243306 424274
rect 243542 424038 243574 424274
rect 242954 421162 243574 424038
rect 245514 446954 246134 452000
rect 248094 451349 248154 453190
rect 248091 451348 248157 451349
rect 248091 451284 248092 451348
rect 248156 451284 248157 451348
rect 248091 451283 248157 451284
rect 245514 446718 245546 446954
rect 245782 446718 245866 446954
rect 246102 446718 246134 446954
rect 245514 426954 246134 446718
rect 245514 426718 245546 426954
rect 245782 426718 245866 426954
rect 246102 426718 246134 426954
rect 245514 421162 246134 426718
rect 249234 450614 249854 452000
rect 250670 451349 250730 453190
rect 253062 452573 253122 453190
rect 255638 452573 255698 453980
rect 258080 453250 258140 454106
rect 260664 453250 260724 454106
rect 257846 453190 258140 453250
rect 260606 453190 260724 453250
rect 263112 453250 263172 454106
rect 265560 453250 265620 454106
rect 268280 453250 268340 454106
rect 270592 453250 270652 454106
rect 263112 453190 263242 453250
rect 265560 453190 265634 453250
rect 268280 453190 268394 453250
rect 253059 452572 253125 452573
rect 253059 452508 253060 452572
rect 253124 452508 253125 452572
rect 253059 452507 253125 452508
rect 255635 452572 255701 452573
rect 255635 452508 255636 452572
rect 255700 452508 255701 452572
rect 255635 452507 255701 452508
rect 250667 451348 250733 451349
rect 250667 451284 250668 451348
rect 250732 451284 250733 451348
rect 250667 451283 250733 451284
rect 249234 450378 249266 450614
rect 249502 450378 249586 450614
rect 249822 450378 249854 450614
rect 249234 430614 249854 450378
rect 249234 430378 249266 430614
rect 249502 430378 249586 430614
rect 249822 430378 249854 430614
rect 249234 421162 249854 430378
rect 251794 433294 252414 452000
rect 251794 433058 251826 433294
rect 252062 433058 252146 433294
rect 252382 433058 252414 433294
rect 251794 421162 252414 433058
rect 252954 434274 253574 452000
rect 252954 434038 252986 434274
rect 253222 434038 253306 434274
rect 253542 434038 253574 434274
rect 252954 421162 253574 434038
rect 255514 436954 256134 452000
rect 257846 451346 257906 453190
rect 260606 452573 260666 453190
rect 263182 452573 263242 453190
rect 265574 452573 265634 453190
rect 268334 452573 268394 453190
rect 270542 453190 270652 453250
rect 273040 453250 273100 454106
rect 275624 453250 275684 454106
rect 277392 453250 277452 454106
rect 273040 453190 273178 453250
rect 275624 453190 275754 453250
rect 270542 452573 270602 453190
rect 273118 452573 273178 453190
rect 275694 452573 275754 453190
rect 277166 453190 277452 453250
rect 278072 453250 278132 454106
rect 278480 453250 278540 454106
rect 279568 453250 279628 454106
rect 280520 453250 280580 454106
rect 278072 453190 278146 453250
rect 260603 452572 260669 452573
rect 260603 452508 260604 452572
rect 260668 452508 260669 452572
rect 260603 452507 260669 452508
rect 263179 452572 263245 452573
rect 263179 452508 263180 452572
rect 263244 452508 263245 452572
rect 263179 452507 263245 452508
rect 265571 452572 265637 452573
rect 265571 452508 265572 452572
rect 265636 452508 265637 452572
rect 265571 452507 265637 452508
rect 268331 452572 268397 452573
rect 268331 452508 268332 452572
rect 268396 452508 268397 452572
rect 268331 452507 268397 452508
rect 270539 452572 270605 452573
rect 270539 452508 270540 452572
rect 270604 452508 270605 452572
rect 270539 452507 270605 452508
rect 273115 452572 273181 452573
rect 273115 452508 273116 452572
rect 273180 452508 273181 452572
rect 273115 452507 273181 452508
rect 275691 452572 275757 452573
rect 275691 452508 275692 452572
rect 275756 452508 275757 452572
rect 275691 452507 275757 452508
rect 277166 452165 277226 453190
rect 278086 452573 278146 453190
rect 278454 453190 278540 453250
rect 279558 453190 279628 453250
rect 280478 453190 280580 453250
rect 280792 453250 280852 454106
rect 282152 453250 282212 454106
rect 280792 453190 280906 453250
rect 278083 452572 278149 452573
rect 278083 452508 278084 452572
rect 278148 452508 278149 452572
rect 278083 452507 278149 452508
rect 277163 452164 277229 452165
rect 277163 452100 277164 452164
rect 277228 452100 277229 452164
rect 277163 452099 277229 452100
rect 258027 451348 258093 451349
rect 258027 451346 258028 451348
rect 257846 451286 258028 451346
rect 258027 451284 258028 451286
rect 258092 451284 258093 451348
rect 258027 451283 258093 451284
rect 255514 436718 255546 436954
rect 255782 436718 255866 436954
rect 256102 436718 256134 436954
rect 255514 421162 256134 436718
rect 259234 440614 259854 452000
rect 259234 440378 259266 440614
rect 259502 440378 259586 440614
rect 259822 440378 259854 440614
rect 259234 421162 259854 440378
rect 261794 443294 262414 452000
rect 261794 443058 261826 443294
rect 262062 443058 262146 443294
rect 262382 443058 262414 443294
rect 261794 423294 262414 443058
rect 261794 423058 261826 423294
rect 262062 423058 262146 423294
rect 262382 423058 262414 423294
rect 261794 421162 262414 423058
rect 262954 444274 263574 452000
rect 262954 444038 262986 444274
rect 263222 444038 263306 444274
rect 263542 444038 263574 444274
rect 262954 424274 263574 444038
rect 262954 424038 262986 424274
rect 263222 424038 263306 424274
rect 263542 424038 263574 424274
rect 262954 421162 263574 424038
rect 265514 446954 266134 452000
rect 265514 446718 265546 446954
rect 265782 446718 265866 446954
rect 266102 446718 266134 446954
rect 265514 426954 266134 446718
rect 265514 426718 265546 426954
rect 265782 426718 265866 426954
rect 266102 426718 266134 426954
rect 265514 421162 266134 426718
rect 269234 450614 269854 452000
rect 269234 450378 269266 450614
rect 269502 450378 269586 450614
rect 269822 450378 269854 450614
rect 269234 430614 269854 450378
rect 269234 430378 269266 430614
rect 269502 430378 269586 430614
rect 269822 430378 269854 430614
rect 269234 421162 269854 430378
rect 271794 433294 272414 452000
rect 271794 433058 271826 433294
rect 272062 433058 272146 433294
rect 272382 433058 272414 433294
rect 271794 421162 272414 433058
rect 272954 434274 273574 452000
rect 272954 434038 272986 434274
rect 273222 434038 273306 434274
rect 273542 434038 273574 434274
rect 272954 421162 273574 434038
rect 275514 436954 276134 452000
rect 278454 451893 278514 453190
rect 279558 453117 279618 453190
rect 279555 453116 279621 453117
rect 279555 453052 279556 453116
rect 279620 453052 279621 453116
rect 279555 453051 279621 453052
rect 280478 452573 280538 453190
rect 280475 452572 280541 452573
rect 280475 452508 280476 452572
rect 280540 452508 280541 452572
rect 280475 452507 280541 452508
rect 280846 452301 280906 453190
rect 282134 453190 282212 453250
rect 282968 453250 283028 454106
rect 283240 453250 283300 454106
rect 284328 453661 284388 454106
rect 284325 453660 284391 453661
rect 284325 453596 284326 453660
rect 284390 453596 284391 453660
rect 284325 453595 284391 453596
rect 285416 453250 285476 454106
rect 282968 453190 283114 453250
rect 282134 452573 282194 453190
rect 283054 452573 283114 453190
rect 283238 453190 283300 453250
rect 285262 453190 285476 453250
rect 285552 453250 285612 454106
rect 286776 453661 286836 454106
rect 286773 453660 286839 453661
rect 286773 453596 286774 453660
rect 286838 453596 286839 453660
rect 286773 453595 286839 453596
rect 287864 453522 287924 454106
rect 288272 453522 288332 454106
rect 288952 453797 289012 454106
rect 288949 453796 289015 453797
rect 288949 453732 288950 453796
rect 289014 453732 289015 453796
rect 288949 453731 289015 453732
rect 290176 453661 290236 454106
rect 290173 453660 290239 453661
rect 290173 453596 290174 453660
rect 290238 453596 290239 453660
rect 290173 453595 290239 453596
rect 287838 453462 287924 453522
rect 288206 453462 288332 453522
rect 290584 453522 290644 454106
rect 291264 453661 291324 454106
rect 291261 453660 291327 453661
rect 291261 453596 291262 453660
rect 291326 453596 291327 453660
rect 291261 453595 291327 453596
rect 292624 453522 292684 454106
rect 293032 453522 293092 454106
rect 293712 453661 293772 454106
rect 294800 453797 294860 454106
rect 294797 453796 294863 453797
rect 294797 453732 294798 453796
rect 294862 453732 294863 453796
rect 294797 453731 294863 453732
rect 293709 453660 293775 453661
rect 293709 453596 293710 453660
rect 293774 453596 293775 453660
rect 293709 453595 293775 453596
rect 290584 453462 290658 453522
rect 285552 453190 285690 453250
rect 282131 452572 282197 452573
rect 282131 452508 282132 452572
rect 282196 452508 282197 452572
rect 282131 452507 282197 452508
rect 283051 452572 283117 452573
rect 283051 452508 283052 452572
rect 283116 452508 283117 452572
rect 283051 452507 283117 452508
rect 283238 452301 283298 453190
rect 285262 452981 285322 453190
rect 285259 452980 285325 452981
rect 285259 452916 285260 452980
rect 285324 452916 285325 452980
rect 285259 452915 285325 452916
rect 285630 452573 285690 453190
rect 285627 452572 285693 452573
rect 285627 452508 285628 452572
rect 285692 452508 285693 452572
rect 285627 452507 285693 452508
rect 287838 452301 287898 453462
rect 288206 452573 288266 453462
rect 290598 452573 290658 453462
rect 292622 453462 292684 453522
rect 292990 453462 293092 453522
rect 295480 453522 295540 454106
rect 295888 453522 295948 454106
rect 297112 453661 297172 454106
rect 297109 453660 297175 453661
rect 297109 453596 297110 453660
rect 297174 453596 297175 453660
rect 297109 453595 297175 453596
rect 295480 453462 295626 453522
rect 295888 453462 295994 453522
rect 292622 452573 292682 453462
rect 292990 452573 293050 453462
rect 295566 452573 295626 453462
rect 295934 452845 295994 453462
rect 298064 453250 298124 454106
rect 298472 453661 298532 454106
rect 299560 453661 299620 454106
rect 298469 453660 298535 453661
rect 298469 453596 298470 453660
rect 298534 453596 298535 453660
rect 298469 453595 298535 453596
rect 299557 453660 299623 453661
rect 299557 453596 299558 453660
rect 299622 453596 299623 453660
rect 299557 453595 299623 453596
rect 300512 453250 300572 454106
rect 298064 453190 298202 453250
rect 295931 452844 295997 452845
rect 295931 452780 295932 452844
rect 295996 452780 295997 452844
rect 295931 452779 295997 452780
rect 298142 452573 298202 453190
rect 300350 453190 300572 453250
rect 300648 453250 300708 454106
rect 302008 453250 302068 454106
rect 302960 453250 303020 454106
rect 300648 453190 300778 453250
rect 300350 452573 300410 453190
rect 288203 452572 288269 452573
rect 288203 452508 288204 452572
rect 288268 452508 288269 452572
rect 288203 452507 288269 452508
rect 290595 452572 290661 452573
rect 290595 452508 290596 452572
rect 290660 452508 290661 452572
rect 290595 452507 290661 452508
rect 292619 452572 292685 452573
rect 292619 452508 292620 452572
rect 292684 452508 292685 452572
rect 292619 452507 292685 452508
rect 292987 452572 293053 452573
rect 292987 452508 292988 452572
rect 293052 452508 293053 452572
rect 292987 452507 293053 452508
rect 295563 452572 295629 452573
rect 295563 452508 295564 452572
rect 295628 452508 295629 452572
rect 295563 452507 295629 452508
rect 298139 452572 298205 452573
rect 298139 452508 298140 452572
rect 298204 452508 298205 452572
rect 298139 452507 298205 452508
rect 300347 452572 300413 452573
rect 300347 452508 300348 452572
rect 300412 452508 300413 452572
rect 300347 452507 300413 452508
rect 300718 452301 300778 453190
rect 302006 453190 302068 453250
rect 302926 453190 303020 453250
rect 303096 453250 303156 454106
rect 304184 453250 304244 454106
rect 305272 453250 305332 454106
rect 305816 453250 305876 454106
rect 306496 453250 306556 454106
rect 303096 453190 303170 453250
rect 304184 453190 304274 453250
rect 305272 453190 305378 453250
rect 305816 453190 305930 453250
rect 302006 452573 302066 453190
rect 302003 452572 302069 452573
rect 302003 452508 302004 452572
rect 302068 452508 302069 452572
rect 302003 452507 302069 452508
rect 302926 452301 302986 453190
rect 303110 452573 303170 453190
rect 304214 452573 304274 453190
rect 305318 452573 305378 453190
rect 303107 452572 303173 452573
rect 303107 452508 303108 452572
rect 303172 452508 303173 452572
rect 303107 452507 303173 452508
rect 304211 452572 304277 452573
rect 304211 452508 304212 452572
rect 304276 452508 304277 452572
rect 304211 452507 304277 452508
rect 305315 452572 305381 452573
rect 305315 452508 305316 452572
rect 305380 452508 305381 452572
rect 305315 452507 305381 452508
rect 305870 452301 305930 453190
rect 306422 453190 306556 453250
rect 307856 453250 307916 454106
rect 308264 453250 308324 454106
rect 307856 453190 307954 453250
rect 306422 452573 306482 453190
rect 307894 452573 307954 453190
rect 308262 453190 308324 453250
rect 308944 453250 309004 454106
rect 310032 453250 310092 454106
rect 311120 453661 311180 454106
rect 312344 453661 312404 454106
rect 311117 453660 311183 453661
rect 311117 453596 311118 453660
rect 311182 453596 311183 453660
rect 311117 453595 311183 453596
rect 312341 453660 312407 453661
rect 312341 453596 312342 453660
rect 312406 453596 312407 453660
rect 312341 453595 312407 453596
rect 313432 453250 313492 454106
rect 314792 453250 314852 454106
rect 316016 453250 316076 454106
rect 316968 453250 317028 454106
rect 308944 453190 309058 453250
rect 306419 452572 306485 452573
rect 306419 452508 306420 452572
rect 306484 452508 306485 452572
rect 306419 452507 306485 452508
rect 307891 452572 307957 452573
rect 307891 452508 307892 452572
rect 307956 452508 307957 452572
rect 307891 452507 307957 452508
rect 280843 452300 280909 452301
rect 280843 452236 280844 452300
rect 280908 452236 280909 452300
rect 280843 452235 280909 452236
rect 283235 452300 283301 452301
rect 283235 452236 283236 452300
rect 283300 452236 283301 452300
rect 283235 452235 283301 452236
rect 287835 452300 287901 452301
rect 287835 452236 287836 452300
rect 287900 452236 287901 452300
rect 287835 452235 287901 452236
rect 300715 452300 300781 452301
rect 300715 452236 300716 452300
rect 300780 452236 300781 452300
rect 300715 452235 300781 452236
rect 302923 452300 302989 452301
rect 302923 452236 302924 452300
rect 302988 452236 302989 452300
rect 302923 452235 302989 452236
rect 305867 452300 305933 452301
rect 305867 452236 305868 452300
rect 305932 452236 305933 452300
rect 305867 452235 305933 452236
rect 278451 451892 278517 451893
rect 278451 451828 278452 451892
rect 278516 451828 278517 451892
rect 278451 451827 278517 451828
rect 275514 436718 275546 436954
rect 275782 436718 275866 436954
rect 276102 436718 276134 436954
rect 275514 421162 276134 436718
rect 279234 440614 279854 452000
rect 279234 440378 279266 440614
rect 279502 440378 279586 440614
rect 279822 440378 279854 440614
rect 279234 421162 279854 440378
rect 281794 443294 282414 452000
rect 281794 443058 281826 443294
rect 282062 443058 282146 443294
rect 282382 443058 282414 443294
rect 281794 423294 282414 443058
rect 281794 423058 281826 423294
rect 282062 423058 282146 423294
rect 282382 423058 282414 423294
rect 281794 421162 282414 423058
rect 282954 444274 283574 452000
rect 282954 444038 282986 444274
rect 283222 444038 283306 444274
rect 283542 444038 283574 444274
rect 282954 424274 283574 444038
rect 282954 424038 282986 424274
rect 283222 424038 283306 424274
rect 283542 424038 283574 424274
rect 282954 421162 283574 424038
rect 285514 446954 286134 452000
rect 285514 446718 285546 446954
rect 285782 446718 285866 446954
rect 286102 446718 286134 446954
rect 285514 426954 286134 446718
rect 285514 426718 285546 426954
rect 285782 426718 285866 426954
rect 286102 426718 286134 426954
rect 285514 421162 286134 426718
rect 289234 450614 289854 452000
rect 289234 450378 289266 450614
rect 289502 450378 289586 450614
rect 289822 450378 289854 450614
rect 289234 430614 289854 450378
rect 289234 430378 289266 430614
rect 289502 430378 289586 430614
rect 289822 430378 289854 430614
rect 289234 421162 289854 430378
rect 291794 433294 292414 452000
rect 291794 433058 291826 433294
rect 292062 433058 292146 433294
rect 292382 433058 292414 433294
rect 291794 421162 292414 433058
rect 292954 434274 293574 452000
rect 292954 434038 292986 434274
rect 293222 434038 293306 434274
rect 293542 434038 293574 434274
rect 292954 421162 293574 434038
rect 295514 436954 296134 452000
rect 295514 436718 295546 436954
rect 295782 436718 295866 436954
rect 296102 436718 296134 436954
rect 295514 421162 296134 436718
rect 299234 440614 299854 452000
rect 299234 440378 299266 440614
rect 299502 440378 299586 440614
rect 299822 440378 299854 440614
rect 299234 421162 299854 440378
rect 301794 443294 302414 452000
rect 301794 443058 301826 443294
rect 302062 443058 302146 443294
rect 302382 443058 302414 443294
rect 301794 423294 302414 443058
rect 301794 423058 301826 423294
rect 302062 423058 302146 423294
rect 302382 423058 302414 423294
rect 301794 421162 302414 423058
rect 302954 444274 303574 452000
rect 302954 444038 302986 444274
rect 303222 444038 303306 444274
rect 303542 444038 303574 444274
rect 302954 424274 303574 444038
rect 302954 424038 302986 424274
rect 303222 424038 303306 424274
rect 303542 424038 303574 424274
rect 302954 421162 303574 424038
rect 305514 446954 306134 452000
rect 308262 451349 308322 453190
rect 308998 452573 309058 453190
rect 309918 453190 310092 453250
rect 313414 453190 313492 453250
rect 314702 453190 314852 453250
rect 315990 453190 316076 453250
rect 316910 453190 317028 453250
rect 318328 453250 318388 454106
rect 319416 453250 319476 454106
rect 320504 453250 320564 454106
rect 318328 453190 318442 453250
rect 319416 453190 319546 453250
rect 309918 452573 309978 453190
rect 313414 452573 313474 453190
rect 314702 452573 314762 453190
rect 315990 452573 316050 453190
rect 316910 452573 316970 453190
rect 318382 452573 318442 453190
rect 308995 452572 309061 452573
rect 308995 452508 308996 452572
rect 309060 452508 309061 452572
rect 308995 452507 309061 452508
rect 309915 452572 309981 452573
rect 309915 452508 309916 452572
rect 309980 452508 309981 452572
rect 309915 452507 309981 452508
rect 313411 452572 313477 452573
rect 313411 452508 313412 452572
rect 313476 452508 313477 452572
rect 313411 452507 313477 452508
rect 314699 452572 314765 452573
rect 314699 452508 314700 452572
rect 314764 452508 314765 452572
rect 314699 452507 314765 452508
rect 315987 452572 316053 452573
rect 315987 452508 315988 452572
rect 316052 452508 316053 452572
rect 315987 452507 316053 452508
rect 316907 452572 316973 452573
rect 316907 452508 316908 452572
rect 316972 452508 316973 452572
rect 316907 452507 316973 452508
rect 318379 452572 318445 452573
rect 318379 452508 318380 452572
rect 318444 452508 318445 452572
rect 318379 452507 318445 452508
rect 319486 452301 319546 453190
rect 320406 453190 320564 453250
rect 320406 452573 320466 453190
rect 320403 452572 320469 452573
rect 320403 452508 320404 452572
rect 320468 452508 320469 452572
rect 320403 452507 320469 452508
rect 319483 452300 319549 452301
rect 319483 452236 319484 452300
rect 319548 452236 319549 452300
rect 319483 452235 319549 452236
rect 308259 451348 308325 451349
rect 308259 451284 308260 451348
rect 308324 451284 308325 451348
rect 308259 451283 308325 451284
rect 305514 446718 305546 446954
rect 305782 446718 305866 446954
rect 306102 446718 306134 446954
rect 305514 426954 306134 446718
rect 305514 426718 305546 426954
rect 305782 426718 305866 426954
rect 306102 426718 306134 426954
rect 305514 421162 306134 426718
rect 309234 450614 309854 452000
rect 309234 450378 309266 450614
rect 309502 450378 309586 450614
rect 309822 450378 309854 450614
rect 309234 430614 309854 450378
rect 309234 430378 309266 430614
rect 309502 430378 309586 430614
rect 309822 430378 309854 430614
rect 309234 421162 309854 430378
rect 311794 433294 312414 452000
rect 311794 433058 311826 433294
rect 312062 433058 312146 433294
rect 312382 433058 312414 433294
rect 311794 421162 312414 433058
rect 312954 434274 313574 452000
rect 312954 434038 312986 434274
rect 313222 434038 313306 434274
rect 313542 434038 313574 434274
rect 312954 421162 313574 434038
rect 315514 436954 316134 452000
rect 315514 436718 315546 436954
rect 315782 436718 315866 436954
rect 316102 436718 316134 436954
rect 315514 421162 316134 436718
rect 319234 440614 319854 452000
rect 319234 440378 319266 440614
rect 319502 440378 319586 440614
rect 319822 440378 319854 440614
rect 319234 421162 319854 440378
rect 321794 443294 322414 452000
rect 321794 443058 321826 443294
rect 322062 443058 322146 443294
rect 322382 443058 322414 443294
rect 321794 423294 322414 443058
rect 321794 423058 321826 423294
rect 322062 423058 322146 423294
rect 322382 423058 322414 423294
rect 321794 421162 322414 423058
rect 322954 444274 323574 452000
rect 322954 444038 322986 444274
rect 323222 444038 323306 444274
rect 323542 444038 323574 444274
rect 322954 424274 323574 444038
rect 322954 424038 322986 424274
rect 323222 424038 323306 424274
rect 323542 424038 323574 424274
rect 322954 421162 323574 424038
rect 325514 446954 326134 452000
rect 325514 446718 325546 446954
rect 325782 446718 325866 446954
rect 326102 446718 326134 446954
rect 325514 426954 326134 446718
rect 325514 426718 325546 426954
rect 325782 426718 325866 426954
rect 326102 426718 326134 426954
rect 325514 421162 326134 426718
rect 329234 450614 329854 452000
rect 329234 450378 329266 450614
rect 329502 450378 329586 450614
rect 329822 450378 329854 450614
rect 329234 430614 329854 450378
rect 329234 430378 329266 430614
rect 329502 430378 329586 430614
rect 329822 430378 329854 430614
rect 329234 421162 329854 430378
rect 331794 433294 332414 452000
rect 331794 433058 331826 433294
rect 332062 433058 332146 433294
rect 332382 433058 332414 433294
rect 331794 421162 332414 433058
rect 332954 434274 333574 452000
rect 332954 434038 332986 434274
rect 333222 434038 333306 434274
rect 333542 434038 333574 434274
rect 332954 421162 333574 434038
rect 335514 436954 336134 452000
rect 336782 447677 336842 574091
rect 336966 447813 337026 575315
rect 337147 543012 337213 543013
rect 337147 542948 337148 543012
rect 337212 542948 337213 543012
rect 337147 542947 337213 542948
rect 336963 447812 337029 447813
rect 336963 447748 336964 447812
rect 337028 447748 337029 447812
rect 336963 447747 337029 447748
rect 336779 447676 336845 447677
rect 336779 447612 336780 447676
rect 336844 447612 336845 447676
rect 336779 447611 336845 447612
rect 335514 436718 335546 436954
rect 335782 436718 335866 436954
rect 336102 436718 336134 436954
rect 335514 421162 336134 436718
rect 337150 421837 337210 542947
rect 338070 439517 338130 610947
rect 338254 447949 338314 612171
rect 339234 600614 339854 620378
rect 339234 600378 339266 600614
rect 339502 600378 339586 600614
rect 339822 600378 339854 600614
rect 339234 580614 339854 600378
rect 339234 580378 339266 580614
rect 339502 580378 339586 580614
rect 339822 580378 339854 580614
rect 339234 560614 339854 580378
rect 339234 560378 339266 560614
rect 339502 560378 339586 560614
rect 339822 560378 339854 560614
rect 338987 543012 339053 543013
rect 338987 542948 338988 543012
rect 339052 542948 339053 543012
rect 338987 542947 339053 542948
rect 338435 462092 338501 462093
rect 338435 462028 338436 462092
rect 338500 462028 338501 462092
rect 338435 462027 338501 462028
rect 338438 461549 338498 462027
rect 338435 461548 338501 461549
rect 338435 461484 338436 461548
rect 338500 461484 338501 461548
rect 338435 461483 338501 461484
rect 338251 447948 338317 447949
rect 338251 447884 338252 447948
rect 338316 447884 338317 447948
rect 338251 447883 338317 447884
rect 338067 439516 338133 439517
rect 338067 439452 338068 439516
rect 338132 439452 338133 439516
rect 338067 439451 338133 439452
rect 338438 425781 338498 461483
rect 338435 425780 338501 425781
rect 338435 425716 338436 425780
rect 338500 425716 338501 425780
rect 338435 425715 338501 425716
rect 338990 421837 339050 542947
rect 339234 540614 339854 560378
rect 339234 540378 339266 540614
rect 339502 540378 339586 540614
rect 339822 540378 339854 540614
rect 339234 520614 339854 540378
rect 339234 520378 339266 520614
rect 339502 520378 339586 520614
rect 339822 520378 339854 520614
rect 339234 500614 339854 520378
rect 339234 500378 339266 500614
rect 339502 500378 339586 500614
rect 339822 500378 339854 500614
rect 339234 480614 339854 500378
rect 339234 480378 339266 480614
rect 339502 480378 339586 480614
rect 339822 480378 339854 480614
rect 339234 460614 339854 480378
rect 339234 460378 339266 460614
rect 339502 460378 339586 460614
rect 339822 460378 339854 460614
rect 339234 440614 339854 460378
rect 339234 440378 339266 440614
rect 339502 440378 339586 440614
rect 339822 440378 339854 440614
rect 337147 421836 337213 421837
rect 337147 421772 337148 421836
rect 337212 421772 337213 421836
rect 337147 421771 337213 421772
rect 338987 421836 339053 421837
rect 338987 421772 338988 421836
rect 339052 421772 339053 421836
rect 338987 421771 339053 421772
rect 339234 421162 339854 440378
rect 340094 421837 340154 659635
rect 341794 643294 342414 663058
rect 341794 643058 341826 643294
rect 342062 643058 342146 643294
rect 342382 643058 342414 643294
rect 341794 623294 342414 643058
rect 341794 623058 341826 623294
rect 342062 623058 342146 623294
rect 342382 623058 342414 623294
rect 341794 603294 342414 623058
rect 341794 603058 341826 603294
rect 342062 603058 342146 603294
rect 342382 603058 342414 603294
rect 341794 583294 342414 603058
rect 341794 583058 341826 583294
rect 342062 583058 342146 583294
rect 342382 583058 342414 583294
rect 341563 576060 341629 576061
rect 341563 575996 341564 576060
rect 341628 575996 341629 576060
rect 341563 575995 341629 575996
rect 341566 543149 341626 575995
rect 341794 563294 342414 583058
rect 341794 563058 341826 563294
rect 342062 563058 342146 563294
rect 342382 563058 342414 563294
rect 341794 543294 342414 563058
rect 341563 543148 341629 543149
rect 341563 543084 341564 543148
rect 341628 543084 341629 543148
rect 341563 543083 341629 543084
rect 341566 428093 341626 543083
rect 341794 543058 341826 543294
rect 342062 543058 342146 543294
rect 342382 543058 342414 543294
rect 341794 523294 342414 543058
rect 341794 523058 341826 523294
rect 342062 523058 342146 523294
rect 342382 523058 342414 523294
rect 341794 503294 342414 523058
rect 341794 503058 341826 503294
rect 342062 503058 342146 503294
rect 342382 503058 342414 503294
rect 341794 483294 342414 503058
rect 341794 483058 341826 483294
rect 342062 483058 342146 483294
rect 342382 483058 342414 483294
rect 341794 463294 342414 483058
rect 341794 463058 341826 463294
rect 342062 463058 342146 463294
rect 342382 463058 342414 463294
rect 341794 443294 342414 463058
rect 341794 443058 341826 443294
rect 342062 443058 342146 443294
rect 342382 443058 342414 443294
rect 341563 428092 341629 428093
rect 341563 428028 341564 428092
rect 341628 428028 341629 428092
rect 341563 428027 341629 428028
rect 341794 423294 342414 443058
rect 341794 423058 341826 423294
rect 342062 423058 342146 423294
rect 342382 423058 342414 423294
rect 340091 421836 340157 421837
rect 340091 421772 340092 421836
rect 340156 421772 340157 421836
rect 340091 421771 340157 421772
rect 341794 421162 342414 423058
rect 342954 684274 343574 711002
rect 352954 710598 353574 711590
rect 352954 710362 352986 710598
rect 353222 710362 353306 710598
rect 353542 710362 353574 710598
rect 352954 710278 353574 710362
rect 352954 710042 352986 710278
rect 353222 710042 353306 710278
rect 353542 710042 353574 710278
rect 349234 708678 349854 709670
rect 349234 708442 349266 708678
rect 349502 708442 349586 708678
rect 349822 708442 349854 708678
rect 349234 708358 349854 708442
rect 349234 708122 349266 708358
rect 349502 708122 349586 708358
rect 349822 708122 349854 708358
rect 342954 684038 342986 684274
rect 343222 684038 343306 684274
rect 343542 684038 343574 684274
rect 342954 664274 343574 684038
rect 342954 664038 342986 664274
rect 343222 664038 343306 664274
rect 343542 664038 343574 664274
rect 342954 644274 343574 664038
rect 342954 644038 342986 644274
rect 343222 644038 343306 644274
rect 343542 644038 343574 644274
rect 342954 624274 343574 644038
rect 342954 624038 342986 624274
rect 343222 624038 343306 624274
rect 343542 624038 343574 624274
rect 342954 604274 343574 624038
rect 342954 604038 342986 604274
rect 343222 604038 343306 604274
rect 343542 604038 343574 604274
rect 342954 584274 343574 604038
rect 342954 584038 342986 584274
rect 343222 584038 343306 584274
rect 343542 584038 343574 584274
rect 342954 564274 343574 584038
rect 342954 564038 342986 564274
rect 343222 564038 343306 564274
rect 343542 564038 343574 564274
rect 342954 544274 343574 564038
rect 342954 544038 342986 544274
rect 343222 544038 343306 544274
rect 343542 544038 343574 544274
rect 342954 524274 343574 544038
rect 342954 524038 342986 524274
rect 343222 524038 343306 524274
rect 343542 524038 343574 524274
rect 342954 504274 343574 524038
rect 342954 504038 342986 504274
rect 343222 504038 343306 504274
rect 343542 504038 343574 504274
rect 342954 484274 343574 504038
rect 342954 484038 342986 484274
rect 343222 484038 343306 484274
rect 343542 484038 343574 484274
rect 342954 464274 343574 484038
rect 342954 464038 342986 464274
rect 343222 464038 343306 464274
rect 343542 464038 343574 464274
rect 342954 444274 343574 464038
rect 342954 444038 342986 444274
rect 343222 444038 343306 444274
rect 343542 444038 343574 444274
rect 342954 424274 343574 444038
rect 342954 424038 342986 424274
rect 343222 424038 343306 424274
rect 343542 424038 343574 424274
rect 342954 421162 343574 424038
rect 345514 706758 346134 707750
rect 345514 706522 345546 706758
rect 345782 706522 345866 706758
rect 346102 706522 346134 706758
rect 345514 706438 346134 706522
rect 345514 706202 345546 706438
rect 345782 706202 345866 706438
rect 346102 706202 346134 706438
rect 345514 686954 346134 706202
rect 345514 686718 345546 686954
rect 345782 686718 345866 686954
rect 346102 686718 346134 686954
rect 345514 666954 346134 686718
rect 345514 666718 345546 666954
rect 345782 666718 345866 666954
rect 346102 666718 346134 666954
rect 345514 646954 346134 666718
rect 345514 646718 345546 646954
rect 345782 646718 345866 646954
rect 346102 646718 346134 646954
rect 345514 626954 346134 646718
rect 345514 626718 345546 626954
rect 345782 626718 345866 626954
rect 346102 626718 346134 626954
rect 345514 606954 346134 626718
rect 345514 606718 345546 606954
rect 345782 606718 345866 606954
rect 346102 606718 346134 606954
rect 345514 586954 346134 606718
rect 345514 586718 345546 586954
rect 345782 586718 345866 586954
rect 346102 586718 346134 586954
rect 345514 566954 346134 586718
rect 345514 566718 345546 566954
rect 345782 566718 345866 566954
rect 346102 566718 346134 566954
rect 345514 546954 346134 566718
rect 345514 546718 345546 546954
rect 345782 546718 345866 546954
rect 346102 546718 346134 546954
rect 345514 526954 346134 546718
rect 345514 526718 345546 526954
rect 345782 526718 345866 526954
rect 346102 526718 346134 526954
rect 345514 506954 346134 526718
rect 345514 506718 345546 506954
rect 345782 506718 345866 506954
rect 346102 506718 346134 506954
rect 345514 486954 346134 506718
rect 345514 486718 345546 486954
rect 345782 486718 345866 486954
rect 346102 486718 346134 486954
rect 345514 466954 346134 486718
rect 345514 466718 345546 466954
rect 345782 466718 345866 466954
rect 346102 466718 346134 466954
rect 345514 446954 346134 466718
rect 345514 446718 345546 446954
rect 345782 446718 345866 446954
rect 346102 446718 346134 446954
rect 345514 426954 346134 446718
rect 345514 426718 345546 426954
rect 345782 426718 345866 426954
rect 346102 426718 346134 426954
rect 345514 421162 346134 426718
rect 349234 690614 349854 708122
rect 349234 690378 349266 690614
rect 349502 690378 349586 690614
rect 349822 690378 349854 690614
rect 349234 670614 349854 690378
rect 349234 670378 349266 670614
rect 349502 670378 349586 670614
rect 349822 670378 349854 670614
rect 349234 650614 349854 670378
rect 349234 650378 349266 650614
rect 349502 650378 349586 650614
rect 349822 650378 349854 650614
rect 349234 630614 349854 650378
rect 349234 630378 349266 630614
rect 349502 630378 349586 630614
rect 349822 630378 349854 630614
rect 349234 610614 349854 630378
rect 349234 610378 349266 610614
rect 349502 610378 349586 610614
rect 349822 610378 349854 610614
rect 349234 590614 349854 610378
rect 349234 590378 349266 590614
rect 349502 590378 349586 590614
rect 349822 590378 349854 590614
rect 349234 570614 349854 590378
rect 349234 570378 349266 570614
rect 349502 570378 349586 570614
rect 349822 570378 349854 570614
rect 349234 550614 349854 570378
rect 349234 550378 349266 550614
rect 349502 550378 349586 550614
rect 349822 550378 349854 550614
rect 349234 530614 349854 550378
rect 349234 530378 349266 530614
rect 349502 530378 349586 530614
rect 349822 530378 349854 530614
rect 349234 510614 349854 530378
rect 349234 510378 349266 510614
rect 349502 510378 349586 510614
rect 349822 510378 349854 510614
rect 349234 490614 349854 510378
rect 349234 490378 349266 490614
rect 349502 490378 349586 490614
rect 349822 490378 349854 490614
rect 349234 470614 349854 490378
rect 349234 470378 349266 470614
rect 349502 470378 349586 470614
rect 349822 470378 349854 470614
rect 349234 450614 349854 470378
rect 349234 450378 349266 450614
rect 349502 450378 349586 450614
rect 349822 450378 349854 450614
rect 349234 430614 349854 450378
rect 349234 430378 349266 430614
rect 349502 430378 349586 430614
rect 349822 430378 349854 430614
rect 349234 421162 349854 430378
rect 351794 705798 352414 705830
rect 351794 705562 351826 705798
rect 352062 705562 352146 705798
rect 352382 705562 352414 705798
rect 351794 705478 352414 705562
rect 351794 705242 351826 705478
rect 352062 705242 352146 705478
rect 352382 705242 352414 705478
rect 351794 693294 352414 705242
rect 351794 693058 351826 693294
rect 352062 693058 352146 693294
rect 352382 693058 352414 693294
rect 351794 673294 352414 693058
rect 351794 673058 351826 673294
rect 352062 673058 352146 673294
rect 352382 673058 352414 673294
rect 351794 653294 352414 673058
rect 351794 653058 351826 653294
rect 352062 653058 352146 653294
rect 352382 653058 352414 653294
rect 351794 633294 352414 653058
rect 351794 633058 351826 633294
rect 352062 633058 352146 633294
rect 352382 633058 352414 633294
rect 351794 613294 352414 633058
rect 351794 613058 351826 613294
rect 352062 613058 352146 613294
rect 352382 613058 352414 613294
rect 351794 593294 352414 613058
rect 351794 593058 351826 593294
rect 352062 593058 352146 593294
rect 352382 593058 352414 593294
rect 351794 573294 352414 593058
rect 351794 573058 351826 573294
rect 352062 573058 352146 573294
rect 352382 573058 352414 573294
rect 351794 553294 352414 573058
rect 351794 553058 351826 553294
rect 352062 553058 352146 553294
rect 352382 553058 352414 553294
rect 351794 533294 352414 553058
rect 351794 533058 351826 533294
rect 352062 533058 352146 533294
rect 352382 533058 352414 533294
rect 351794 513294 352414 533058
rect 351794 513058 351826 513294
rect 352062 513058 352146 513294
rect 352382 513058 352414 513294
rect 351794 493294 352414 513058
rect 351794 493058 351826 493294
rect 352062 493058 352146 493294
rect 352382 493058 352414 493294
rect 351794 473294 352414 493058
rect 351794 473058 351826 473294
rect 352062 473058 352146 473294
rect 352382 473058 352414 473294
rect 351794 453294 352414 473058
rect 351794 453058 351826 453294
rect 352062 453058 352146 453294
rect 352382 453058 352414 453294
rect 351794 433294 352414 453058
rect 351794 433058 351826 433294
rect 352062 433058 352146 433294
rect 352382 433058 352414 433294
rect 351794 421162 352414 433058
rect 352954 694274 353574 710042
rect 362954 711558 363574 711590
rect 362954 711322 362986 711558
rect 363222 711322 363306 711558
rect 363542 711322 363574 711558
rect 362954 711238 363574 711322
rect 362954 711002 362986 711238
rect 363222 711002 363306 711238
rect 363542 711002 363574 711238
rect 359234 709638 359854 709670
rect 359234 709402 359266 709638
rect 359502 709402 359586 709638
rect 359822 709402 359854 709638
rect 359234 709318 359854 709402
rect 359234 709082 359266 709318
rect 359502 709082 359586 709318
rect 359822 709082 359854 709318
rect 352954 694038 352986 694274
rect 353222 694038 353306 694274
rect 353542 694038 353574 694274
rect 352954 674274 353574 694038
rect 352954 674038 352986 674274
rect 353222 674038 353306 674274
rect 353542 674038 353574 674274
rect 352954 654274 353574 674038
rect 352954 654038 352986 654274
rect 353222 654038 353306 654274
rect 353542 654038 353574 654274
rect 352954 634274 353574 654038
rect 352954 634038 352986 634274
rect 353222 634038 353306 634274
rect 353542 634038 353574 634274
rect 352954 614274 353574 634038
rect 352954 614038 352986 614274
rect 353222 614038 353306 614274
rect 353542 614038 353574 614274
rect 352954 594274 353574 614038
rect 352954 594038 352986 594274
rect 353222 594038 353306 594274
rect 353542 594038 353574 594274
rect 352954 574274 353574 594038
rect 352954 574038 352986 574274
rect 353222 574038 353306 574274
rect 353542 574038 353574 574274
rect 352954 554274 353574 574038
rect 352954 554038 352986 554274
rect 353222 554038 353306 554274
rect 353542 554038 353574 554274
rect 352954 534274 353574 554038
rect 352954 534038 352986 534274
rect 353222 534038 353306 534274
rect 353542 534038 353574 534274
rect 352954 514274 353574 534038
rect 352954 514038 352986 514274
rect 353222 514038 353306 514274
rect 353542 514038 353574 514274
rect 352954 494274 353574 514038
rect 352954 494038 352986 494274
rect 353222 494038 353306 494274
rect 353542 494038 353574 494274
rect 352954 474274 353574 494038
rect 352954 474038 352986 474274
rect 353222 474038 353306 474274
rect 353542 474038 353574 474274
rect 352954 454274 353574 474038
rect 352954 454038 352986 454274
rect 353222 454038 353306 454274
rect 353542 454038 353574 454274
rect 352954 434274 353574 454038
rect 352954 434038 352986 434274
rect 353222 434038 353306 434274
rect 353542 434038 353574 434274
rect 352954 421162 353574 434038
rect 355514 707718 356134 707750
rect 355514 707482 355546 707718
rect 355782 707482 355866 707718
rect 356102 707482 356134 707718
rect 355514 707398 356134 707482
rect 355514 707162 355546 707398
rect 355782 707162 355866 707398
rect 356102 707162 356134 707398
rect 355514 696954 356134 707162
rect 355514 696718 355546 696954
rect 355782 696718 355866 696954
rect 356102 696718 356134 696954
rect 355514 676954 356134 696718
rect 355514 676718 355546 676954
rect 355782 676718 355866 676954
rect 356102 676718 356134 676954
rect 355514 656954 356134 676718
rect 355514 656718 355546 656954
rect 355782 656718 355866 656954
rect 356102 656718 356134 656954
rect 355514 636954 356134 656718
rect 355514 636718 355546 636954
rect 355782 636718 355866 636954
rect 356102 636718 356134 636954
rect 355514 616954 356134 636718
rect 355514 616718 355546 616954
rect 355782 616718 355866 616954
rect 356102 616718 356134 616954
rect 355514 596954 356134 616718
rect 355514 596718 355546 596954
rect 355782 596718 355866 596954
rect 356102 596718 356134 596954
rect 355514 576954 356134 596718
rect 355514 576718 355546 576954
rect 355782 576718 355866 576954
rect 356102 576718 356134 576954
rect 355514 556954 356134 576718
rect 355514 556718 355546 556954
rect 355782 556718 355866 556954
rect 356102 556718 356134 556954
rect 355514 536954 356134 556718
rect 355514 536718 355546 536954
rect 355782 536718 355866 536954
rect 356102 536718 356134 536954
rect 355514 516954 356134 536718
rect 355514 516718 355546 516954
rect 355782 516718 355866 516954
rect 356102 516718 356134 516954
rect 355514 496954 356134 516718
rect 355514 496718 355546 496954
rect 355782 496718 355866 496954
rect 356102 496718 356134 496954
rect 355514 476954 356134 496718
rect 355514 476718 355546 476954
rect 355782 476718 355866 476954
rect 356102 476718 356134 476954
rect 355514 456954 356134 476718
rect 355514 456718 355546 456954
rect 355782 456718 355866 456954
rect 356102 456718 356134 456954
rect 355514 436954 356134 456718
rect 355514 436718 355546 436954
rect 355782 436718 355866 436954
rect 356102 436718 356134 436954
rect 355514 421162 356134 436718
rect 359234 700614 359854 709082
rect 359234 700378 359266 700614
rect 359502 700378 359586 700614
rect 359822 700378 359854 700614
rect 359234 680614 359854 700378
rect 359234 680378 359266 680614
rect 359502 680378 359586 680614
rect 359822 680378 359854 680614
rect 359234 660614 359854 680378
rect 359234 660378 359266 660614
rect 359502 660378 359586 660614
rect 359822 660378 359854 660614
rect 359234 640614 359854 660378
rect 359234 640378 359266 640614
rect 359502 640378 359586 640614
rect 359822 640378 359854 640614
rect 359234 620614 359854 640378
rect 359234 620378 359266 620614
rect 359502 620378 359586 620614
rect 359822 620378 359854 620614
rect 359234 600614 359854 620378
rect 359234 600378 359266 600614
rect 359502 600378 359586 600614
rect 359822 600378 359854 600614
rect 359234 580614 359854 600378
rect 359234 580378 359266 580614
rect 359502 580378 359586 580614
rect 359822 580378 359854 580614
rect 359234 560614 359854 580378
rect 359234 560378 359266 560614
rect 359502 560378 359586 560614
rect 359822 560378 359854 560614
rect 359234 540614 359854 560378
rect 359234 540378 359266 540614
rect 359502 540378 359586 540614
rect 359822 540378 359854 540614
rect 359234 520614 359854 540378
rect 359234 520378 359266 520614
rect 359502 520378 359586 520614
rect 359822 520378 359854 520614
rect 359234 500614 359854 520378
rect 359234 500378 359266 500614
rect 359502 500378 359586 500614
rect 359822 500378 359854 500614
rect 359234 480614 359854 500378
rect 359234 480378 359266 480614
rect 359502 480378 359586 480614
rect 359822 480378 359854 480614
rect 359234 460614 359854 480378
rect 359234 460378 359266 460614
rect 359502 460378 359586 460614
rect 359822 460378 359854 460614
rect 359234 440614 359854 460378
rect 359234 440378 359266 440614
rect 359502 440378 359586 440614
rect 359822 440378 359854 440614
rect 359234 421162 359854 440378
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 683294 362414 704282
rect 361794 683058 361826 683294
rect 362062 683058 362146 683294
rect 362382 683058 362414 683294
rect 361794 663294 362414 683058
rect 361794 663058 361826 663294
rect 362062 663058 362146 663294
rect 362382 663058 362414 663294
rect 361794 643294 362414 663058
rect 361794 643058 361826 643294
rect 362062 643058 362146 643294
rect 362382 643058 362414 643294
rect 361794 623294 362414 643058
rect 361794 623058 361826 623294
rect 362062 623058 362146 623294
rect 362382 623058 362414 623294
rect 361794 603294 362414 623058
rect 361794 603058 361826 603294
rect 362062 603058 362146 603294
rect 362382 603058 362414 603294
rect 361794 583294 362414 603058
rect 361794 583058 361826 583294
rect 362062 583058 362146 583294
rect 362382 583058 362414 583294
rect 361794 563294 362414 583058
rect 361794 563058 361826 563294
rect 362062 563058 362146 563294
rect 362382 563058 362414 563294
rect 361794 543294 362414 563058
rect 361794 543058 361826 543294
rect 362062 543058 362146 543294
rect 362382 543058 362414 543294
rect 361794 523294 362414 543058
rect 361794 523058 361826 523294
rect 362062 523058 362146 523294
rect 362382 523058 362414 523294
rect 361794 503294 362414 523058
rect 361794 503058 361826 503294
rect 362062 503058 362146 503294
rect 362382 503058 362414 503294
rect 361794 483294 362414 503058
rect 361794 483058 361826 483294
rect 362062 483058 362146 483294
rect 362382 483058 362414 483294
rect 361794 463294 362414 483058
rect 361794 463058 361826 463294
rect 362062 463058 362146 463294
rect 362382 463058 362414 463294
rect 361794 443294 362414 463058
rect 361794 443058 361826 443294
rect 362062 443058 362146 443294
rect 362382 443058 362414 443294
rect 361794 423294 362414 443058
rect 361794 423058 361826 423294
rect 362062 423058 362146 423294
rect 362382 423058 362414 423294
rect 361794 421162 362414 423058
rect 362954 684274 363574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 362954 684038 362986 684274
rect 363222 684038 363306 684274
rect 363542 684038 363574 684274
rect 362954 664274 363574 684038
rect 362954 664038 362986 664274
rect 363222 664038 363306 664274
rect 363542 664038 363574 664274
rect 362954 644274 363574 664038
rect 362954 644038 362986 644274
rect 363222 644038 363306 644274
rect 363542 644038 363574 644274
rect 362954 624274 363574 644038
rect 362954 624038 362986 624274
rect 363222 624038 363306 624274
rect 363542 624038 363574 624274
rect 362954 604274 363574 624038
rect 362954 604038 362986 604274
rect 363222 604038 363306 604274
rect 363542 604038 363574 604274
rect 362954 584274 363574 604038
rect 362954 584038 362986 584274
rect 363222 584038 363306 584274
rect 363542 584038 363574 584274
rect 362954 564274 363574 584038
rect 362954 564038 362986 564274
rect 363222 564038 363306 564274
rect 363542 564038 363574 564274
rect 362954 544274 363574 564038
rect 362954 544038 362986 544274
rect 363222 544038 363306 544274
rect 363542 544038 363574 544274
rect 362954 524274 363574 544038
rect 362954 524038 362986 524274
rect 363222 524038 363306 524274
rect 363542 524038 363574 524274
rect 362954 504274 363574 524038
rect 362954 504038 362986 504274
rect 363222 504038 363306 504274
rect 363542 504038 363574 504274
rect 362954 484274 363574 504038
rect 362954 484038 362986 484274
rect 363222 484038 363306 484274
rect 363542 484038 363574 484274
rect 362954 464274 363574 484038
rect 362954 464038 362986 464274
rect 363222 464038 363306 464274
rect 363542 464038 363574 464274
rect 362954 444274 363574 464038
rect 362954 444038 362986 444274
rect 363222 444038 363306 444274
rect 363542 444038 363574 444274
rect 362954 424274 363574 444038
rect 362954 424038 362986 424274
rect 363222 424038 363306 424274
rect 363542 424038 363574 424274
rect 362954 421162 363574 424038
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 365514 686954 366134 706202
rect 365514 686718 365546 686954
rect 365782 686718 365866 686954
rect 366102 686718 366134 686954
rect 365514 666954 366134 686718
rect 365514 666718 365546 666954
rect 365782 666718 365866 666954
rect 366102 666718 366134 666954
rect 365514 646954 366134 666718
rect 365514 646718 365546 646954
rect 365782 646718 365866 646954
rect 366102 646718 366134 646954
rect 365514 626954 366134 646718
rect 365514 626718 365546 626954
rect 365782 626718 365866 626954
rect 366102 626718 366134 626954
rect 365514 606954 366134 626718
rect 365514 606718 365546 606954
rect 365782 606718 365866 606954
rect 366102 606718 366134 606954
rect 365514 586954 366134 606718
rect 365514 586718 365546 586954
rect 365782 586718 365866 586954
rect 366102 586718 366134 586954
rect 365514 566954 366134 586718
rect 365514 566718 365546 566954
rect 365782 566718 365866 566954
rect 366102 566718 366134 566954
rect 365514 546954 366134 566718
rect 365514 546718 365546 546954
rect 365782 546718 365866 546954
rect 366102 546718 366134 546954
rect 365514 526954 366134 546718
rect 365514 526718 365546 526954
rect 365782 526718 365866 526954
rect 366102 526718 366134 526954
rect 365514 506954 366134 526718
rect 365514 506718 365546 506954
rect 365782 506718 365866 506954
rect 366102 506718 366134 506954
rect 365514 486954 366134 506718
rect 365514 486718 365546 486954
rect 365782 486718 365866 486954
rect 366102 486718 366134 486954
rect 365514 466954 366134 486718
rect 365514 466718 365546 466954
rect 365782 466718 365866 466954
rect 366102 466718 366134 466954
rect 365514 446954 366134 466718
rect 365514 446718 365546 446954
rect 365782 446718 365866 446954
rect 366102 446718 366134 446954
rect 365514 426954 366134 446718
rect 365514 426718 365546 426954
rect 365782 426718 365866 426954
rect 366102 426718 366134 426954
rect 365514 421162 366134 426718
rect 369234 690614 369854 708122
rect 369234 690378 369266 690614
rect 369502 690378 369586 690614
rect 369822 690378 369854 690614
rect 369234 670614 369854 690378
rect 369234 670378 369266 670614
rect 369502 670378 369586 670614
rect 369822 670378 369854 670614
rect 369234 650614 369854 670378
rect 369234 650378 369266 650614
rect 369502 650378 369586 650614
rect 369822 650378 369854 650614
rect 369234 630614 369854 650378
rect 369234 630378 369266 630614
rect 369502 630378 369586 630614
rect 369822 630378 369854 630614
rect 369234 610614 369854 630378
rect 369234 610378 369266 610614
rect 369502 610378 369586 610614
rect 369822 610378 369854 610614
rect 369234 590614 369854 610378
rect 369234 590378 369266 590614
rect 369502 590378 369586 590614
rect 369822 590378 369854 590614
rect 369234 570614 369854 590378
rect 369234 570378 369266 570614
rect 369502 570378 369586 570614
rect 369822 570378 369854 570614
rect 369234 550614 369854 570378
rect 369234 550378 369266 550614
rect 369502 550378 369586 550614
rect 369822 550378 369854 550614
rect 369234 530614 369854 550378
rect 369234 530378 369266 530614
rect 369502 530378 369586 530614
rect 369822 530378 369854 530614
rect 369234 510614 369854 530378
rect 369234 510378 369266 510614
rect 369502 510378 369586 510614
rect 369822 510378 369854 510614
rect 369234 490614 369854 510378
rect 369234 490378 369266 490614
rect 369502 490378 369586 490614
rect 369822 490378 369854 490614
rect 369234 470614 369854 490378
rect 369234 470378 369266 470614
rect 369502 470378 369586 470614
rect 369822 470378 369854 470614
rect 369234 450614 369854 470378
rect 369234 450378 369266 450614
rect 369502 450378 369586 450614
rect 369822 450378 369854 450614
rect 369234 430614 369854 450378
rect 369234 430378 369266 430614
rect 369502 430378 369586 430614
rect 369822 430378 369854 430614
rect 369234 421162 369854 430378
rect 371794 705798 372414 705830
rect 371794 705562 371826 705798
rect 372062 705562 372146 705798
rect 372382 705562 372414 705798
rect 371794 705478 372414 705562
rect 371794 705242 371826 705478
rect 372062 705242 372146 705478
rect 372382 705242 372414 705478
rect 371794 693294 372414 705242
rect 371794 693058 371826 693294
rect 372062 693058 372146 693294
rect 372382 693058 372414 693294
rect 371794 673294 372414 693058
rect 371794 673058 371826 673294
rect 372062 673058 372146 673294
rect 372382 673058 372414 673294
rect 371794 653294 372414 673058
rect 371794 653058 371826 653294
rect 372062 653058 372146 653294
rect 372382 653058 372414 653294
rect 371794 633294 372414 653058
rect 371794 633058 371826 633294
rect 372062 633058 372146 633294
rect 372382 633058 372414 633294
rect 371794 613294 372414 633058
rect 371794 613058 371826 613294
rect 372062 613058 372146 613294
rect 372382 613058 372414 613294
rect 371794 593294 372414 613058
rect 371794 593058 371826 593294
rect 372062 593058 372146 593294
rect 372382 593058 372414 593294
rect 371794 573294 372414 593058
rect 371794 573058 371826 573294
rect 372062 573058 372146 573294
rect 372382 573058 372414 573294
rect 371794 553294 372414 573058
rect 371794 553058 371826 553294
rect 372062 553058 372146 553294
rect 372382 553058 372414 553294
rect 371794 533294 372414 553058
rect 371794 533058 371826 533294
rect 372062 533058 372146 533294
rect 372382 533058 372414 533294
rect 371794 513294 372414 533058
rect 371794 513058 371826 513294
rect 372062 513058 372146 513294
rect 372382 513058 372414 513294
rect 371794 493294 372414 513058
rect 371794 493058 371826 493294
rect 372062 493058 372146 493294
rect 372382 493058 372414 493294
rect 371794 473294 372414 493058
rect 371794 473058 371826 473294
rect 372062 473058 372146 473294
rect 372382 473058 372414 473294
rect 371794 453294 372414 473058
rect 371794 453058 371826 453294
rect 372062 453058 372146 453294
rect 372382 453058 372414 453294
rect 371794 433294 372414 453058
rect 371794 433058 371826 433294
rect 372062 433058 372146 433294
rect 372382 433058 372414 433294
rect 371794 421162 372414 433058
rect 372954 694274 373574 710042
rect 382954 711558 383574 711590
rect 382954 711322 382986 711558
rect 383222 711322 383306 711558
rect 383542 711322 383574 711558
rect 382954 711238 383574 711322
rect 382954 711002 382986 711238
rect 383222 711002 383306 711238
rect 383542 711002 383574 711238
rect 379234 709638 379854 709670
rect 379234 709402 379266 709638
rect 379502 709402 379586 709638
rect 379822 709402 379854 709638
rect 379234 709318 379854 709402
rect 379234 709082 379266 709318
rect 379502 709082 379586 709318
rect 379822 709082 379854 709318
rect 372954 694038 372986 694274
rect 373222 694038 373306 694274
rect 373542 694038 373574 694274
rect 372954 674274 373574 694038
rect 372954 674038 372986 674274
rect 373222 674038 373306 674274
rect 373542 674038 373574 674274
rect 372954 654274 373574 674038
rect 372954 654038 372986 654274
rect 373222 654038 373306 654274
rect 373542 654038 373574 654274
rect 372954 634274 373574 654038
rect 372954 634038 372986 634274
rect 373222 634038 373306 634274
rect 373542 634038 373574 634274
rect 372954 614274 373574 634038
rect 372954 614038 372986 614274
rect 373222 614038 373306 614274
rect 373542 614038 373574 614274
rect 372954 594274 373574 614038
rect 372954 594038 372986 594274
rect 373222 594038 373306 594274
rect 373542 594038 373574 594274
rect 372954 574274 373574 594038
rect 372954 574038 372986 574274
rect 373222 574038 373306 574274
rect 373542 574038 373574 574274
rect 372954 554274 373574 574038
rect 372954 554038 372986 554274
rect 373222 554038 373306 554274
rect 373542 554038 373574 554274
rect 372954 534274 373574 554038
rect 372954 534038 372986 534274
rect 373222 534038 373306 534274
rect 373542 534038 373574 534274
rect 372954 514274 373574 534038
rect 372954 514038 372986 514274
rect 373222 514038 373306 514274
rect 373542 514038 373574 514274
rect 372954 494274 373574 514038
rect 372954 494038 372986 494274
rect 373222 494038 373306 494274
rect 373542 494038 373574 494274
rect 372954 474274 373574 494038
rect 372954 474038 372986 474274
rect 373222 474038 373306 474274
rect 373542 474038 373574 474274
rect 372954 454274 373574 474038
rect 372954 454038 372986 454274
rect 373222 454038 373306 454274
rect 373542 454038 373574 454274
rect 372954 434274 373574 454038
rect 372954 434038 372986 434274
rect 373222 434038 373306 434274
rect 373542 434038 373574 434274
rect 372954 421162 373574 434038
rect 375514 707718 376134 707750
rect 375514 707482 375546 707718
rect 375782 707482 375866 707718
rect 376102 707482 376134 707718
rect 375514 707398 376134 707482
rect 375514 707162 375546 707398
rect 375782 707162 375866 707398
rect 376102 707162 376134 707398
rect 375514 696954 376134 707162
rect 375514 696718 375546 696954
rect 375782 696718 375866 696954
rect 376102 696718 376134 696954
rect 375514 676954 376134 696718
rect 375514 676718 375546 676954
rect 375782 676718 375866 676954
rect 376102 676718 376134 676954
rect 375514 656954 376134 676718
rect 375514 656718 375546 656954
rect 375782 656718 375866 656954
rect 376102 656718 376134 656954
rect 375514 636954 376134 656718
rect 375514 636718 375546 636954
rect 375782 636718 375866 636954
rect 376102 636718 376134 636954
rect 375514 616954 376134 636718
rect 375514 616718 375546 616954
rect 375782 616718 375866 616954
rect 376102 616718 376134 616954
rect 375514 596954 376134 616718
rect 375514 596718 375546 596954
rect 375782 596718 375866 596954
rect 376102 596718 376134 596954
rect 375514 576954 376134 596718
rect 375514 576718 375546 576954
rect 375782 576718 375866 576954
rect 376102 576718 376134 576954
rect 375514 556954 376134 576718
rect 375514 556718 375546 556954
rect 375782 556718 375866 556954
rect 376102 556718 376134 556954
rect 375514 536954 376134 556718
rect 375514 536718 375546 536954
rect 375782 536718 375866 536954
rect 376102 536718 376134 536954
rect 375514 516954 376134 536718
rect 375514 516718 375546 516954
rect 375782 516718 375866 516954
rect 376102 516718 376134 516954
rect 375514 496954 376134 516718
rect 375514 496718 375546 496954
rect 375782 496718 375866 496954
rect 376102 496718 376134 496954
rect 375514 476954 376134 496718
rect 375514 476718 375546 476954
rect 375782 476718 375866 476954
rect 376102 476718 376134 476954
rect 375514 456954 376134 476718
rect 375514 456718 375546 456954
rect 375782 456718 375866 456954
rect 376102 456718 376134 456954
rect 375514 436954 376134 456718
rect 375514 436718 375546 436954
rect 375782 436718 375866 436954
rect 376102 436718 376134 436954
rect 375514 421162 376134 436718
rect 379234 700614 379854 709082
rect 379234 700378 379266 700614
rect 379502 700378 379586 700614
rect 379822 700378 379854 700614
rect 379234 680614 379854 700378
rect 379234 680378 379266 680614
rect 379502 680378 379586 680614
rect 379822 680378 379854 680614
rect 379234 660614 379854 680378
rect 379234 660378 379266 660614
rect 379502 660378 379586 660614
rect 379822 660378 379854 660614
rect 379234 640614 379854 660378
rect 379234 640378 379266 640614
rect 379502 640378 379586 640614
rect 379822 640378 379854 640614
rect 379234 620614 379854 640378
rect 379234 620378 379266 620614
rect 379502 620378 379586 620614
rect 379822 620378 379854 620614
rect 379234 600614 379854 620378
rect 379234 600378 379266 600614
rect 379502 600378 379586 600614
rect 379822 600378 379854 600614
rect 379234 580614 379854 600378
rect 379234 580378 379266 580614
rect 379502 580378 379586 580614
rect 379822 580378 379854 580614
rect 379234 560614 379854 580378
rect 379234 560378 379266 560614
rect 379502 560378 379586 560614
rect 379822 560378 379854 560614
rect 379234 540614 379854 560378
rect 379234 540378 379266 540614
rect 379502 540378 379586 540614
rect 379822 540378 379854 540614
rect 379234 520614 379854 540378
rect 379234 520378 379266 520614
rect 379502 520378 379586 520614
rect 379822 520378 379854 520614
rect 379234 500614 379854 520378
rect 379234 500378 379266 500614
rect 379502 500378 379586 500614
rect 379822 500378 379854 500614
rect 379234 480614 379854 500378
rect 379234 480378 379266 480614
rect 379502 480378 379586 480614
rect 379822 480378 379854 480614
rect 379234 460614 379854 480378
rect 379234 460378 379266 460614
rect 379502 460378 379586 460614
rect 379822 460378 379854 460614
rect 379234 440614 379854 460378
rect 379234 440378 379266 440614
rect 379502 440378 379586 440614
rect 379822 440378 379854 440614
rect 379234 421162 379854 440378
rect 381794 704838 382414 705830
rect 381794 704602 381826 704838
rect 382062 704602 382146 704838
rect 382382 704602 382414 704838
rect 381794 704518 382414 704602
rect 381794 704282 381826 704518
rect 382062 704282 382146 704518
rect 382382 704282 382414 704518
rect 381794 683294 382414 704282
rect 381794 683058 381826 683294
rect 382062 683058 382146 683294
rect 382382 683058 382414 683294
rect 381794 663294 382414 683058
rect 381794 663058 381826 663294
rect 382062 663058 382146 663294
rect 382382 663058 382414 663294
rect 381794 643294 382414 663058
rect 381794 643058 381826 643294
rect 382062 643058 382146 643294
rect 382382 643058 382414 643294
rect 381794 623294 382414 643058
rect 381794 623058 381826 623294
rect 382062 623058 382146 623294
rect 382382 623058 382414 623294
rect 381794 603294 382414 623058
rect 381794 603058 381826 603294
rect 382062 603058 382146 603294
rect 382382 603058 382414 603294
rect 381794 583294 382414 603058
rect 381794 583058 381826 583294
rect 382062 583058 382146 583294
rect 382382 583058 382414 583294
rect 381794 563294 382414 583058
rect 381794 563058 381826 563294
rect 382062 563058 382146 563294
rect 382382 563058 382414 563294
rect 381794 543294 382414 563058
rect 381794 543058 381826 543294
rect 382062 543058 382146 543294
rect 382382 543058 382414 543294
rect 381794 523294 382414 543058
rect 381794 523058 381826 523294
rect 382062 523058 382146 523294
rect 382382 523058 382414 523294
rect 381794 503294 382414 523058
rect 381794 503058 381826 503294
rect 382062 503058 382146 503294
rect 382382 503058 382414 503294
rect 381794 483294 382414 503058
rect 381794 483058 381826 483294
rect 382062 483058 382146 483294
rect 382382 483058 382414 483294
rect 381794 463294 382414 483058
rect 381794 463058 381826 463294
rect 382062 463058 382146 463294
rect 382382 463058 382414 463294
rect 381794 443294 382414 463058
rect 381794 443058 381826 443294
rect 382062 443058 382146 443294
rect 382382 443058 382414 443294
rect 381794 423294 382414 443058
rect 381794 423058 381826 423294
rect 382062 423058 382146 423294
rect 382382 423058 382414 423294
rect 381794 421162 382414 423058
rect 382954 684274 383574 711002
rect 392954 710598 393574 711590
rect 392954 710362 392986 710598
rect 393222 710362 393306 710598
rect 393542 710362 393574 710598
rect 392954 710278 393574 710362
rect 392954 710042 392986 710278
rect 393222 710042 393306 710278
rect 393542 710042 393574 710278
rect 389234 708678 389854 709670
rect 389234 708442 389266 708678
rect 389502 708442 389586 708678
rect 389822 708442 389854 708678
rect 389234 708358 389854 708442
rect 389234 708122 389266 708358
rect 389502 708122 389586 708358
rect 389822 708122 389854 708358
rect 382954 684038 382986 684274
rect 383222 684038 383306 684274
rect 383542 684038 383574 684274
rect 382954 664274 383574 684038
rect 382954 664038 382986 664274
rect 383222 664038 383306 664274
rect 383542 664038 383574 664274
rect 382954 644274 383574 664038
rect 382954 644038 382986 644274
rect 383222 644038 383306 644274
rect 383542 644038 383574 644274
rect 382954 624274 383574 644038
rect 382954 624038 382986 624274
rect 383222 624038 383306 624274
rect 383542 624038 383574 624274
rect 382954 604274 383574 624038
rect 382954 604038 382986 604274
rect 383222 604038 383306 604274
rect 383542 604038 383574 604274
rect 382954 584274 383574 604038
rect 382954 584038 382986 584274
rect 383222 584038 383306 584274
rect 383542 584038 383574 584274
rect 382954 564274 383574 584038
rect 382954 564038 382986 564274
rect 383222 564038 383306 564274
rect 383542 564038 383574 564274
rect 382954 544274 383574 564038
rect 382954 544038 382986 544274
rect 383222 544038 383306 544274
rect 383542 544038 383574 544274
rect 382954 524274 383574 544038
rect 382954 524038 382986 524274
rect 383222 524038 383306 524274
rect 383542 524038 383574 524274
rect 382954 504274 383574 524038
rect 382954 504038 382986 504274
rect 383222 504038 383306 504274
rect 383542 504038 383574 504274
rect 382954 484274 383574 504038
rect 382954 484038 382986 484274
rect 383222 484038 383306 484274
rect 383542 484038 383574 484274
rect 382954 464274 383574 484038
rect 382954 464038 382986 464274
rect 383222 464038 383306 464274
rect 383542 464038 383574 464274
rect 382954 444274 383574 464038
rect 382954 444038 382986 444274
rect 383222 444038 383306 444274
rect 383542 444038 383574 444274
rect 382954 424274 383574 444038
rect 382954 424038 382986 424274
rect 383222 424038 383306 424274
rect 383542 424038 383574 424274
rect 382954 421162 383574 424038
rect 385514 706758 386134 707750
rect 385514 706522 385546 706758
rect 385782 706522 385866 706758
rect 386102 706522 386134 706758
rect 385514 706438 386134 706522
rect 385514 706202 385546 706438
rect 385782 706202 385866 706438
rect 386102 706202 386134 706438
rect 385514 686954 386134 706202
rect 385514 686718 385546 686954
rect 385782 686718 385866 686954
rect 386102 686718 386134 686954
rect 385514 666954 386134 686718
rect 385514 666718 385546 666954
rect 385782 666718 385866 666954
rect 386102 666718 386134 666954
rect 385514 646954 386134 666718
rect 385514 646718 385546 646954
rect 385782 646718 385866 646954
rect 386102 646718 386134 646954
rect 385514 626954 386134 646718
rect 385514 626718 385546 626954
rect 385782 626718 385866 626954
rect 386102 626718 386134 626954
rect 385514 606954 386134 626718
rect 385514 606718 385546 606954
rect 385782 606718 385866 606954
rect 386102 606718 386134 606954
rect 385514 586954 386134 606718
rect 385514 586718 385546 586954
rect 385782 586718 385866 586954
rect 386102 586718 386134 586954
rect 385514 566954 386134 586718
rect 385514 566718 385546 566954
rect 385782 566718 385866 566954
rect 386102 566718 386134 566954
rect 385514 546954 386134 566718
rect 385514 546718 385546 546954
rect 385782 546718 385866 546954
rect 386102 546718 386134 546954
rect 385514 526954 386134 546718
rect 385514 526718 385546 526954
rect 385782 526718 385866 526954
rect 386102 526718 386134 526954
rect 385514 506954 386134 526718
rect 385514 506718 385546 506954
rect 385782 506718 385866 506954
rect 386102 506718 386134 506954
rect 385514 486954 386134 506718
rect 385514 486718 385546 486954
rect 385782 486718 385866 486954
rect 386102 486718 386134 486954
rect 385514 466954 386134 486718
rect 385514 466718 385546 466954
rect 385782 466718 385866 466954
rect 386102 466718 386134 466954
rect 385514 446954 386134 466718
rect 385514 446718 385546 446954
rect 385782 446718 385866 446954
rect 386102 446718 386134 446954
rect 385514 426954 386134 446718
rect 385514 426718 385546 426954
rect 385782 426718 385866 426954
rect 386102 426718 386134 426954
rect 385514 421162 386134 426718
rect 389234 690614 389854 708122
rect 389234 690378 389266 690614
rect 389502 690378 389586 690614
rect 389822 690378 389854 690614
rect 389234 670614 389854 690378
rect 389234 670378 389266 670614
rect 389502 670378 389586 670614
rect 389822 670378 389854 670614
rect 389234 650614 389854 670378
rect 389234 650378 389266 650614
rect 389502 650378 389586 650614
rect 389822 650378 389854 650614
rect 389234 630614 389854 650378
rect 389234 630378 389266 630614
rect 389502 630378 389586 630614
rect 389822 630378 389854 630614
rect 389234 610614 389854 630378
rect 389234 610378 389266 610614
rect 389502 610378 389586 610614
rect 389822 610378 389854 610614
rect 389234 590614 389854 610378
rect 389234 590378 389266 590614
rect 389502 590378 389586 590614
rect 389822 590378 389854 590614
rect 389234 570614 389854 590378
rect 389234 570378 389266 570614
rect 389502 570378 389586 570614
rect 389822 570378 389854 570614
rect 389234 550614 389854 570378
rect 389234 550378 389266 550614
rect 389502 550378 389586 550614
rect 389822 550378 389854 550614
rect 389234 530614 389854 550378
rect 389234 530378 389266 530614
rect 389502 530378 389586 530614
rect 389822 530378 389854 530614
rect 389234 510614 389854 530378
rect 389234 510378 389266 510614
rect 389502 510378 389586 510614
rect 389822 510378 389854 510614
rect 389234 490614 389854 510378
rect 389234 490378 389266 490614
rect 389502 490378 389586 490614
rect 389822 490378 389854 490614
rect 389234 470614 389854 490378
rect 389234 470378 389266 470614
rect 389502 470378 389586 470614
rect 389822 470378 389854 470614
rect 389234 450614 389854 470378
rect 389234 450378 389266 450614
rect 389502 450378 389586 450614
rect 389822 450378 389854 450614
rect 389234 430614 389854 450378
rect 389234 430378 389266 430614
rect 389502 430378 389586 430614
rect 389822 430378 389854 430614
rect 389234 421162 389854 430378
rect 391794 705798 392414 705830
rect 391794 705562 391826 705798
rect 392062 705562 392146 705798
rect 392382 705562 392414 705798
rect 391794 705478 392414 705562
rect 391794 705242 391826 705478
rect 392062 705242 392146 705478
rect 392382 705242 392414 705478
rect 391794 693294 392414 705242
rect 391794 693058 391826 693294
rect 392062 693058 392146 693294
rect 392382 693058 392414 693294
rect 391794 673294 392414 693058
rect 391794 673058 391826 673294
rect 392062 673058 392146 673294
rect 392382 673058 392414 673294
rect 391794 653294 392414 673058
rect 391794 653058 391826 653294
rect 392062 653058 392146 653294
rect 392382 653058 392414 653294
rect 391794 633294 392414 653058
rect 391794 633058 391826 633294
rect 392062 633058 392146 633294
rect 392382 633058 392414 633294
rect 391794 613294 392414 633058
rect 391794 613058 391826 613294
rect 392062 613058 392146 613294
rect 392382 613058 392414 613294
rect 391794 593294 392414 613058
rect 391794 593058 391826 593294
rect 392062 593058 392146 593294
rect 392382 593058 392414 593294
rect 391794 573294 392414 593058
rect 391794 573058 391826 573294
rect 392062 573058 392146 573294
rect 392382 573058 392414 573294
rect 391794 553294 392414 573058
rect 391794 553058 391826 553294
rect 392062 553058 392146 553294
rect 392382 553058 392414 553294
rect 391794 533294 392414 553058
rect 391794 533058 391826 533294
rect 392062 533058 392146 533294
rect 392382 533058 392414 533294
rect 391794 513294 392414 533058
rect 391794 513058 391826 513294
rect 392062 513058 392146 513294
rect 392382 513058 392414 513294
rect 391794 493294 392414 513058
rect 391794 493058 391826 493294
rect 392062 493058 392146 493294
rect 392382 493058 392414 493294
rect 391794 473294 392414 493058
rect 391794 473058 391826 473294
rect 392062 473058 392146 473294
rect 392382 473058 392414 473294
rect 391794 453294 392414 473058
rect 391794 453058 391826 453294
rect 392062 453058 392146 453294
rect 392382 453058 392414 453294
rect 391794 433294 392414 453058
rect 391794 433058 391826 433294
rect 392062 433058 392146 433294
rect 392382 433058 392414 433294
rect 391794 421162 392414 433058
rect 392954 694274 393574 710042
rect 402954 711558 403574 711590
rect 402954 711322 402986 711558
rect 403222 711322 403306 711558
rect 403542 711322 403574 711558
rect 402954 711238 403574 711322
rect 402954 711002 402986 711238
rect 403222 711002 403306 711238
rect 403542 711002 403574 711238
rect 399234 709638 399854 709670
rect 399234 709402 399266 709638
rect 399502 709402 399586 709638
rect 399822 709402 399854 709638
rect 399234 709318 399854 709402
rect 399234 709082 399266 709318
rect 399502 709082 399586 709318
rect 399822 709082 399854 709318
rect 392954 694038 392986 694274
rect 393222 694038 393306 694274
rect 393542 694038 393574 694274
rect 392954 674274 393574 694038
rect 392954 674038 392986 674274
rect 393222 674038 393306 674274
rect 393542 674038 393574 674274
rect 392954 654274 393574 674038
rect 392954 654038 392986 654274
rect 393222 654038 393306 654274
rect 393542 654038 393574 654274
rect 392954 634274 393574 654038
rect 392954 634038 392986 634274
rect 393222 634038 393306 634274
rect 393542 634038 393574 634274
rect 392954 614274 393574 634038
rect 392954 614038 392986 614274
rect 393222 614038 393306 614274
rect 393542 614038 393574 614274
rect 392954 594274 393574 614038
rect 392954 594038 392986 594274
rect 393222 594038 393306 594274
rect 393542 594038 393574 594274
rect 392954 574274 393574 594038
rect 392954 574038 392986 574274
rect 393222 574038 393306 574274
rect 393542 574038 393574 574274
rect 392954 554274 393574 574038
rect 392954 554038 392986 554274
rect 393222 554038 393306 554274
rect 393542 554038 393574 554274
rect 392954 534274 393574 554038
rect 392954 534038 392986 534274
rect 393222 534038 393306 534274
rect 393542 534038 393574 534274
rect 392954 514274 393574 534038
rect 392954 514038 392986 514274
rect 393222 514038 393306 514274
rect 393542 514038 393574 514274
rect 392954 494274 393574 514038
rect 392954 494038 392986 494274
rect 393222 494038 393306 494274
rect 393542 494038 393574 494274
rect 392954 474274 393574 494038
rect 392954 474038 392986 474274
rect 393222 474038 393306 474274
rect 393542 474038 393574 474274
rect 392954 454274 393574 474038
rect 392954 454038 392986 454274
rect 393222 454038 393306 454274
rect 393542 454038 393574 454274
rect 392954 434274 393574 454038
rect 392954 434038 392986 434274
rect 393222 434038 393306 434274
rect 393542 434038 393574 434274
rect 392954 421162 393574 434038
rect 395514 707718 396134 707750
rect 395514 707482 395546 707718
rect 395782 707482 395866 707718
rect 396102 707482 396134 707718
rect 395514 707398 396134 707482
rect 395514 707162 395546 707398
rect 395782 707162 395866 707398
rect 396102 707162 396134 707398
rect 395514 696954 396134 707162
rect 395514 696718 395546 696954
rect 395782 696718 395866 696954
rect 396102 696718 396134 696954
rect 395514 676954 396134 696718
rect 395514 676718 395546 676954
rect 395782 676718 395866 676954
rect 396102 676718 396134 676954
rect 395514 656954 396134 676718
rect 395514 656718 395546 656954
rect 395782 656718 395866 656954
rect 396102 656718 396134 656954
rect 395514 636954 396134 656718
rect 395514 636718 395546 636954
rect 395782 636718 395866 636954
rect 396102 636718 396134 636954
rect 395514 616954 396134 636718
rect 395514 616718 395546 616954
rect 395782 616718 395866 616954
rect 396102 616718 396134 616954
rect 395514 596954 396134 616718
rect 395514 596718 395546 596954
rect 395782 596718 395866 596954
rect 396102 596718 396134 596954
rect 395514 576954 396134 596718
rect 395514 576718 395546 576954
rect 395782 576718 395866 576954
rect 396102 576718 396134 576954
rect 395514 556954 396134 576718
rect 395514 556718 395546 556954
rect 395782 556718 395866 556954
rect 396102 556718 396134 556954
rect 395514 536954 396134 556718
rect 395514 536718 395546 536954
rect 395782 536718 395866 536954
rect 396102 536718 396134 536954
rect 395514 516954 396134 536718
rect 395514 516718 395546 516954
rect 395782 516718 395866 516954
rect 396102 516718 396134 516954
rect 395514 496954 396134 516718
rect 395514 496718 395546 496954
rect 395782 496718 395866 496954
rect 396102 496718 396134 496954
rect 395514 476954 396134 496718
rect 395514 476718 395546 476954
rect 395782 476718 395866 476954
rect 396102 476718 396134 476954
rect 395514 456954 396134 476718
rect 395514 456718 395546 456954
rect 395782 456718 395866 456954
rect 396102 456718 396134 456954
rect 395514 436954 396134 456718
rect 395514 436718 395546 436954
rect 395782 436718 395866 436954
rect 396102 436718 396134 436954
rect 395514 421162 396134 436718
rect 399234 700614 399854 709082
rect 399234 700378 399266 700614
rect 399502 700378 399586 700614
rect 399822 700378 399854 700614
rect 399234 680614 399854 700378
rect 399234 680378 399266 680614
rect 399502 680378 399586 680614
rect 399822 680378 399854 680614
rect 399234 660614 399854 680378
rect 399234 660378 399266 660614
rect 399502 660378 399586 660614
rect 399822 660378 399854 660614
rect 399234 640614 399854 660378
rect 399234 640378 399266 640614
rect 399502 640378 399586 640614
rect 399822 640378 399854 640614
rect 399234 620614 399854 640378
rect 399234 620378 399266 620614
rect 399502 620378 399586 620614
rect 399822 620378 399854 620614
rect 399234 600614 399854 620378
rect 399234 600378 399266 600614
rect 399502 600378 399586 600614
rect 399822 600378 399854 600614
rect 399234 580614 399854 600378
rect 399234 580378 399266 580614
rect 399502 580378 399586 580614
rect 399822 580378 399854 580614
rect 399234 560614 399854 580378
rect 399234 560378 399266 560614
rect 399502 560378 399586 560614
rect 399822 560378 399854 560614
rect 399234 540614 399854 560378
rect 399234 540378 399266 540614
rect 399502 540378 399586 540614
rect 399822 540378 399854 540614
rect 399234 520614 399854 540378
rect 399234 520378 399266 520614
rect 399502 520378 399586 520614
rect 399822 520378 399854 520614
rect 399234 500614 399854 520378
rect 399234 500378 399266 500614
rect 399502 500378 399586 500614
rect 399822 500378 399854 500614
rect 399234 480614 399854 500378
rect 399234 480378 399266 480614
rect 399502 480378 399586 480614
rect 399822 480378 399854 480614
rect 399234 460614 399854 480378
rect 399234 460378 399266 460614
rect 399502 460378 399586 460614
rect 399822 460378 399854 460614
rect 399234 440614 399854 460378
rect 399234 440378 399266 440614
rect 399502 440378 399586 440614
rect 399822 440378 399854 440614
rect 399234 421162 399854 440378
rect 401794 704838 402414 705830
rect 401794 704602 401826 704838
rect 402062 704602 402146 704838
rect 402382 704602 402414 704838
rect 401794 704518 402414 704602
rect 401794 704282 401826 704518
rect 402062 704282 402146 704518
rect 402382 704282 402414 704518
rect 401794 683294 402414 704282
rect 401794 683058 401826 683294
rect 402062 683058 402146 683294
rect 402382 683058 402414 683294
rect 401794 663294 402414 683058
rect 401794 663058 401826 663294
rect 402062 663058 402146 663294
rect 402382 663058 402414 663294
rect 401794 643294 402414 663058
rect 401794 643058 401826 643294
rect 402062 643058 402146 643294
rect 402382 643058 402414 643294
rect 401794 623294 402414 643058
rect 401794 623058 401826 623294
rect 402062 623058 402146 623294
rect 402382 623058 402414 623294
rect 401794 603294 402414 623058
rect 401794 603058 401826 603294
rect 402062 603058 402146 603294
rect 402382 603058 402414 603294
rect 401794 583294 402414 603058
rect 401794 583058 401826 583294
rect 402062 583058 402146 583294
rect 402382 583058 402414 583294
rect 401794 563294 402414 583058
rect 401794 563058 401826 563294
rect 402062 563058 402146 563294
rect 402382 563058 402414 563294
rect 401794 543294 402414 563058
rect 401794 543058 401826 543294
rect 402062 543058 402146 543294
rect 402382 543058 402414 543294
rect 401794 523294 402414 543058
rect 401794 523058 401826 523294
rect 402062 523058 402146 523294
rect 402382 523058 402414 523294
rect 401794 503294 402414 523058
rect 401794 503058 401826 503294
rect 402062 503058 402146 503294
rect 402382 503058 402414 503294
rect 401794 483294 402414 503058
rect 401794 483058 401826 483294
rect 402062 483058 402146 483294
rect 402382 483058 402414 483294
rect 401794 463294 402414 483058
rect 401794 463058 401826 463294
rect 402062 463058 402146 463294
rect 402382 463058 402414 463294
rect 401794 443294 402414 463058
rect 401794 443058 401826 443294
rect 402062 443058 402146 443294
rect 402382 443058 402414 443294
rect 401794 423294 402414 443058
rect 401794 423058 401826 423294
rect 402062 423058 402146 423294
rect 402382 423058 402414 423294
rect 401794 421162 402414 423058
rect 402954 684274 403574 711002
rect 412954 710598 413574 711590
rect 412954 710362 412986 710598
rect 413222 710362 413306 710598
rect 413542 710362 413574 710598
rect 412954 710278 413574 710362
rect 412954 710042 412986 710278
rect 413222 710042 413306 710278
rect 413542 710042 413574 710278
rect 409234 708678 409854 709670
rect 409234 708442 409266 708678
rect 409502 708442 409586 708678
rect 409822 708442 409854 708678
rect 409234 708358 409854 708442
rect 409234 708122 409266 708358
rect 409502 708122 409586 708358
rect 409822 708122 409854 708358
rect 402954 684038 402986 684274
rect 403222 684038 403306 684274
rect 403542 684038 403574 684274
rect 402954 664274 403574 684038
rect 402954 664038 402986 664274
rect 403222 664038 403306 664274
rect 403542 664038 403574 664274
rect 402954 644274 403574 664038
rect 402954 644038 402986 644274
rect 403222 644038 403306 644274
rect 403542 644038 403574 644274
rect 402954 624274 403574 644038
rect 402954 624038 402986 624274
rect 403222 624038 403306 624274
rect 403542 624038 403574 624274
rect 402954 604274 403574 624038
rect 402954 604038 402986 604274
rect 403222 604038 403306 604274
rect 403542 604038 403574 604274
rect 402954 584274 403574 604038
rect 402954 584038 402986 584274
rect 403222 584038 403306 584274
rect 403542 584038 403574 584274
rect 402954 564274 403574 584038
rect 402954 564038 402986 564274
rect 403222 564038 403306 564274
rect 403542 564038 403574 564274
rect 402954 544274 403574 564038
rect 402954 544038 402986 544274
rect 403222 544038 403306 544274
rect 403542 544038 403574 544274
rect 402954 524274 403574 544038
rect 402954 524038 402986 524274
rect 403222 524038 403306 524274
rect 403542 524038 403574 524274
rect 402954 504274 403574 524038
rect 402954 504038 402986 504274
rect 403222 504038 403306 504274
rect 403542 504038 403574 504274
rect 402954 484274 403574 504038
rect 402954 484038 402986 484274
rect 403222 484038 403306 484274
rect 403542 484038 403574 484274
rect 402954 464274 403574 484038
rect 402954 464038 402986 464274
rect 403222 464038 403306 464274
rect 403542 464038 403574 464274
rect 402954 444274 403574 464038
rect 402954 444038 402986 444274
rect 403222 444038 403306 444274
rect 403542 444038 403574 444274
rect 402954 424274 403574 444038
rect 402954 424038 402986 424274
rect 403222 424038 403306 424274
rect 403542 424038 403574 424274
rect 402954 421162 403574 424038
rect 405514 706758 406134 707750
rect 405514 706522 405546 706758
rect 405782 706522 405866 706758
rect 406102 706522 406134 706758
rect 405514 706438 406134 706522
rect 405514 706202 405546 706438
rect 405782 706202 405866 706438
rect 406102 706202 406134 706438
rect 405514 686954 406134 706202
rect 405514 686718 405546 686954
rect 405782 686718 405866 686954
rect 406102 686718 406134 686954
rect 405514 666954 406134 686718
rect 405514 666718 405546 666954
rect 405782 666718 405866 666954
rect 406102 666718 406134 666954
rect 405514 646954 406134 666718
rect 409234 690614 409854 708122
rect 409234 690378 409266 690614
rect 409502 690378 409586 690614
rect 409822 690378 409854 690614
rect 409234 670614 409854 690378
rect 409234 670378 409266 670614
rect 409502 670378 409586 670614
rect 409822 670378 409854 670614
rect 409234 659500 409854 670378
rect 411794 705798 412414 705830
rect 411794 705562 411826 705798
rect 412062 705562 412146 705798
rect 412382 705562 412414 705798
rect 411794 705478 412414 705562
rect 411794 705242 411826 705478
rect 412062 705242 412146 705478
rect 412382 705242 412414 705478
rect 411794 693294 412414 705242
rect 411794 693058 411826 693294
rect 412062 693058 412146 693294
rect 412382 693058 412414 693294
rect 411794 673294 412414 693058
rect 411794 673058 411826 673294
rect 412062 673058 412146 673294
rect 412382 673058 412414 673294
rect 411794 659500 412414 673058
rect 412954 694274 413574 710042
rect 422954 711558 423574 711590
rect 422954 711322 422986 711558
rect 423222 711322 423306 711558
rect 423542 711322 423574 711558
rect 422954 711238 423574 711322
rect 422954 711002 422986 711238
rect 423222 711002 423306 711238
rect 423542 711002 423574 711238
rect 419234 709638 419854 709670
rect 419234 709402 419266 709638
rect 419502 709402 419586 709638
rect 419822 709402 419854 709638
rect 419234 709318 419854 709402
rect 419234 709082 419266 709318
rect 419502 709082 419586 709318
rect 419822 709082 419854 709318
rect 412954 694038 412986 694274
rect 413222 694038 413306 694274
rect 413542 694038 413574 694274
rect 412954 674274 413574 694038
rect 412954 674038 412986 674274
rect 413222 674038 413306 674274
rect 413542 674038 413574 674274
rect 412954 659500 413574 674038
rect 415514 707718 416134 707750
rect 415514 707482 415546 707718
rect 415782 707482 415866 707718
rect 416102 707482 416134 707718
rect 415514 707398 416134 707482
rect 415514 707162 415546 707398
rect 415782 707162 415866 707398
rect 416102 707162 416134 707398
rect 415514 696954 416134 707162
rect 415514 696718 415546 696954
rect 415782 696718 415866 696954
rect 416102 696718 416134 696954
rect 415514 676954 416134 696718
rect 415514 676718 415546 676954
rect 415782 676718 415866 676954
rect 416102 676718 416134 676954
rect 415514 659500 416134 676718
rect 419234 700614 419854 709082
rect 419234 700378 419266 700614
rect 419502 700378 419586 700614
rect 419822 700378 419854 700614
rect 419234 680614 419854 700378
rect 419234 680378 419266 680614
rect 419502 680378 419586 680614
rect 419822 680378 419854 680614
rect 419234 660614 419854 680378
rect 419234 660378 419266 660614
rect 419502 660378 419586 660614
rect 419822 660378 419854 660614
rect 419234 659500 419854 660378
rect 421794 704838 422414 705830
rect 421794 704602 421826 704838
rect 422062 704602 422146 704838
rect 422382 704602 422414 704838
rect 421794 704518 422414 704602
rect 421794 704282 421826 704518
rect 422062 704282 422146 704518
rect 422382 704282 422414 704518
rect 421794 683294 422414 704282
rect 421794 683058 421826 683294
rect 422062 683058 422146 683294
rect 422382 683058 422414 683294
rect 421794 663294 422414 683058
rect 421794 663058 421826 663294
rect 422062 663058 422146 663294
rect 422382 663058 422414 663294
rect 421794 659500 422414 663058
rect 422954 684274 423574 711002
rect 432954 710598 433574 711590
rect 432954 710362 432986 710598
rect 433222 710362 433306 710598
rect 433542 710362 433574 710598
rect 432954 710278 433574 710362
rect 432954 710042 432986 710278
rect 433222 710042 433306 710278
rect 433542 710042 433574 710278
rect 429234 708678 429854 709670
rect 429234 708442 429266 708678
rect 429502 708442 429586 708678
rect 429822 708442 429854 708678
rect 429234 708358 429854 708442
rect 429234 708122 429266 708358
rect 429502 708122 429586 708358
rect 429822 708122 429854 708358
rect 422954 684038 422986 684274
rect 423222 684038 423306 684274
rect 423542 684038 423574 684274
rect 422954 664274 423574 684038
rect 422954 664038 422986 664274
rect 423222 664038 423306 664274
rect 423542 664038 423574 664274
rect 422954 659500 423574 664038
rect 425514 706758 426134 707750
rect 425514 706522 425546 706758
rect 425782 706522 425866 706758
rect 426102 706522 426134 706758
rect 425514 706438 426134 706522
rect 425514 706202 425546 706438
rect 425782 706202 425866 706438
rect 426102 706202 426134 706438
rect 425514 686954 426134 706202
rect 425514 686718 425546 686954
rect 425782 686718 425866 686954
rect 426102 686718 426134 686954
rect 425514 666954 426134 686718
rect 425514 666718 425546 666954
rect 425782 666718 425866 666954
rect 426102 666718 426134 666954
rect 425514 659500 426134 666718
rect 429234 690614 429854 708122
rect 429234 690378 429266 690614
rect 429502 690378 429586 690614
rect 429822 690378 429854 690614
rect 429234 670614 429854 690378
rect 429234 670378 429266 670614
rect 429502 670378 429586 670614
rect 429822 670378 429854 670614
rect 429234 659500 429854 670378
rect 431794 705798 432414 705830
rect 431794 705562 431826 705798
rect 432062 705562 432146 705798
rect 432382 705562 432414 705798
rect 431794 705478 432414 705562
rect 431794 705242 431826 705478
rect 432062 705242 432146 705478
rect 432382 705242 432414 705478
rect 431794 693294 432414 705242
rect 431794 693058 431826 693294
rect 432062 693058 432146 693294
rect 432382 693058 432414 693294
rect 431794 673294 432414 693058
rect 431794 673058 431826 673294
rect 432062 673058 432146 673294
rect 432382 673058 432414 673294
rect 431794 659500 432414 673058
rect 432954 694274 433574 710042
rect 442954 711558 443574 711590
rect 442954 711322 442986 711558
rect 443222 711322 443306 711558
rect 443542 711322 443574 711558
rect 442954 711238 443574 711322
rect 442954 711002 442986 711238
rect 443222 711002 443306 711238
rect 443542 711002 443574 711238
rect 439234 709638 439854 709670
rect 439234 709402 439266 709638
rect 439502 709402 439586 709638
rect 439822 709402 439854 709638
rect 439234 709318 439854 709402
rect 439234 709082 439266 709318
rect 439502 709082 439586 709318
rect 439822 709082 439854 709318
rect 432954 694038 432986 694274
rect 433222 694038 433306 694274
rect 433542 694038 433574 694274
rect 432954 674274 433574 694038
rect 432954 674038 432986 674274
rect 433222 674038 433306 674274
rect 433542 674038 433574 674274
rect 432954 659500 433574 674038
rect 435514 707718 436134 707750
rect 435514 707482 435546 707718
rect 435782 707482 435866 707718
rect 436102 707482 436134 707718
rect 435514 707398 436134 707482
rect 435514 707162 435546 707398
rect 435782 707162 435866 707398
rect 436102 707162 436134 707398
rect 435514 696954 436134 707162
rect 435514 696718 435546 696954
rect 435782 696718 435866 696954
rect 436102 696718 436134 696954
rect 435514 676954 436134 696718
rect 435514 676718 435546 676954
rect 435782 676718 435866 676954
rect 436102 676718 436134 676954
rect 435514 659500 436134 676718
rect 439234 700614 439854 709082
rect 439234 700378 439266 700614
rect 439502 700378 439586 700614
rect 439822 700378 439854 700614
rect 439234 680614 439854 700378
rect 439234 680378 439266 680614
rect 439502 680378 439586 680614
rect 439822 680378 439854 680614
rect 439234 660614 439854 680378
rect 439234 660378 439266 660614
rect 439502 660378 439586 660614
rect 439822 660378 439854 660614
rect 439234 659500 439854 660378
rect 441794 704838 442414 705830
rect 441794 704602 441826 704838
rect 442062 704602 442146 704838
rect 442382 704602 442414 704838
rect 441794 704518 442414 704602
rect 441794 704282 441826 704518
rect 442062 704282 442146 704518
rect 442382 704282 442414 704518
rect 441794 683294 442414 704282
rect 441794 683058 441826 683294
rect 442062 683058 442146 683294
rect 442382 683058 442414 683294
rect 441794 663294 442414 683058
rect 441794 663058 441826 663294
rect 442062 663058 442146 663294
rect 442382 663058 442414 663294
rect 441794 659500 442414 663058
rect 442954 684274 443574 711002
rect 452954 710598 453574 711590
rect 452954 710362 452986 710598
rect 453222 710362 453306 710598
rect 453542 710362 453574 710598
rect 452954 710278 453574 710362
rect 452954 710042 452986 710278
rect 453222 710042 453306 710278
rect 453542 710042 453574 710278
rect 449234 708678 449854 709670
rect 449234 708442 449266 708678
rect 449502 708442 449586 708678
rect 449822 708442 449854 708678
rect 449234 708358 449854 708442
rect 449234 708122 449266 708358
rect 449502 708122 449586 708358
rect 449822 708122 449854 708358
rect 442954 684038 442986 684274
rect 443222 684038 443306 684274
rect 443542 684038 443574 684274
rect 442954 664274 443574 684038
rect 442954 664038 442986 664274
rect 443222 664038 443306 664274
rect 443542 664038 443574 664274
rect 442954 659500 443574 664038
rect 445514 706758 446134 707750
rect 445514 706522 445546 706758
rect 445782 706522 445866 706758
rect 446102 706522 446134 706758
rect 445514 706438 446134 706522
rect 445514 706202 445546 706438
rect 445782 706202 445866 706438
rect 446102 706202 446134 706438
rect 445514 686954 446134 706202
rect 445514 686718 445546 686954
rect 445782 686718 445866 686954
rect 446102 686718 446134 686954
rect 445514 666954 446134 686718
rect 445514 666718 445546 666954
rect 445782 666718 445866 666954
rect 446102 666718 446134 666954
rect 445514 659500 446134 666718
rect 449234 690614 449854 708122
rect 449234 690378 449266 690614
rect 449502 690378 449586 690614
rect 449822 690378 449854 690614
rect 449234 670614 449854 690378
rect 449234 670378 449266 670614
rect 449502 670378 449586 670614
rect 449822 670378 449854 670614
rect 449234 659500 449854 670378
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 693294 452414 705242
rect 451794 693058 451826 693294
rect 452062 693058 452146 693294
rect 452382 693058 452414 693294
rect 451794 673294 452414 693058
rect 451794 673058 451826 673294
rect 452062 673058 452146 673294
rect 452382 673058 452414 673294
rect 451794 659500 452414 673058
rect 452954 694274 453574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 452954 694038 452986 694274
rect 453222 694038 453306 694274
rect 453542 694038 453574 694274
rect 452954 674274 453574 694038
rect 452954 674038 452986 674274
rect 453222 674038 453306 674274
rect 453542 674038 453574 674274
rect 452954 659500 453574 674038
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 455514 696954 456134 707162
rect 455514 696718 455546 696954
rect 455782 696718 455866 696954
rect 456102 696718 456134 696954
rect 455514 676954 456134 696718
rect 455514 676718 455546 676954
rect 455782 676718 455866 676954
rect 456102 676718 456134 676954
rect 455514 659500 456134 676718
rect 459234 700614 459854 709082
rect 459234 700378 459266 700614
rect 459502 700378 459586 700614
rect 459822 700378 459854 700614
rect 459234 680614 459854 700378
rect 459234 680378 459266 680614
rect 459502 680378 459586 680614
rect 459822 680378 459854 680614
rect 459234 660614 459854 680378
rect 459234 660378 459266 660614
rect 459502 660378 459586 660614
rect 459822 660378 459854 660614
rect 459234 659500 459854 660378
rect 461794 704838 462414 705830
rect 461794 704602 461826 704838
rect 462062 704602 462146 704838
rect 462382 704602 462414 704838
rect 461794 704518 462414 704602
rect 461794 704282 461826 704518
rect 462062 704282 462146 704518
rect 462382 704282 462414 704518
rect 461794 683294 462414 704282
rect 461794 683058 461826 683294
rect 462062 683058 462146 683294
rect 462382 683058 462414 683294
rect 461794 663294 462414 683058
rect 461794 663058 461826 663294
rect 462062 663058 462146 663294
rect 462382 663058 462414 663294
rect 461794 659500 462414 663058
rect 462954 684274 463574 711002
rect 472954 710598 473574 711590
rect 472954 710362 472986 710598
rect 473222 710362 473306 710598
rect 473542 710362 473574 710598
rect 472954 710278 473574 710362
rect 472954 710042 472986 710278
rect 473222 710042 473306 710278
rect 473542 710042 473574 710278
rect 469234 708678 469854 709670
rect 469234 708442 469266 708678
rect 469502 708442 469586 708678
rect 469822 708442 469854 708678
rect 469234 708358 469854 708442
rect 469234 708122 469266 708358
rect 469502 708122 469586 708358
rect 469822 708122 469854 708358
rect 462954 684038 462986 684274
rect 463222 684038 463306 684274
rect 463542 684038 463574 684274
rect 462954 664274 463574 684038
rect 462954 664038 462986 664274
rect 463222 664038 463306 664274
rect 463542 664038 463574 664274
rect 462954 659500 463574 664038
rect 465514 706758 466134 707750
rect 465514 706522 465546 706758
rect 465782 706522 465866 706758
rect 466102 706522 466134 706758
rect 465514 706438 466134 706522
rect 465514 706202 465546 706438
rect 465782 706202 465866 706438
rect 466102 706202 466134 706438
rect 465514 686954 466134 706202
rect 465514 686718 465546 686954
rect 465782 686718 465866 686954
rect 466102 686718 466134 686954
rect 465514 666954 466134 686718
rect 465514 666718 465546 666954
rect 465782 666718 465866 666954
rect 466102 666718 466134 666954
rect 465514 659500 466134 666718
rect 469234 690614 469854 708122
rect 469234 690378 469266 690614
rect 469502 690378 469586 690614
rect 469822 690378 469854 690614
rect 469234 670614 469854 690378
rect 469234 670378 469266 670614
rect 469502 670378 469586 670614
rect 469822 670378 469854 670614
rect 469234 659500 469854 670378
rect 471794 705798 472414 705830
rect 471794 705562 471826 705798
rect 472062 705562 472146 705798
rect 472382 705562 472414 705798
rect 471794 705478 472414 705562
rect 471794 705242 471826 705478
rect 472062 705242 472146 705478
rect 472382 705242 472414 705478
rect 471794 693294 472414 705242
rect 471794 693058 471826 693294
rect 472062 693058 472146 693294
rect 472382 693058 472414 693294
rect 471794 673294 472414 693058
rect 471794 673058 471826 673294
rect 472062 673058 472146 673294
rect 472382 673058 472414 673294
rect 471794 659500 472414 673058
rect 472954 694274 473574 710042
rect 482954 711558 483574 711590
rect 482954 711322 482986 711558
rect 483222 711322 483306 711558
rect 483542 711322 483574 711558
rect 482954 711238 483574 711322
rect 482954 711002 482986 711238
rect 483222 711002 483306 711238
rect 483542 711002 483574 711238
rect 479234 709638 479854 709670
rect 479234 709402 479266 709638
rect 479502 709402 479586 709638
rect 479822 709402 479854 709638
rect 479234 709318 479854 709402
rect 479234 709082 479266 709318
rect 479502 709082 479586 709318
rect 479822 709082 479854 709318
rect 472954 694038 472986 694274
rect 473222 694038 473306 694274
rect 473542 694038 473574 694274
rect 472954 674274 473574 694038
rect 472954 674038 472986 674274
rect 473222 674038 473306 674274
rect 473542 674038 473574 674274
rect 472954 659500 473574 674038
rect 475514 707718 476134 707750
rect 475514 707482 475546 707718
rect 475782 707482 475866 707718
rect 476102 707482 476134 707718
rect 475514 707398 476134 707482
rect 475514 707162 475546 707398
rect 475782 707162 475866 707398
rect 476102 707162 476134 707398
rect 475514 696954 476134 707162
rect 475514 696718 475546 696954
rect 475782 696718 475866 696954
rect 476102 696718 476134 696954
rect 475514 676954 476134 696718
rect 475514 676718 475546 676954
rect 475782 676718 475866 676954
rect 476102 676718 476134 676954
rect 475514 659500 476134 676718
rect 479234 700614 479854 709082
rect 479234 700378 479266 700614
rect 479502 700378 479586 700614
rect 479822 700378 479854 700614
rect 479234 680614 479854 700378
rect 479234 680378 479266 680614
rect 479502 680378 479586 680614
rect 479822 680378 479854 680614
rect 479234 660614 479854 680378
rect 479234 660378 479266 660614
rect 479502 660378 479586 660614
rect 479822 660378 479854 660614
rect 479234 659500 479854 660378
rect 481794 704838 482414 705830
rect 481794 704602 481826 704838
rect 482062 704602 482146 704838
rect 482382 704602 482414 704838
rect 481794 704518 482414 704602
rect 481794 704282 481826 704518
rect 482062 704282 482146 704518
rect 482382 704282 482414 704518
rect 481794 683294 482414 704282
rect 481794 683058 481826 683294
rect 482062 683058 482146 683294
rect 482382 683058 482414 683294
rect 481794 663294 482414 683058
rect 481794 663058 481826 663294
rect 482062 663058 482146 663294
rect 482382 663058 482414 663294
rect 481794 659500 482414 663058
rect 482954 684274 483574 711002
rect 492954 710598 493574 711590
rect 492954 710362 492986 710598
rect 493222 710362 493306 710598
rect 493542 710362 493574 710598
rect 492954 710278 493574 710362
rect 492954 710042 492986 710278
rect 493222 710042 493306 710278
rect 493542 710042 493574 710278
rect 489234 708678 489854 709670
rect 489234 708442 489266 708678
rect 489502 708442 489586 708678
rect 489822 708442 489854 708678
rect 489234 708358 489854 708442
rect 489234 708122 489266 708358
rect 489502 708122 489586 708358
rect 489822 708122 489854 708358
rect 482954 684038 482986 684274
rect 483222 684038 483306 684274
rect 483542 684038 483574 684274
rect 482954 664274 483574 684038
rect 482954 664038 482986 664274
rect 483222 664038 483306 664274
rect 483542 664038 483574 664274
rect 482954 659500 483574 664038
rect 485514 706758 486134 707750
rect 485514 706522 485546 706758
rect 485782 706522 485866 706758
rect 486102 706522 486134 706758
rect 485514 706438 486134 706522
rect 485514 706202 485546 706438
rect 485782 706202 485866 706438
rect 486102 706202 486134 706438
rect 485514 686954 486134 706202
rect 485514 686718 485546 686954
rect 485782 686718 485866 686954
rect 486102 686718 486134 686954
rect 485514 666954 486134 686718
rect 485514 666718 485546 666954
rect 485782 666718 485866 666954
rect 486102 666718 486134 666954
rect 485514 659500 486134 666718
rect 489234 690614 489854 708122
rect 489234 690378 489266 690614
rect 489502 690378 489586 690614
rect 489822 690378 489854 690614
rect 489234 670614 489854 690378
rect 489234 670378 489266 670614
rect 489502 670378 489586 670614
rect 489822 670378 489854 670614
rect 488947 659700 489013 659701
rect 488947 659636 488948 659700
rect 489012 659636 489013 659700
rect 488947 659635 489013 659636
rect 488950 657930 489010 659635
rect 489234 659500 489854 670378
rect 491794 705798 492414 705830
rect 491794 705562 491826 705798
rect 492062 705562 492146 705798
rect 492382 705562 492414 705798
rect 491794 705478 492414 705562
rect 491794 705242 491826 705478
rect 492062 705242 492146 705478
rect 492382 705242 492414 705478
rect 491794 693294 492414 705242
rect 491794 693058 491826 693294
rect 492062 693058 492146 693294
rect 492382 693058 492414 693294
rect 491794 673294 492414 693058
rect 491794 673058 491826 673294
rect 492062 673058 492146 673294
rect 492382 673058 492414 673294
rect 491794 659500 492414 673058
rect 492954 694274 493574 710042
rect 502954 711558 503574 711590
rect 502954 711322 502986 711558
rect 503222 711322 503306 711558
rect 503542 711322 503574 711558
rect 502954 711238 503574 711322
rect 502954 711002 502986 711238
rect 503222 711002 503306 711238
rect 503542 711002 503574 711238
rect 499234 709638 499854 709670
rect 499234 709402 499266 709638
rect 499502 709402 499586 709638
rect 499822 709402 499854 709638
rect 499234 709318 499854 709402
rect 499234 709082 499266 709318
rect 499502 709082 499586 709318
rect 499822 709082 499854 709318
rect 492954 694038 492986 694274
rect 493222 694038 493306 694274
rect 493542 694038 493574 694274
rect 492954 674274 493574 694038
rect 492954 674038 492986 674274
rect 493222 674038 493306 674274
rect 493542 674038 493574 674274
rect 492954 659500 493574 674038
rect 495514 707718 496134 707750
rect 495514 707482 495546 707718
rect 495782 707482 495866 707718
rect 496102 707482 496134 707718
rect 495514 707398 496134 707482
rect 495514 707162 495546 707398
rect 495782 707162 495866 707398
rect 496102 707162 496134 707398
rect 495514 696954 496134 707162
rect 495514 696718 495546 696954
rect 495782 696718 495866 696954
rect 496102 696718 496134 696954
rect 495514 676954 496134 696718
rect 495514 676718 495546 676954
rect 495782 676718 495866 676954
rect 496102 676718 496134 676954
rect 495514 659500 496134 676718
rect 499234 700614 499854 709082
rect 499234 700378 499266 700614
rect 499502 700378 499586 700614
rect 499822 700378 499854 700614
rect 499234 680614 499854 700378
rect 499234 680378 499266 680614
rect 499502 680378 499586 680614
rect 499822 680378 499854 680614
rect 499234 660614 499854 680378
rect 499234 660378 499266 660614
rect 499502 660378 499586 660614
rect 499822 660378 499854 660614
rect 499234 659500 499854 660378
rect 501794 704838 502414 705830
rect 501794 704602 501826 704838
rect 502062 704602 502146 704838
rect 502382 704602 502414 704838
rect 501794 704518 502414 704602
rect 501794 704282 501826 704518
rect 502062 704282 502146 704518
rect 502382 704282 502414 704518
rect 501794 683294 502414 704282
rect 501794 683058 501826 683294
rect 502062 683058 502146 683294
rect 502382 683058 502414 683294
rect 501794 663294 502414 683058
rect 501794 663058 501826 663294
rect 502062 663058 502146 663294
rect 502382 663058 502414 663294
rect 499987 659700 500053 659701
rect 499987 659636 499988 659700
rect 500052 659636 500053 659700
rect 499987 659635 500053 659636
rect 499990 657930 500050 659635
rect 501794 659500 502414 663058
rect 502954 684274 503574 711002
rect 512954 710598 513574 711590
rect 512954 710362 512986 710598
rect 513222 710362 513306 710598
rect 513542 710362 513574 710598
rect 512954 710278 513574 710362
rect 512954 710042 512986 710278
rect 513222 710042 513306 710278
rect 513542 710042 513574 710278
rect 509234 708678 509854 709670
rect 509234 708442 509266 708678
rect 509502 708442 509586 708678
rect 509822 708442 509854 708678
rect 509234 708358 509854 708442
rect 509234 708122 509266 708358
rect 509502 708122 509586 708358
rect 509822 708122 509854 708358
rect 502954 684038 502986 684274
rect 503222 684038 503306 684274
rect 503542 684038 503574 684274
rect 502954 664274 503574 684038
rect 502954 664038 502986 664274
rect 503222 664038 503306 664274
rect 503542 664038 503574 664274
rect 502954 659500 503574 664038
rect 505514 706758 506134 707750
rect 505514 706522 505546 706758
rect 505782 706522 505866 706758
rect 506102 706522 506134 706758
rect 505514 706438 506134 706522
rect 505514 706202 505546 706438
rect 505782 706202 505866 706438
rect 506102 706202 506134 706438
rect 505514 686954 506134 706202
rect 505514 686718 505546 686954
rect 505782 686718 505866 686954
rect 506102 686718 506134 686954
rect 505514 666954 506134 686718
rect 505514 666718 505546 666954
rect 505782 666718 505866 666954
rect 506102 666718 506134 666954
rect 505514 659500 506134 666718
rect 509234 690614 509854 708122
rect 509234 690378 509266 690614
rect 509502 690378 509586 690614
rect 509822 690378 509854 690614
rect 509234 670614 509854 690378
rect 509234 670378 509266 670614
rect 509502 670378 509586 670614
rect 509822 670378 509854 670614
rect 488950 657870 489492 657930
rect 499990 657870 500100 657930
rect 489432 657394 489492 657870
rect 500040 657394 500100 657870
rect 410272 653294 410620 653456
rect 410272 653058 410328 653294
rect 410564 653058 410620 653294
rect 410272 652896 410620 653058
rect 505336 653294 505684 653456
rect 505336 653058 505392 653294
rect 505628 653058 505684 653294
rect 505336 652896 505684 653058
rect 405514 646718 405546 646954
rect 405782 646718 405866 646954
rect 406102 646718 406134 646954
rect 405514 626954 406134 646718
rect 509234 650614 509854 670378
rect 509234 650378 509266 650614
rect 509502 650378 509586 650614
rect 509822 650378 509854 650614
rect 410952 643294 411300 643456
rect 410952 643058 411008 643294
rect 411244 643058 411300 643294
rect 410952 642896 411300 643058
rect 504656 643294 505004 643456
rect 504656 643058 504712 643294
rect 504948 643058 505004 643294
rect 504656 642896 505004 643058
rect 410272 633294 410620 633456
rect 410272 633058 410328 633294
rect 410564 633058 410620 633294
rect 410272 632896 410620 633058
rect 505336 633294 505684 633456
rect 505336 633058 505392 633294
rect 505628 633058 505684 633294
rect 505336 632896 505684 633058
rect 405514 626718 405546 626954
rect 405782 626718 405866 626954
rect 406102 626718 406134 626954
rect 405514 606954 406134 626718
rect 509234 630614 509854 650378
rect 509234 630378 509266 630614
rect 509502 630378 509586 630614
rect 509822 630378 509854 630614
rect 410952 623294 411300 623456
rect 410952 623058 411008 623294
rect 411244 623058 411300 623294
rect 410952 622896 411300 623058
rect 504656 623294 505004 623456
rect 504656 623058 504712 623294
rect 504948 623058 505004 623294
rect 504656 622896 505004 623058
rect 410272 613294 410620 613456
rect 410272 613058 410328 613294
rect 410564 613058 410620 613294
rect 410272 612896 410620 613058
rect 505336 613294 505684 613456
rect 505336 613058 505392 613294
rect 505628 613058 505684 613294
rect 505336 612896 505684 613058
rect 405514 606718 405546 606954
rect 405782 606718 405866 606954
rect 406102 606718 406134 606954
rect 405514 586954 406134 606718
rect 509234 610614 509854 630378
rect 509234 610378 509266 610614
rect 509502 610378 509586 610614
rect 509822 610378 509854 610614
rect 410952 603294 411300 603456
rect 410952 603058 411008 603294
rect 411244 603058 411300 603294
rect 410952 602896 411300 603058
rect 504656 603294 505004 603456
rect 504656 603058 504712 603294
rect 504948 603058 505004 603294
rect 504656 602896 505004 603058
rect 410272 593294 410620 593456
rect 410272 593058 410328 593294
rect 410564 593058 410620 593294
rect 410272 592896 410620 593058
rect 505336 593294 505684 593456
rect 505336 593058 505392 593294
rect 505628 593058 505684 593294
rect 505336 592896 505684 593058
rect 405514 586718 405546 586954
rect 405782 586718 405866 586954
rect 406102 586718 406134 586954
rect 405514 566954 406134 586718
rect 509234 590614 509854 610378
rect 509234 590378 509266 590614
rect 509502 590378 509586 590614
rect 509822 590378 509854 590614
rect 410952 583294 411300 583456
rect 410952 583058 411008 583294
rect 411244 583058 411300 583294
rect 410952 582896 411300 583058
rect 504656 583294 505004 583456
rect 504656 583058 504712 583294
rect 504948 583058 505004 583294
rect 504656 582896 505004 583058
rect 415856 577690 415916 578000
rect 425512 577690 425572 578000
rect 415534 577630 415916 577690
rect 425286 577630 425572 577690
rect 426736 577690 426796 578000
rect 427824 577690 427884 578000
rect 429184 577690 429244 578000
rect 430136 577690 430196 578000
rect 431360 577690 431420 578000
rect 426736 577630 430196 577690
rect 431358 577630 431420 577690
rect 432584 577690 432644 578000
rect 433672 577690 433732 578000
rect 435032 577690 435092 578000
rect 432584 577630 432706 577690
rect 433672 577630 433810 577690
rect 415534 576870 415594 577630
rect 415350 576810 415594 576870
rect 405514 566718 405546 566954
rect 405782 566718 405866 566954
rect 406102 566718 406134 566954
rect 405514 546954 406134 566718
rect 405514 546718 405546 546954
rect 405782 546718 405866 546954
rect 406102 546718 406134 546954
rect 405514 526954 406134 546718
rect 409234 570614 409854 576000
rect 409234 570378 409266 570614
rect 409502 570378 409586 570614
rect 409822 570378 409854 570614
rect 409234 550614 409854 570378
rect 409234 550378 409266 550614
rect 409502 550378 409586 550614
rect 409822 550378 409854 550614
rect 409234 539308 409854 550378
rect 411794 573294 412414 576000
rect 411794 573058 411826 573294
rect 412062 573058 412146 573294
rect 412382 573058 412414 573294
rect 411794 553294 412414 573058
rect 411794 553058 411826 553294
rect 412062 553058 412146 553294
rect 412382 553058 412414 553294
rect 411794 539308 412414 553058
rect 412954 574274 413574 576000
rect 415350 575381 415410 576810
rect 415347 575380 415413 575381
rect 415347 575316 415348 575380
rect 415412 575316 415413 575380
rect 415347 575315 415413 575316
rect 412954 574038 412986 574274
rect 413222 574038 413306 574274
rect 413542 574038 413574 574274
rect 412954 554274 413574 574038
rect 412954 554038 412986 554274
rect 413222 554038 413306 554274
rect 413542 554038 413574 554274
rect 412954 539308 413574 554038
rect 415514 556954 416134 576000
rect 415514 556718 415546 556954
rect 415782 556718 415866 556954
rect 416102 556718 416134 556954
rect 415514 539308 416134 556718
rect 419234 560614 419854 576000
rect 419234 560378 419266 560614
rect 419502 560378 419586 560614
rect 419822 560378 419854 560614
rect 419234 540614 419854 560378
rect 419234 540378 419266 540614
rect 419502 540378 419586 540614
rect 419822 540378 419854 540614
rect 419234 539308 419854 540378
rect 421794 563294 422414 576000
rect 421794 563058 421826 563294
rect 422062 563058 422146 563294
rect 422382 563058 422414 563294
rect 421794 543294 422414 563058
rect 421794 543058 421826 543294
rect 422062 543058 422146 543294
rect 422382 543058 422414 543294
rect 421794 539308 422414 543058
rect 422954 564274 423574 576000
rect 425286 575381 425346 577630
rect 425283 575380 425349 575381
rect 425283 575316 425284 575380
rect 425348 575316 425349 575380
rect 425283 575315 425349 575316
rect 422954 564038 422986 564274
rect 423222 564038 423306 564274
rect 423542 564038 423574 564274
rect 422954 544274 423574 564038
rect 422954 544038 422986 544274
rect 423222 544038 423306 544274
rect 423542 544038 423574 544274
rect 422954 539308 423574 544038
rect 425514 566954 426134 576000
rect 426758 575245 426818 577630
rect 426755 575244 426821 575245
rect 426755 575180 426756 575244
rect 426820 575180 426821 575244
rect 426755 575179 426821 575180
rect 425514 566718 425546 566954
rect 425782 566718 425866 566954
rect 426102 566718 426134 566954
rect 425514 546954 426134 566718
rect 425514 546718 425546 546954
rect 425782 546718 425866 546954
rect 426102 546718 426134 546954
rect 425514 539308 426134 546718
rect 429234 570614 429854 576000
rect 431358 574973 431418 577630
rect 431355 574972 431421 574973
rect 431355 574908 431356 574972
rect 431420 574908 431421 574972
rect 431355 574907 431421 574908
rect 429234 570378 429266 570614
rect 429502 570378 429586 570614
rect 429822 570378 429854 570614
rect 429234 550614 429854 570378
rect 429234 550378 429266 550614
rect 429502 550378 429586 550614
rect 429822 550378 429854 550614
rect 429234 539308 429854 550378
rect 431794 573294 432414 576000
rect 432646 574837 432706 577630
rect 432643 574836 432709 574837
rect 432643 574772 432644 574836
rect 432708 574772 432709 574836
rect 432643 574771 432709 574772
rect 431794 573058 431826 573294
rect 432062 573058 432146 573294
rect 432382 573058 432414 573294
rect 431794 553294 432414 573058
rect 431794 553058 431826 553294
rect 432062 553058 432146 553294
rect 432382 553058 432414 553294
rect 431794 539308 432414 553058
rect 432954 574274 433574 576000
rect 433750 574429 433810 577630
rect 434854 577630 435092 577690
rect 436120 577690 436180 578000
rect 437208 577690 437268 578000
rect 437888 577690 437948 578000
rect 436120 577630 436386 577690
rect 437208 577630 437306 577690
rect 433747 574428 433813 574429
rect 433747 574364 433748 574428
rect 433812 574364 433813 574428
rect 433747 574363 433813 574364
rect 432954 574038 432986 574274
rect 433222 574038 433306 574274
rect 433542 574038 433574 574274
rect 434854 574157 434914 577630
rect 434851 574156 434917 574157
rect 434851 574092 434852 574156
rect 434916 574092 434917 574156
rect 434851 574091 434917 574092
rect 432954 554274 433574 574038
rect 432954 554038 432986 554274
rect 433222 554038 433306 554274
rect 433542 554038 433574 554274
rect 432954 539308 433574 554038
rect 435514 556954 436134 576000
rect 436326 574293 436386 577630
rect 436323 574292 436389 574293
rect 436323 574228 436324 574292
rect 436388 574228 436389 574292
rect 436323 574227 436389 574228
rect 437246 574157 437306 577630
rect 437798 577630 437948 577690
rect 438296 577690 438356 578000
rect 439248 577690 439308 578000
rect 438296 577630 438410 577690
rect 437798 574157 437858 577630
rect 438350 575245 438410 577630
rect 439086 577630 439308 577690
rect 439656 577690 439716 578000
rect 440336 577690 440396 578000
rect 440744 577690 440804 578000
rect 439656 577630 440066 577690
rect 440336 577630 440434 577690
rect 438347 575244 438413 575245
rect 438347 575180 438348 575244
rect 438412 575180 438413 575244
rect 438347 575179 438413 575180
rect 439086 574157 439146 577630
rect 437243 574156 437309 574157
rect 437243 574092 437244 574156
rect 437308 574092 437309 574156
rect 437243 574091 437309 574092
rect 437795 574156 437861 574157
rect 437795 574092 437796 574156
rect 437860 574092 437861 574156
rect 437795 574091 437861 574092
rect 439083 574156 439149 574157
rect 439083 574092 439084 574156
rect 439148 574092 439149 574156
rect 439083 574091 439149 574092
rect 435514 556718 435546 556954
rect 435782 556718 435866 556954
rect 436102 556718 436134 556954
rect 435514 539308 436134 556718
rect 439234 560614 439854 576000
rect 440006 574837 440066 577630
rect 440003 574836 440069 574837
rect 440003 574772 440004 574836
rect 440068 574772 440069 574836
rect 440003 574771 440069 574772
rect 440374 574157 440434 577630
rect 440742 577630 440804 577690
rect 441832 577690 441892 578000
rect 441968 577690 442028 578000
rect 443056 577690 443116 578000
rect 441832 577630 441906 577690
rect 441968 577630 442090 577690
rect 440742 574293 440802 577630
rect 441846 577013 441906 577630
rect 441843 577012 441909 577013
rect 441843 576948 441844 577012
rect 441908 576948 441909 577012
rect 441843 576947 441909 576948
rect 442030 576870 442090 577630
rect 442950 577630 443116 577690
rect 443192 577690 443252 578000
rect 444144 577690 444204 578000
rect 443192 577630 443746 577690
rect 442030 576810 442642 576870
rect 440739 574292 440805 574293
rect 440739 574228 440740 574292
rect 440804 574228 440805 574292
rect 440739 574227 440805 574228
rect 440371 574156 440437 574157
rect 440371 574092 440372 574156
rect 440436 574092 440437 574156
rect 440371 574091 440437 574092
rect 439234 560378 439266 560614
rect 439502 560378 439586 560614
rect 439822 560378 439854 560614
rect 439234 540614 439854 560378
rect 439234 540378 439266 540614
rect 439502 540378 439586 540614
rect 439822 540378 439854 540614
rect 439234 539308 439854 540378
rect 441794 563294 442414 576000
rect 442582 574157 442642 576810
rect 442950 576330 443010 577630
rect 442766 576270 443010 576330
rect 442766 575109 442826 576270
rect 442763 575108 442829 575109
rect 442763 575044 442764 575108
rect 442828 575044 442829 575108
rect 442763 575043 442829 575044
rect 442579 574156 442645 574157
rect 442579 574092 442580 574156
rect 442644 574092 442645 574156
rect 442579 574091 442645 574092
rect 441794 563058 441826 563294
rect 442062 563058 442146 563294
rect 442382 563058 442414 563294
rect 441794 543294 442414 563058
rect 441794 543058 441826 543294
rect 442062 543058 442146 543294
rect 442382 543058 442414 543294
rect 441794 539308 442414 543058
rect 442954 564274 443574 576000
rect 443686 574157 443746 577630
rect 444054 577630 444204 577690
rect 444416 577690 444476 578000
rect 445504 577829 445564 578000
rect 445155 577828 445221 577829
rect 445155 577764 445156 577828
rect 445220 577764 445221 577828
rect 445155 577763 445221 577764
rect 445501 577828 445567 577829
rect 445501 577764 445502 577828
rect 445566 577764 445567 577828
rect 445501 577763 445567 577764
rect 444416 577630 444482 577690
rect 444054 574293 444114 577630
rect 444051 574292 444117 574293
rect 444051 574228 444052 574292
rect 444116 574228 444117 574292
rect 444051 574227 444117 574228
rect 444422 574157 444482 577630
rect 445158 574837 445218 577763
rect 445640 577690 445700 578000
rect 445342 577630 445700 577690
rect 446592 577690 446652 578000
rect 446864 577690 446924 578000
rect 447680 577690 447740 578000
rect 446592 577630 446690 577690
rect 445155 574836 445221 574837
rect 445155 574772 445156 574836
rect 445220 574772 445221 574836
rect 445155 574771 445221 574772
rect 445342 574293 445402 577630
rect 445339 574292 445405 574293
rect 445339 574228 445340 574292
rect 445404 574228 445405 574292
rect 445339 574227 445405 574228
rect 443683 574156 443749 574157
rect 443683 574092 443684 574156
rect 443748 574092 443749 574156
rect 443683 574091 443749 574092
rect 444419 574156 444485 574157
rect 444419 574092 444420 574156
rect 444484 574092 444485 574156
rect 444419 574091 444485 574092
rect 442954 564038 442986 564274
rect 443222 564038 443306 564274
rect 443542 564038 443574 564274
rect 442954 544274 443574 564038
rect 442954 544038 442986 544274
rect 443222 544038 443306 544274
rect 443542 544038 443574 544274
rect 442954 539308 443574 544038
rect 445514 566954 446134 576000
rect 446630 574293 446690 577630
rect 446814 577630 446924 577690
rect 447550 577630 447740 577690
rect 447816 577690 447876 578000
rect 448904 577690 448964 578000
rect 449312 577690 449372 578000
rect 447816 577630 447978 577690
rect 446627 574292 446693 574293
rect 446627 574228 446628 574292
rect 446692 574228 446693 574292
rect 446627 574227 446693 574228
rect 446814 574157 446874 577630
rect 447550 574293 447610 577630
rect 447547 574292 447613 574293
rect 447547 574228 447548 574292
rect 447612 574228 447613 574292
rect 447547 574227 447613 574228
rect 447918 574157 447978 577630
rect 448838 577630 448964 577690
rect 449206 577630 449372 577690
rect 450264 577690 450324 578000
rect 450672 577690 450732 578000
rect 451352 577690 451412 578000
rect 451896 577690 451956 578000
rect 450264 577630 450370 577690
rect 450672 577630 450738 577690
rect 451352 577630 451474 577690
rect 448838 575109 448898 577630
rect 449206 576870 449266 577630
rect 449022 576810 449266 576870
rect 448835 575108 448901 575109
rect 448835 575044 448836 575108
rect 448900 575044 448901 575108
rect 448835 575043 448901 575044
rect 449022 574157 449082 576810
rect 446811 574156 446877 574157
rect 446811 574092 446812 574156
rect 446876 574092 446877 574156
rect 446811 574091 446877 574092
rect 447915 574156 447981 574157
rect 447915 574092 447916 574156
rect 447980 574092 447981 574156
rect 447915 574091 447981 574092
rect 449019 574156 449085 574157
rect 449019 574092 449020 574156
rect 449084 574092 449085 574156
rect 449019 574091 449085 574092
rect 445514 566718 445546 566954
rect 445782 566718 445866 566954
rect 446102 566718 446134 566954
rect 445514 546954 446134 566718
rect 445514 546718 445546 546954
rect 445782 546718 445866 546954
rect 446102 546718 446134 546954
rect 445514 539308 446134 546718
rect 449234 570614 449854 576000
rect 450310 574293 450370 577630
rect 450307 574292 450373 574293
rect 450307 574228 450308 574292
rect 450372 574228 450373 574292
rect 450307 574227 450373 574228
rect 450678 574157 450738 577630
rect 451414 574565 451474 577630
rect 451598 577630 451956 577690
rect 452440 577690 452500 578000
rect 453120 577690 453180 578000
rect 452440 577630 452578 577690
rect 451411 574564 451477 574565
rect 451411 574500 451412 574564
rect 451476 574500 451477 574564
rect 451411 574499 451477 574500
rect 451598 574157 451658 577630
rect 450675 574156 450741 574157
rect 450675 574092 450676 574156
rect 450740 574092 450741 574156
rect 450675 574091 450741 574092
rect 451595 574156 451661 574157
rect 451595 574092 451596 574156
rect 451660 574092 451661 574156
rect 451595 574091 451661 574092
rect 449234 570378 449266 570614
rect 449502 570378 449586 570614
rect 449822 570378 449854 570614
rect 449234 550614 449854 570378
rect 449234 550378 449266 550614
rect 449502 550378 449586 550614
rect 449822 550378 449854 550614
rect 449234 539308 449854 550378
rect 451794 573294 452414 576000
rect 452518 574701 452578 577630
rect 452702 577630 453180 577690
rect 453528 577690 453588 578000
rect 454344 577690 454404 578000
rect 454888 577690 454948 578000
rect 455568 577690 455628 578000
rect 453528 577630 453866 577690
rect 454344 577630 454418 577690
rect 454888 577630 454970 577690
rect 452515 574700 452581 574701
rect 452515 574636 452516 574700
rect 452580 574636 452581 574700
rect 452515 574635 452581 574636
rect 452702 574293 452762 577630
rect 452699 574292 452765 574293
rect 452699 574228 452700 574292
rect 452764 574228 452765 574292
rect 452699 574227 452765 574228
rect 452954 574274 453574 576000
rect 451794 573058 451826 573294
rect 452062 573058 452146 573294
rect 452382 573058 452414 573294
rect 451794 553294 452414 573058
rect 451794 553058 451826 553294
rect 452062 553058 452146 553294
rect 452382 553058 452414 553294
rect 451794 539308 452414 553058
rect 452954 574038 452986 574274
rect 453222 574038 453306 574274
rect 453542 574038 453574 574274
rect 453806 574157 453866 577630
rect 454358 574157 454418 577630
rect 454910 574293 454970 577630
rect 455462 577630 455628 577690
rect 455976 577690 456036 578000
rect 456656 577690 456716 578000
rect 455976 577630 456442 577690
rect 455462 576197 455522 577630
rect 455459 576196 455525 576197
rect 455459 576132 455460 576196
rect 455524 576132 455525 576196
rect 455459 576131 455525 576132
rect 454907 574292 454973 574293
rect 454907 574228 454908 574292
rect 454972 574228 454973 574292
rect 454907 574227 454973 574228
rect 453803 574156 453869 574157
rect 453803 574092 453804 574156
rect 453868 574092 453869 574156
rect 453803 574091 453869 574092
rect 454355 574156 454421 574157
rect 454355 574092 454356 574156
rect 454420 574092 454421 574156
rect 454355 574091 454421 574092
rect 452954 554274 453574 574038
rect 452954 554038 452986 554274
rect 453222 554038 453306 554274
rect 453542 554038 453574 554274
rect 452954 539308 453574 554038
rect 455514 556954 456134 576000
rect 456382 574565 456442 577630
rect 456566 577630 456716 577690
rect 457064 577690 457124 578000
rect 457880 577690 457940 578000
rect 458288 577690 458348 578000
rect 459104 577690 459164 578000
rect 459376 577690 459436 578000
rect 457064 577630 457178 577690
rect 456379 574564 456445 574565
rect 456379 574500 456380 574564
rect 456444 574500 456445 574564
rect 456379 574499 456445 574500
rect 456566 574157 456626 577630
rect 457118 574293 457178 577630
rect 457854 577630 457940 577690
rect 458222 577630 458348 577690
rect 458958 577630 459164 577690
rect 459326 577630 459436 577690
rect 460600 577690 460660 578000
rect 460736 577690 460796 578000
rect 461416 577690 461476 578000
rect 461824 577690 461884 578000
rect 462912 577690 462972 578000
rect 460600 577630 460674 577690
rect 460736 577630 460858 577690
rect 457115 574292 457181 574293
rect 457115 574228 457116 574292
rect 457180 574228 457181 574292
rect 457115 574227 457181 574228
rect 457854 574157 457914 577630
rect 458222 574429 458282 577630
rect 458219 574428 458285 574429
rect 458219 574364 458220 574428
rect 458284 574364 458285 574428
rect 458219 574363 458285 574364
rect 458958 574157 459018 577630
rect 459326 576197 459386 577630
rect 459323 576196 459389 576197
rect 459323 576132 459324 576196
rect 459388 576132 459389 576196
rect 459323 576131 459389 576132
rect 456563 574156 456629 574157
rect 456563 574092 456564 574156
rect 456628 574092 456629 574156
rect 456563 574091 456629 574092
rect 457851 574156 457917 574157
rect 457851 574092 457852 574156
rect 457916 574092 457917 574156
rect 457851 574091 457917 574092
rect 458955 574156 459021 574157
rect 458955 574092 458956 574156
rect 459020 574092 459021 574156
rect 458955 574091 459021 574092
rect 455514 556718 455546 556954
rect 455782 556718 455866 556954
rect 456102 556718 456134 556954
rect 455514 539308 456134 556718
rect 459234 560614 459854 576000
rect 460614 574157 460674 577630
rect 460798 574429 460858 577630
rect 461350 577630 461476 577690
rect 461718 577630 461884 577690
rect 462822 577630 462972 577690
rect 463184 577690 463244 578000
rect 464000 577690 464060 578000
rect 464408 577690 464468 578000
rect 465224 577690 465284 578000
rect 465632 577690 465692 578000
rect 466584 577690 466644 578000
rect 463184 577630 463250 577690
rect 460795 574428 460861 574429
rect 460795 574364 460796 574428
rect 460860 574364 460861 574428
rect 460795 574363 460861 574364
rect 461350 574293 461410 577630
rect 461718 576870 461778 577630
rect 462822 577013 462882 577630
rect 462819 577012 462885 577013
rect 462819 576948 462820 577012
rect 462884 576948 462885 577012
rect 462819 576947 462885 576948
rect 463190 576870 463250 577630
rect 461534 576810 461778 576870
rect 462638 576810 463250 576870
rect 463926 577630 464060 577690
rect 464294 577630 464468 577690
rect 465030 577630 465284 577690
rect 465398 577630 465692 577690
rect 466502 577630 466644 577690
rect 466856 577690 466916 578000
rect 467672 577690 467732 578000
rect 466856 577630 466930 577690
rect 461347 574292 461413 574293
rect 461347 574228 461348 574292
rect 461412 574228 461413 574292
rect 461347 574227 461413 574228
rect 461534 574157 461594 576810
rect 460611 574156 460677 574157
rect 460611 574092 460612 574156
rect 460676 574092 460677 574156
rect 460611 574091 460677 574092
rect 461531 574156 461597 574157
rect 461531 574092 461532 574156
rect 461596 574092 461597 574156
rect 461531 574091 461597 574092
rect 459234 560378 459266 560614
rect 459502 560378 459586 560614
rect 459822 560378 459854 560614
rect 459234 540614 459854 560378
rect 459234 540378 459266 540614
rect 459502 540378 459586 540614
rect 459822 540378 459854 540614
rect 459234 539308 459854 540378
rect 461794 563294 462414 576000
rect 462638 574157 462698 576810
rect 462635 574156 462701 574157
rect 462635 574092 462636 574156
rect 462700 574092 462701 574156
rect 462635 574091 462701 574092
rect 461794 563058 461826 563294
rect 462062 563058 462146 563294
rect 462382 563058 462414 563294
rect 461794 543294 462414 563058
rect 461794 543058 461826 543294
rect 462062 543058 462146 543294
rect 462382 543058 462414 543294
rect 461794 539308 462414 543058
rect 462954 564274 463574 576000
rect 463926 574565 463986 577630
rect 463923 574564 463989 574565
rect 463923 574500 463924 574564
rect 463988 574500 463989 574564
rect 463923 574499 463989 574500
rect 464294 574157 464354 577630
rect 465030 574429 465090 577630
rect 465398 576870 465458 577630
rect 465214 576810 465458 576870
rect 465027 574428 465093 574429
rect 465027 574364 465028 574428
rect 465092 574364 465093 574428
rect 465027 574363 465093 574364
rect 465214 574293 465274 576810
rect 465211 574292 465277 574293
rect 465211 574228 465212 574292
rect 465276 574228 465277 574292
rect 465211 574227 465277 574228
rect 464291 574156 464357 574157
rect 464291 574092 464292 574156
rect 464356 574092 464357 574156
rect 464291 574091 464357 574092
rect 462954 564038 462986 564274
rect 463222 564038 463306 564274
rect 463542 564038 463574 564274
rect 462954 544274 463574 564038
rect 462954 544038 462986 544274
rect 463222 544038 463306 544274
rect 463542 544038 463574 544274
rect 462954 539308 463574 544038
rect 465514 566954 466134 576000
rect 466502 574157 466562 577630
rect 466870 574157 466930 577630
rect 467606 577630 467732 577690
rect 467606 575245 467666 577630
rect 467808 577010 467868 578000
rect 469304 577690 469364 578000
rect 467790 576950 467868 577010
rect 469262 577630 469364 577690
rect 470528 577690 470588 578000
rect 471888 577690 471948 578000
rect 473112 577690 473172 578000
rect 474336 577690 474396 578000
rect 475560 577690 475620 578000
rect 470528 577630 470794 577690
rect 467603 575244 467669 575245
rect 467603 575180 467604 575244
rect 467668 575180 467669 575244
rect 467603 575179 467669 575180
rect 467790 574157 467850 576950
rect 469262 576197 469322 577630
rect 470734 576870 470794 577630
rect 470366 576810 470794 576870
rect 471470 577630 471948 577690
rect 472758 577630 473172 577690
rect 474230 577630 474396 577690
rect 475334 577630 475620 577690
rect 476784 577690 476844 578000
rect 492696 577829 492756 578000
rect 492693 577828 492759 577829
rect 492693 577764 492694 577828
rect 492758 577764 492759 577828
rect 492693 577763 492759 577764
rect 492627 577692 492693 577693
rect 476784 577630 476866 577690
rect 469259 576196 469325 576197
rect 469259 576132 469260 576196
rect 469324 576132 469325 576196
rect 469259 576131 469325 576132
rect 466499 574156 466565 574157
rect 466499 574092 466500 574156
rect 466564 574092 466565 574156
rect 466499 574091 466565 574092
rect 466867 574156 466933 574157
rect 466867 574092 466868 574156
rect 466932 574092 466933 574156
rect 466867 574091 466933 574092
rect 467787 574156 467853 574157
rect 467787 574092 467788 574156
rect 467852 574092 467853 574156
rect 467787 574091 467853 574092
rect 465514 566718 465546 566954
rect 465782 566718 465866 566954
rect 466102 566718 466134 566954
rect 465514 546954 466134 566718
rect 465514 546718 465546 546954
rect 465782 546718 465866 546954
rect 466102 546718 466134 546954
rect 465514 539308 466134 546718
rect 469234 570614 469854 576000
rect 470366 574154 470426 576810
rect 471470 574293 471530 577630
rect 471467 574292 471533 574293
rect 471467 574228 471468 574292
rect 471532 574228 471533 574292
rect 471467 574227 471533 574228
rect 470547 574156 470613 574157
rect 470547 574154 470548 574156
rect 470366 574094 470548 574154
rect 470547 574092 470548 574094
rect 470612 574092 470613 574156
rect 470547 574091 470613 574092
rect 469234 570378 469266 570614
rect 469502 570378 469586 570614
rect 469822 570378 469854 570614
rect 469234 550614 469854 570378
rect 469234 550378 469266 550614
rect 469502 550378 469586 550614
rect 469822 550378 469854 550614
rect 469234 539308 469854 550378
rect 471794 573294 472414 576000
rect 472758 574157 472818 577630
rect 472954 574274 473574 576000
rect 472755 574156 472821 574157
rect 472755 574092 472756 574156
rect 472820 574092 472821 574156
rect 472755 574091 472821 574092
rect 471794 573058 471826 573294
rect 472062 573058 472146 573294
rect 472382 573058 472414 573294
rect 471794 553294 472414 573058
rect 471794 553058 471826 553294
rect 472062 553058 472146 553294
rect 472382 553058 472414 553294
rect 471794 539308 472414 553058
rect 472954 574038 472986 574274
rect 473222 574038 473306 574274
rect 473542 574038 473574 574274
rect 474230 574157 474290 577630
rect 475334 574157 475394 577630
rect 474227 574156 474293 574157
rect 474227 574092 474228 574156
rect 474292 574092 474293 574156
rect 474227 574091 474293 574092
rect 475331 574156 475397 574157
rect 475331 574092 475332 574156
rect 475396 574092 475397 574156
rect 475331 574091 475397 574092
rect 472954 554274 473574 574038
rect 472954 554038 472986 554274
rect 473222 554038 473306 554274
rect 473542 554038 473574 554274
rect 472954 539308 473574 554038
rect 475514 556954 476134 576000
rect 476806 574157 476866 577630
rect 492627 577628 492628 577692
rect 492692 577628 492693 577692
rect 492832 577690 492892 578000
rect 492627 577627 492693 577628
rect 492814 577630 492892 577690
rect 492968 577690 493028 578000
rect 493104 577829 493164 578000
rect 493101 577828 493167 577829
rect 493101 577764 493102 577828
rect 493166 577764 493167 577828
rect 493101 577763 493167 577764
rect 492968 577630 493058 577690
rect 476803 574156 476869 574157
rect 476803 574092 476804 574156
rect 476868 574092 476869 574156
rect 476803 574091 476869 574092
rect 475514 556718 475546 556954
rect 475782 556718 475866 556954
rect 476102 556718 476134 556954
rect 475514 539308 476134 556718
rect 479234 560614 479854 576000
rect 479234 560378 479266 560614
rect 479502 560378 479586 560614
rect 479822 560378 479854 560614
rect 479234 540614 479854 560378
rect 479234 540378 479266 540614
rect 479502 540378 479586 540614
rect 479822 540378 479854 540614
rect 479234 539308 479854 540378
rect 481794 563294 482414 576000
rect 481794 563058 481826 563294
rect 482062 563058 482146 563294
rect 482382 563058 482414 563294
rect 481794 543294 482414 563058
rect 481794 543058 481826 543294
rect 482062 543058 482146 543294
rect 482382 543058 482414 543294
rect 481794 539308 482414 543058
rect 482954 564274 483574 576000
rect 482954 564038 482986 564274
rect 483222 564038 483306 564274
rect 483542 564038 483574 564274
rect 482954 544274 483574 564038
rect 482954 544038 482986 544274
rect 483222 544038 483306 544274
rect 483542 544038 483574 544274
rect 482954 539308 483574 544038
rect 485514 566954 486134 576000
rect 485514 566718 485546 566954
rect 485782 566718 485866 566954
rect 486102 566718 486134 566954
rect 485514 546954 486134 566718
rect 485514 546718 485546 546954
rect 485782 546718 485866 546954
rect 486102 546718 486134 546954
rect 485514 539308 486134 546718
rect 489234 570614 489854 576000
rect 489234 570378 489266 570614
rect 489502 570378 489586 570614
rect 489822 570378 489854 570614
rect 489234 550614 489854 570378
rect 489234 550378 489266 550614
rect 489502 550378 489586 550614
rect 489822 550378 489854 550614
rect 489234 539308 489854 550378
rect 491794 573294 492414 576000
rect 492630 574429 492690 577627
rect 492627 574428 492693 574429
rect 492627 574364 492628 574428
rect 492692 574364 492693 574428
rect 492627 574363 492693 574364
rect 492627 574292 492693 574293
rect 492627 574228 492628 574292
rect 492692 574290 492693 574292
rect 492814 574290 492874 577630
rect 492998 576877 493058 577630
rect 492995 576876 493061 576877
rect 492995 576812 492996 576876
rect 493060 576812 493061 576876
rect 492995 576811 493061 576812
rect 492692 574230 492874 574290
rect 492954 574274 493574 576000
rect 492692 574228 492693 574230
rect 492627 574227 492693 574228
rect 491794 573058 491826 573294
rect 492062 573058 492146 573294
rect 492382 573058 492414 573294
rect 491794 553294 492414 573058
rect 491794 553058 491826 553294
rect 492062 553058 492146 553294
rect 492382 553058 492414 553294
rect 491794 539308 492414 553058
rect 492954 574038 492986 574274
rect 493222 574038 493306 574274
rect 493542 574038 493574 574274
rect 492954 554274 493574 574038
rect 492954 554038 492986 554274
rect 493222 554038 493306 554274
rect 493542 554038 493574 554274
rect 492954 539308 493574 554038
rect 495514 556954 496134 576000
rect 495514 556718 495546 556954
rect 495782 556718 495866 556954
rect 496102 556718 496134 556954
rect 495514 539308 496134 556718
rect 499234 560614 499854 576000
rect 499234 560378 499266 560614
rect 499502 560378 499586 560614
rect 499822 560378 499854 560614
rect 499234 540614 499854 560378
rect 499234 540378 499266 540614
rect 499502 540378 499586 540614
rect 499822 540378 499854 540614
rect 499234 539308 499854 540378
rect 501794 563294 502414 576000
rect 501794 563058 501826 563294
rect 502062 563058 502146 563294
rect 502382 563058 502414 563294
rect 501794 543294 502414 563058
rect 501794 543058 501826 543294
rect 502062 543058 502146 543294
rect 502382 543058 502414 543294
rect 501794 539308 502414 543058
rect 502954 564274 503574 576000
rect 502954 564038 502986 564274
rect 503222 564038 503306 564274
rect 503542 564038 503574 564274
rect 502954 544274 503574 564038
rect 502954 544038 502986 544274
rect 503222 544038 503306 544274
rect 503542 544038 503574 544274
rect 502954 539308 503574 544038
rect 505514 566954 506134 576000
rect 505514 566718 505546 566954
rect 505782 566718 505866 566954
rect 506102 566718 506134 566954
rect 505514 546954 506134 566718
rect 505514 546718 505546 546954
rect 505782 546718 505866 546954
rect 506102 546718 506134 546954
rect 505514 539308 506134 546718
rect 509234 570614 509854 590378
rect 509234 570378 509266 570614
rect 509502 570378 509586 570614
rect 509822 570378 509854 570614
rect 509234 550614 509854 570378
rect 509234 550378 509266 550614
rect 509502 550378 509586 550614
rect 509822 550378 509854 550614
rect 509234 539308 509854 550378
rect 511794 705798 512414 705830
rect 511794 705562 511826 705798
rect 512062 705562 512146 705798
rect 512382 705562 512414 705798
rect 511794 705478 512414 705562
rect 511794 705242 511826 705478
rect 512062 705242 512146 705478
rect 512382 705242 512414 705478
rect 511794 693294 512414 705242
rect 511794 693058 511826 693294
rect 512062 693058 512146 693294
rect 512382 693058 512414 693294
rect 511794 673294 512414 693058
rect 511794 673058 511826 673294
rect 512062 673058 512146 673294
rect 512382 673058 512414 673294
rect 511794 653294 512414 673058
rect 511794 653058 511826 653294
rect 512062 653058 512146 653294
rect 512382 653058 512414 653294
rect 511794 633294 512414 653058
rect 511794 633058 511826 633294
rect 512062 633058 512146 633294
rect 512382 633058 512414 633294
rect 511794 613294 512414 633058
rect 511794 613058 511826 613294
rect 512062 613058 512146 613294
rect 512382 613058 512414 613294
rect 511794 593294 512414 613058
rect 511794 593058 511826 593294
rect 512062 593058 512146 593294
rect 512382 593058 512414 593294
rect 511794 573294 512414 593058
rect 511794 573058 511826 573294
rect 512062 573058 512146 573294
rect 512382 573058 512414 573294
rect 511794 553294 512414 573058
rect 511794 553058 511826 553294
rect 512062 553058 512146 553294
rect 512382 553058 512414 553294
rect 511794 539308 512414 553058
rect 512954 694274 513574 710042
rect 522954 711558 523574 711590
rect 522954 711322 522986 711558
rect 523222 711322 523306 711558
rect 523542 711322 523574 711558
rect 522954 711238 523574 711322
rect 522954 711002 522986 711238
rect 523222 711002 523306 711238
rect 523542 711002 523574 711238
rect 519234 709638 519854 709670
rect 519234 709402 519266 709638
rect 519502 709402 519586 709638
rect 519822 709402 519854 709638
rect 519234 709318 519854 709402
rect 519234 709082 519266 709318
rect 519502 709082 519586 709318
rect 519822 709082 519854 709318
rect 512954 694038 512986 694274
rect 513222 694038 513306 694274
rect 513542 694038 513574 694274
rect 512954 674274 513574 694038
rect 512954 674038 512986 674274
rect 513222 674038 513306 674274
rect 513542 674038 513574 674274
rect 512954 654274 513574 674038
rect 512954 654038 512986 654274
rect 513222 654038 513306 654274
rect 513542 654038 513574 654274
rect 512954 634274 513574 654038
rect 512954 634038 512986 634274
rect 513222 634038 513306 634274
rect 513542 634038 513574 634274
rect 512954 614274 513574 634038
rect 512954 614038 512986 614274
rect 513222 614038 513306 614274
rect 513542 614038 513574 614274
rect 512954 594274 513574 614038
rect 512954 594038 512986 594274
rect 513222 594038 513306 594274
rect 513542 594038 513574 594274
rect 512954 574274 513574 594038
rect 512954 574038 512986 574274
rect 513222 574038 513306 574274
rect 513542 574038 513574 574274
rect 512954 554274 513574 574038
rect 512954 554038 512986 554274
rect 513222 554038 513306 554274
rect 513542 554038 513574 554274
rect 512954 539308 513574 554038
rect 515514 707718 516134 707750
rect 515514 707482 515546 707718
rect 515782 707482 515866 707718
rect 516102 707482 516134 707718
rect 515514 707398 516134 707482
rect 515514 707162 515546 707398
rect 515782 707162 515866 707398
rect 516102 707162 516134 707398
rect 515514 696954 516134 707162
rect 515514 696718 515546 696954
rect 515782 696718 515866 696954
rect 516102 696718 516134 696954
rect 515514 676954 516134 696718
rect 515514 676718 515546 676954
rect 515782 676718 515866 676954
rect 516102 676718 516134 676954
rect 515514 656954 516134 676718
rect 515514 656718 515546 656954
rect 515782 656718 515866 656954
rect 516102 656718 516134 656954
rect 515514 636954 516134 656718
rect 515514 636718 515546 636954
rect 515782 636718 515866 636954
rect 516102 636718 516134 636954
rect 515514 616954 516134 636718
rect 515514 616718 515546 616954
rect 515782 616718 515866 616954
rect 516102 616718 516134 616954
rect 515514 596954 516134 616718
rect 515514 596718 515546 596954
rect 515782 596718 515866 596954
rect 516102 596718 516134 596954
rect 515514 576954 516134 596718
rect 515514 576718 515546 576954
rect 515782 576718 515866 576954
rect 516102 576718 516134 576954
rect 515514 556954 516134 576718
rect 515514 556718 515546 556954
rect 515782 556718 515866 556954
rect 516102 556718 516134 556954
rect 515514 539308 516134 556718
rect 519234 700614 519854 709082
rect 519234 700378 519266 700614
rect 519502 700378 519586 700614
rect 519822 700378 519854 700614
rect 519234 680614 519854 700378
rect 519234 680378 519266 680614
rect 519502 680378 519586 680614
rect 519822 680378 519854 680614
rect 519234 660614 519854 680378
rect 519234 660378 519266 660614
rect 519502 660378 519586 660614
rect 519822 660378 519854 660614
rect 519234 640614 519854 660378
rect 519234 640378 519266 640614
rect 519502 640378 519586 640614
rect 519822 640378 519854 640614
rect 519234 620614 519854 640378
rect 519234 620378 519266 620614
rect 519502 620378 519586 620614
rect 519822 620378 519854 620614
rect 519234 600614 519854 620378
rect 519234 600378 519266 600614
rect 519502 600378 519586 600614
rect 519822 600378 519854 600614
rect 519234 580614 519854 600378
rect 519234 580378 519266 580614
rect 519502 580378 519586 580614
rect 519822 580378 519854 580614
rect 519234 560614 519854 580378
rect 519234 560378 519266 560614
rect 519502 560378 519586 560614
rect 519822 560378 519854 560614
rect 519234 540614 519854 560378
rect 519234 540378 519266 540614
rect 519502 540378 519586 540614
rect 519822 540378 519854 540614
rect 519234 539308 519854 540378
rect 521794 704838 522414 705830
rect 521794 704602 521826 704838
rect 522062 704602 522146 704838
rect 522382 704602 522414 704838
rect 521794 704518 522414 704602
rect 521794 704282 521826 704518
rect 522062 704282 522146 704518
rect 522382 704282 522414 704518
rect 521794 683294 522414 704282
rect 521794 683058 521826 683294
rect 522062 683058 522146 683294
rect 522382 683058 522414 683294
rect 521794 663294 522414 683058
rect 521794 663058 521826 663294
rect 522062 663058 522146 663294
rect 522382 663058 522414 663294
rect 521794 643294 522414 663058
rect 521794 643058 521826 643294
rect 522062 643058 522146 643294
rect 522382 643058 522414 643294
rect 521794 623294 522414 643058
rect 521794 623058 521826 623294
rect 522062 623058 522146 623294
rect 522382 623058 522414 623294
rect 521794 603294 522414 623058
rect 521794 603058 521826 603294
rect 522062 603058 522146 603294
rect 522382 603058 522414 603294
rect 521794 583294 522414 603058
rect 521794 583058 521826 583294
rect 522062 583058 522146 583294
rect 522382 583058 522414 583294
rect 521794 563294 522414 583058
rect 521794 563058 521826 563294
rect 522062 563058 522146 563294
rect 522382 563058 522414 563294
rect 521794 543294 522414 563058
rect 521794 543058 521826 543294
rect 522062 543058 522146 543294
rect 522382 543058 522414 543294
rect 521794 539308 522414 543058
rect 522954 684274 523574 711002
rect 532954 710598 533574 711590
rect 532954 710362 532986 710598
rect 533222 710362 533306 710598
rect 533542 710362 533574 710598
rect 532954 710278 533574 710362
rect 532954 710042 532986 710278
rect 533222 710042 533306 710278
rect 533542 710042 533574 710278
rect 529234 708678 529854 709670
rect 529234 708442 529266 708678
rect 529502 708442 529586 708678
rect 529822 708442 529854 708678
rect 529234 708358 529854 708442
rect 529234 708122 529266 708358
rect 529502 708122 529586 708358
rect 529822 708122 529854 708358
rect 522954 684038 522986 684274
rect 523222 684038 523306 684274
rect 523542 684038 523574 684274
rect 522954 664274 523574 684038
rect 522954 664038 522986 664274
rect 523222 664038 523306 664274
rect 523542 664038 523574 664274
rect 522954 644274 523574 664038
rect 522954 644038 522986 644274
rect 523222 644038 523306 644274
rect 523542 644038 523574 644274
rect 522954 624274 523574 644038
rect 522954 624038 522986 624274
rect 523222 624038 523306 624274
rect 523542 624038 523574 624274
rect 522954 604274 523574 624038
rect 522954 604038 522986 604274
rect 523222 604038 523306 604274
rect 523542 604038 523574 604274
rect 522954 584274 523574 604038
rect 522954 584038 522986 584274
rect 523222 584038 523306 584274
rect 523542 584038 523574 584274
rect 522954 564274 523574 584038
rect 522954 564038 522986 564274
rect 523222 564038 523306 564274
rect 523542 564038 523574 564274
rect 522954 544274 523574 564038
rect 522954 544038 522986 544274
rect 523222 544038 523306 544274
rect 523542 544038 523574 544274
rect 522954 539308 523574 544038
rect 525514 706758 526134 707750
rect 525514 706522 525546 706758
rect 525782 706522 525866 706758
rect 526102 706522 526134 706758
rect 525514 706438 526134 706522
rect 525514 706202 525546 706438
rect 525782 706202 525866 706438
rect 526102 706202 526134 706438
rect 525514 686954 526134 706202
rect 525514 686718 525546 686954
rect 525782 686718 525866 686954
rect 526102 686718 526134 686954
rect 525514 666954 526134 686718
rect 525514 666718 525546 666954
rect 525782 666718 525866 666954
rect 526102 666718 526134 666954
rect 525514 646954 526134 666718
rect 525514 646718 525546 646954
rect 525782 646718 525866 646954
rect 526102 646718 526134 646954
rect 525514 626954 526134 646718
rect 525514 626718 525546 626954
rect 525782 626718 525866 626954
rect 526102 626718 526134 626954
rect 525514 606954 526134 626718
rect 525514 606718 525546 606954
rect 525782 606718 525866 606954
rect 526102 606718 526134 606954
rect 525514 586954 526134 606718
rect 525514 586718 525546 586954
rect 525782 586718 525866 586954
rect 526102 586718 526134 586954
rect 525514 566954 526134 586718
rect 525514 566718 525546 566954
rect 525782 566718 525866 566954
rect 526102 566718 526134 566954
rect 525514 546954 526134 566718
rect 525514 546718 525546 546954
rect 525782 546718 525866 546954
rect 526102 546718 526134 546954
rect 525514 539308 526134 546718
rect 529234 690614 529854 708122
rect 529234 690378 529266 690614
rect 529502 690378 529586 690614
rect 529822 690378 529854 690614
rect 529234 670614 529854 690378
rect 529234 670378 529266 670614
rect 529502 670378 529586 670614
rect 529822 670378 529854 670614
rect 529234 650614 529854 670378
rect 529234 650378 529266 650614
rect 529502 650378 529586 650614
rect 529822 650378 529854 650614
rect 529234 630614 529854 650378
rect 529234 630378 529266 630614
rect 529502 630378 529586 630614
rect 529822 630378 529854 630614
rect 529234 610614 529854 630378
rect 529234 610378 529266 610614
rect 529502 610378 529586 610614
rect 529822 610378 529854 610614
rect 529234 590614 529854 610378
rect 529234 590378 529266 590614
rect 529502 590378 529586 590614
rect 529822 590378 529854 590614
rect 529234 570614 529854 590378
rect 529234 570378 529266 570614
rect 529502 570378 529586 570614
rect 529822 570378 529854 570614
rect 529234 550614 529854 570378
rect 529234 550378 529266 550614
rect 529502 550378 529586 550614
rect 529822 550378 529854 550614
rect 528323 540292 528389 540293
rect 528323 540228 528324 540292
rect 528388 540228 528389 540292
rect 528323 540227 528389 540228
rect 528326 537570 528386 540227
rect 529059 539748 529125 539749
rect 529059 539684 529060 539748
rect 529124 539684 529125 539748
rect 529059 539683 529125 539684
rect 529062 538230 529122 539683
rect 529234 539308 529854 550378
rect 531794 705798 532414 705830
rect 531794 705562 531826 705798
rect 532062 705562 532146 705798
rect 532382 705562 532414 705798
rect 531794 705478 532414 705562
rect 531794 705242 531826 705478
rect 532062 705242 532146 705478
rect 532382 705242 532414 705478
rect 531794 693294 532414 705242
rect 531794 693058 531826 693294
rect 532062 693058 532146 693294
rect 532382 693058 532414 693294
rect 531794 673294 532414 693058
rect 531794 673058 531826 673294
rect 532062 673058 532146 673294
rect 532382 673058 532414 673294
rect 531794 653294 532414 673058
rect 531794 653058 531826 653294
rect 532062 653058 532146 653294
rect 532382 653058 532414 653294
rect 531794 633294 532414 653058
rect 531794 633058 531826 633294
rect 532062 633058 532146 633294
rect 532382 633058 532414 633294
rect 531794 613294 532414 633058
rect 531794 613058 531826 613294
rect 532062 613058 532146 613294
rect 532382 613058 532414 613294
rect 531794 593294 532414 613058
rect 531794 593058 531826 593294
rect 532062 593058 532146 593294
rect 532382 593058 532414 593294
rect 531794 573294 532414 593058
rect 531794 573058 531826 573294
rect 532062 573058 532146 573294
rect 532382 573058 532414 573294
rect 531794 553294 532414 573058
rect 531794 553058 531826 553294
rect 532062 553058 532146 553294
rect 532382 553058 532414 553294
rect 531794 539308 532414 553058
rect 532954 694274 533574 710042
rect 542954 711558 543574 711590
rect 542954 711322 542986 711558
rect 543222 711322 543306 711558
rect 543542 711322 543574 711558
rect 542954 711238 543574 711322
rect 542954 711002 542986 711238
rect 543222 711002 543306 711238
rect 543542 711002 543574 711238
rect 539234 709638 539854 709670
rect 539234 709402 539266 709638
rect 539502 709402 539586 709638
rect 539822 709402 539854 709638
rect 539234 709318 539854 709402
rect 539234 709082 539266 709318
rect 539502 709082 539586 709318
rect 539822 709082 539854 709318
rect 532954 694038 532986 694274
rect 533222 694038 533306 694274
rect 533542 694038 533574 694274
rect 532954 674274 533574 694038
rect 532954 674038 532986 674274
rect 533222 674038 533306 674274
rect 533542 674038 533574 674274
rect 532954 654274 533574 674038
rect 532954 654038 532986 654274
rect 533222 654038 533306 654274
rect 533542 654038 533574 654274
rect 532954 634274 533574 654038
rect 532954 634038 532986 634274
rect 533222 634038 533306 634274
rect 533542 634038 533574 634274
rect 532954 614274 533574 634038
rect 532954 614038 532986 614274
rect 533222 614038 533306 614274
rect 533542 614038 533574 614274
rect 532954 594274 533574 614038
rect 532954 594038 532986 594274
rect 533222 594038 533306 594274
rect 533542 594038 533574 594274
rect 532954 574274 533574 594038
rect 532954 574038 532986 574274
rect 533222 574038 533306 574274
rect 533542 574038 533574 574274
rect 532954 554274 533574 574038
rect 532954 554038 532986 554274
rect 533222 554038 533306 554274
rect 533542 554038 533574 554274
rect 532954 539308 533574 554038
rect 535514 707718 536134 707750
rect 535514 707482 535546 707718
rect 535782 707482 535866 707718
rect 536102 707482 536134 707718
rect 535514 707398 536134 707482
rect 535514 707162 535546 707398
rect 535782 707162 535866 707398
rect 536102 707162 536134 707398
rect 535514 696954 536134 707162
rect 535514 696718 535546 696954
rect 535782 696718 535866 696954
rect 536102 696718 536134 696954
rect 535514 676954 536134 696718
rect 535514 676718 535546 676954
rect 535782 676718 535866 676954
rect 536102 676718 536134 676954
rect 535514 656954 536134 676718
rect 535514 656718 535546 656954
rect 535782 656718 535866 656954
rect 536102 656718 536134 656954
rect 535514 636954 536134 656718
rect 535514 636718 535546 636954
rect 535782 636718 535866 636954
rect 536102 636718 536134 636954
rect 535514 616954 536134 636718
rect 535514 616718 535546 616954
rect 535782 616718 535866 616954
rect 536102 616718 536134 616954
rect 535514 596954 536134 616718
rect 535514 596718 535546 596954
rect 535782 596718 535866 596954
rect 536102 596718 536134 596954
rect 535514 576954 536134 596718
rect 535514 576718 535546 576954
rect 535782 576718 535866 576954
rect 536102 576718 536134 576954
rect 535514 556954 536134 576718
rect 535514 556718 535546 556954
rect 535782 556718 535866 556954
rect 536102 556718 536134 556954
rect 535514 539308 536134 556718
rect 539234 700614 539854 709082
rect 539234 700378 539266 700614
rect 539502 700378 539586 700614
rect 539822 700378 539854 700614
rect 539234 680614 539854 700378
rect 539234 680378 539266 680614
rect 539502 680378 539586 680614
rect 539822 680378 539854 680614
rect 539234 660614 539854 680378
rect 539234 660378 539266 660614
rect 539502 660378 539586 660614
rect 539822 660378 539854 660614
rect 539234 640614 539854 660378
rect 539234 640378 539266 640614
rect 539502 640378 539586 640614
rect 539822 640378 539854 640614
rect 539234 620614 539854 640378
rect 539234 620378 539266 620614
rect 539502 620378 539586 620614
rect 539822 620378 539854 620614
rect 539234 600614 539854 620378
rect 539234 600378 539266 600614
rect 539502 600378 539586 600614
rect 539822 600378 539854 600614
rect 539234 580614 539854 600378
rect 539234 580378 539266 580614
rect 539502 580378 539586 580614
rect 539822 580378 539854 580614
rect 539234 560614 539854 580378
rect 539234 560378 539266 560614
rect 539502 560378 539586 560614
rect 539822 560378 539854 560614
rect 539234 540614 539854 560378
rect 539234 540378 539266 540614
rect 539502 540378 539586 540614
rect 539822 540378 539854 540614
rect 539234 539308 539854 540378
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 683294 542414 704282
rect 541794 683058 541826 683294
rect 542062 683058 542146 683294
rect 542382 683058 542414 683294
rect 541794 663294 542414 683058
rect 541794 663058 541826 663294
rect 542062 663058 542146 663294
rect 542382 663058 542414 663294
rect 541794 643294 542414 663058
rect 541794 643058 541826 643294
rect 542062 643058 542146 643294
rect 542382 643058 542414 643294
rect 541794 623294 542414 643058
rect 541794 623058 541826 623294
rect 542062 623058 542146 623294
rect 542382 623058 542414 623294
rect 541794 603294 542414 623058
rect 541794 603058 541826 603294
rect 542062 603058 542146 603294
rect 542382 603058 542414 603294
rect 541794 583294 542414 603058
rect 541794 583058 541826 583294
rect 542062 583058 542146 583294
rect 542382 583058 542414 583294
rect 541794 563294 542414 583058
rect 541794 563058 541826 563294
rect 542062 563058 542146 563294
rect 542382 563058 542414 563294
rect 541794 543294 542414 563058
rect 541794 543058 541826 543294
rect 542062 543058 542146 543294
rect 542382 543058 542414 543294
rect 541794 539308 542414 543058
rect 542954 684274 543574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 542954 684038 542986 684274
rect 543222 684038 543306 684274
rect 543542 684038 543574 684274
rect 542954 664274 543574 684038
rect 542954 664038 542986 664274
rect 543222 664038 543306 664274
rect 543542 664038 543574 664274
rect 542954 644274 543574 664038
rect 542954 644038 542986 644274
rect 543222 644038 543306 644274
rect 543542 644038 543574 644274
rect 542954 624274 543574 644038
rect 542954 624038 542986 624274
rect 543222 624038 543306 624274
rect 543542 624038 543574 624274
rect 542954 604274 543574 624038
rect 542954 604038 542986 604274
rect 543222 604038 543306 604274
rect 543542 604038 543574 604274
rect 542954 584274 543574 604038
rect 542954 584038 542986 584274
rect 543222 584038 543306 584274
rect 543542 584038 543574 584274
rect 542954 564274 543574 584038
rect 542954 564038 542986 564274
rect 543222 564038 543306 564274
rect 543542 564038 543574 564274
rect 542954 544274 543574 564038
rect 542954 544038 542986 544274
rect 543222 544038 543306 544274
rect 543542 544038 543574 544274
rect 542954 539308 543574 544038
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 545514 686954 546134 706202
rect 545514 686718 545546 686954
rect 545782 686718 545866 686954
rect 546102 686718 546134 686954
rect 545514 666954 546134 686718
rect 545514 666718 545546 666954
rect 545782 666718 545866 666954
rect 546102 666718 546134 666954
rect 545514 646954 546134 666718
rect 545514 646718 545546 646954
rect 545782 646718 545866 646954
rect 546102 646718 546134 646954
rect 545514 626954 546134 646718
rect 545514 626718 545546 626954
rect 545782 626718 545866 626954
rect 546102 626718 546134 626954
rect 545514 606954 546134 626718
rect 545514 606718 545546 606954
rect 545782 606718 545866 606954
rect 546102 606718 546134 606954
rect 545514 586954 546134 606718
rect 545514 586718 545546 586954
rect 545782 586718 545866 586954
rect 546102 586718 546134 586954
rect 545514 566954 546134 586718
rect 545514 566718 545546 566954
rect 545782 566718 545866 566954
rect 546102 566718 546134 566954
rect 545514 546954 546134 566718
rect 545514 546718 545546 546954
rect 545782 546718 545866 546954
rect 546102 546718 546134 546954
rect 545514 539308 546134 546718
rect 549234 690614 549854 708122
rect 549234 690378 549266 690614
rect 549502 690378 549586 690614
rect 549822 690378 549854 690614
rect 549234 670614 549854 690378
rect 549234 670378 549266 670614
rect 549502 670378 549586 670614
rect 549822 670378 549854 670614
rect 549234 650614 549854 670378
rect 549234 650378 549266 650614
rect 549502 650378 549586 650614
rect 549822 650378 549854 650614
rect 549234 630614 549854 650378
rect 549234 630378 549266 630614
rect 549502 630378 549586 630614
rect 549822 630378 549854 630614
rect 549234 610614 549854 630378
rect 549234 610378 549266 610614
rect 549502 610378 549586 610614
rect 549822 610378 549854 610614
rect 549234 590614 549854 610378
rect 549234 590378 549266 590614
rect 549502 590378 549586 590614
rect 549822 590378 549854 590614
rect 549234 570614 549854 590378
rect 549234 570378 549266 570614
rect 549502 570378 549586 570614
rect 549822 570378 549854 570614
rect 549234 550614 549854 570378
rect 549234 550378 549266 550614
rect 549502 550378 549586 550614
rect 549822 550378 549854 550614
rect 540835 538796 540901 538797
rect 540835 538732 540836 538796
rect 540900 538732 540901 538796
rect 540835 538731 540901 538732
rect 529062 538170 529674 538230
rect 529614 537570 529674 538170
rect 540838 537570 540898 538731
rect 528326 537510 528524 537570
rect 529614 537510 529748 537570
rect 540838 537510 540900 537570
rect 528464 537202 528524 537510
rect 529688 537202 529748 537510
rect 540840 537202 540900 537510
rect 410272 533294 410620 533456
rect 410272 533058 410328 533294
rect 410564 533058 410620 533294
rect 410272 532896 410620 533058
rect 546000 533294 546348 533456
rect 546000 533058 546056 533294
rect 546292 533058 546348 533294
rect 546000 532896 546348 533058
rect 405514 526718 405546 526954
rect 405782 526718 405866 526954
rect 406102 526718 406134 526954
rect 405514 506954 406134 526718
rect 549234 530614 549854 550378
rect 549234 530378 549266 530614
rect 549502 530378 549586 530614
rect 549822 530378 549854 530614
rect 410952 523294 411300 523456
rect 410952 523058 411008 523294
rect 411244 523058 411300 523294
rect 410952 522896 411300 523058
rect 545320 523294 545668 523456
rect 545320 523058 545376 523294
rect 545612 523058 545668 523294
rect 545320 522896 545668 523058
rect 410272 513294 410620 513456
rect 410272 513058 410328 513294
rect 410564 513058 410620 513294
rect 410272 512896 410620 513058
rect 546000 513294 546348 513456
rect 546000 513058 546056 513294
rect 546292 513058 546348 513294
rect 546000 512896 546348 513058
rect 405514 506718 405546 506954
rect 405782 506718 405866 506954
rect 406102 506718 406134 506954
rect 405514 486954 406134 506718
rect 549234 510614 549854 530378
rect 549234 510378 549266 510614
rect 549502 510378 549586 510614
rect 549822 510378 549854 510614
rect 410952 503294 411300 503456
rect 410952 503058 411008 503294
rect 411244 503058 411300 503294
rect 410952 502896 411300 503058
rect 545320 503294 545668 503456
rect 545320 503058 545376 503294
rect 545612 503058 545668 503294
rect 545320 502896 545668 503058
rect 410272 493294 410620 493456
rect 410272 493058 410328 493294
rect 410564 493058 410620 493294
rect 410272 492896 410620 493058
rect 546000 493294 546348 493456
rect 546000 493058 546056 493294
rect 546292 493058 546348 493294
rect 546000 492896 546348 493058
rect 405514 486718 405546 486954
rect 405782 486718 405866 486954
rect 406102 486718 406134 486954
rect 405514 466954 406134 486718
rect 549234 490614 549854 510378
rect 549234 490378 549266 490614
rect 549502 490378 549586 490614
rect 549822 490378 549854 490614
rect 410952 483294 411300 483456
rect 410952 483058 411008 483294
rect 411244 483058 411300 483294
rect 410952 482896 411300 483058
rect 545320 483294 545668 483456
rect 545320 483058 545376 483294
rect 545612 483058 545668 483294
rect 545320 482896 545668 483058
rect 410272 473294 410620 473456
rect 410272 473058 410328 473294
rect 410564 473058 410620 473294
rect 410272 472896 410620 473058
rect 546000 473294 546348 473456
rect 546000 473058 546056 473294
rect 546292 473058 546348 473294
rect 546000 472896 546348 473058
rect 405514 466718 405546 466954
rect 405782 466718 405866 466954
rect 406102 466718 406134 466954
rect 405514 446954 406134 466718
rect 549234 470614 549854 490378
rect 549234 470378 549266 470614
rect 549502 470378 549586 470614
rect 549822 470378 549854 470614
rect 410952 463294 411300 463456
rect 410952 463058 411008 463294
rect 411244 463058 411300 463294
rect 410952 462896 411300 463058
rect 545320 463294 545668 463456
rect 545320 463058 545376 463294
rect 545612 463058 545668 463294
rect 545320 462896 545668 463058
rect 426056 453250 426116 454106
rect 427144 453250 427204 454106
rect 428232 453250 428292 454106
rect 429592 453797 429652 454106
rect 430544 453797 430604 454106
rect 431768 453797 431828 454106
rect 429589 453796 429655 453797
rect 429589 453732 429590 453796
rect 429654 453732 429655 453796
rect 429589 453731 429655 453732
rect 430541 453796 430607 453797
rect 430541 453732 430542 453796
rect 430606 453732 430607 453796
rect 430541 453731 430607 453732
rect 431765 453796 431831 453797
rect 431765 453732 431766 453796
rect 431830 453732 431831 453796
rect 433128 453794 433188 454106
rect 434216 453794 434276 454106
rect 435440 453794 435500 454106
rect 436528 453794 436588 454106
rect 431765 453731 431831 453732
rect 433014 453734 433188 453794
rect 434118 453734 434276 453794
rect 435406 453734 435500 453794
rect 436510 453734 436588 453794
rect 429592 453250 429652 453731
rect 426022 453190 426116 453250
rect 427126 453190 427204 453250
rect 428230 453190 428292 453250
rect 429518 453190 429652 453250
rect 426022 452573 426082 453190
rect 427126 452573 427186 453190
rect 428230 452573 428290 453190
rect 429518 452573 429578 453190
rect 433014 452573 433074 453734
rect 434118 452573 434178 453734
rect 435406 452573 435466 453734
rect 436510 452573 436570 453734
rect 437616 453250 437676 454106
rect 437614 453190 437676 453250
rect 438296 453250 438356 454106
rect 438704 453250 438764 454106
rect 440064 453250 440124 454106
rect 440744 453250 440804 454106
rect 438296 453190 438410 453250
rect 438704 453190 438778 453250
rect 426019 452572 426085 452573
rect 426019 452508 426020 452572
rect 426084 452508 426085 452572
rect 426019 452507 426085 452508
rect 427123 452572 427189 452573
rect 427123 452508 427124 452572
rect 427188 452508 427189 452572
rect 427123 452507 427189 452508
rect 428227 452572 428293 452573
rect 428227 452508 428228 452572
rect 428292 452508 428293 452572
rect 428227 452507 428293 452508
rect 429515 452572 429581 452573
rect 429515 452508 429516 452572
rect 429580 452508 429581 452572
rect 429515 452507 429581 452508
rect 433011 452572 433077 452573
rect 433011 452508 433012 452572
rect 433076 452508 433077 452572
rect 433011 452507 433077 452508
rect 434115 452572 434181 452573
rect 434115 452508 434116 452572
rect 434180 452508 434181 452572
rect 434115 452507 434181 452508
rect 435403 452572 435469 452573
rect 435403 452508 435404 452572
rect 435468 452508 435469 452572
rect 435403 452507 435469 452508
rect 436507 452572 436573 452573
rect 436507 452508 436508 452572
rect 436572 452508 436573 452572
rect 436507 452507 436573 452508
rect 405514 446718 405546 446954
rect 405782 446718 405866 446954
rect 406102 446718 406134 446954
rect 405514 426954 406134 446718
rect 405514 426718 405546 426954
rect 405782 426718 405866 426954
rect 406102 426718 406134 426954
rect 405514 421162 406134 426718
rect 409234 450614 409854 452000
rect 409234 450378 409266 450614
rect 409502 450378 409586 450614
rect 409822 450378 409854 450614
rect 409234 430614 409854 450378
rect 409234 430378 409266 430614
rect 409502 430378 409586 430614
rect 409822 430378 409854 430614
rect 409234 421162 409854 430378
rect 411794 433294 412414 452000
rect 411794 433058 411826 433294
rect 412062 433058 412146 433294
rect 412382 433058 412414 433294
rect 411794 421162 412414 433058
rect 412954 434274 413574 452000
rect 412954 434038 412986 434274
rect 413222 434038 413306 434274
rect 413542 434038 413574 434274
rect 412954 421162 413574 434038
rect 415514 436954 416134 452000
rect 415514 436718 415546 436954
rect 415782 436718 415866 436954
rect 416102 436718 416134 436954
rect 415514 421162 416134 436718
rect 419234 440614 419854 452000
rect 419234 440378 419266 440614
rect 419502 440378 419586 440614
rect 419822 440378 419854 440614
rect 419234 421162 419854 440378
rect 421794 443294 422414 452000
rect 421794 443058 421826 443294
rect 422062 443058 422146 443294
rect 422382 443058 422414 443294
rect 421794 423294 422414 443058
rect 421794 423058 421826 423294
rect 422062 423058 422146 423294
rect 422382 423058 422414 423294
rect 421794 421162 422414 423058
rect 422954 444274 423574 452000
rect 422954 444038 422986 444274
rect 423222 444038 423306 444274
rect 423542 444038 423574 444274
rect 422954 424274 423574 444038
rect 422954 424038 422986 424274
rect 423222 424038 423306 424274
rect 423542 424038 423574 424274
rect 422954 421162 423574 424038
rect 425514 446954 426134 452000
rect 425514 446718 425546 446954
rect 425782 446718 425866 446954
rect 426102 446718 426134 446954
rect 425514 426954 426134 446718
rect 425514 426718 425546 426954
rect 425782 426718 425866 426954
rect 426102 426718 426134 426954
rect 425514 421162 426134 426718
rect 429234 450614 429854 452000
rect 429234 450378 429266 450614
rect 429502 450378 429586 450614
rect 429822 450378 429854 450614
rect 429234 430614 429854 450378
rect 429234 430378 429266 430614
rect 429502 430378 429586 430614
rect 429822 430378 429854 430614
rect 429234 421162 429854 430378
rect 431794 433294 432414 452000
rect 431794 433058 431826 433294
rect 432062 433058 432146 433294
rect 432382 433058 432414 433294
rect 431794 421162 432414 433058
rect 432954 434274 433574 452000
rect 432954 434038 432986 434274
rect 433222 434038 433306 434274
rect 433542 434038 433574 434274
rect 432954 421162 433574 434038
rect 435514 436954 436134 452000
rect 437614 451349 437674 453190
rect 438350 452301 438410 453190
rect 438347 452300 438413 452301
rect 438347 452236 438348 452300
rect 438412 452236 438413 452300
rect 438347 452235 438413 452236
rect 438718 451621 438778 453190
rect 440006 453190 440124 453250
rect 440742 453190 440804 453250
rect 441288 453250 441348 454106
rect 442376 453250 442436 454106
rect 443464 453250 443524 454106
rect 443600 453661 443660 454106
rect 443597 453660 443663 453661
rect 443597 453596 443598 453660
rect 443662 453596 443663 453660
rect 443597 453595 443663 453596
rect 444552 453250 444612 454106
rect 445912 453250 445972 454106
rect 441288 453190 441354 453250
rect 442376 453190 442458 453250
rect 443464 453190 443562 453250
rect 444552 453190 444666 453250
rect 438715 451620 438781 451621
rect 438715 451556 438716 451620
rect 438780 451556 438781 451620
rect 438715 451555 438781 451556
rect 437611 451348 437677 451349
rect 437611 451284 437612 451348
rect 437676 451284 437677 451348
rect 437611 451283 437677 451284
rect 435514 436718 435546 436954
rect 435782 436718 435866 436954
rect 436102 436718 436134 436954
rect 435514 421162 436134 436718
rect 439234 440614 439854 452000
rect 440006 451349 440066 453190
rect 440742 451349 440802 453190
rect 441294 451621 441354 453190
rect 442398 452165 442458 453190
rect 443502 452165 443562 453190
rect 442395 452164 442461 452165
rect 442395 452100 442396 452164
rect 442460 452100 442461 452164
rect 442395 452099 442461 452100
rect 443499 452164 443565 452165
rect 443499 452100 443500 452164
rect 443564 452100 443565 452164
rect 443499 452099 443565 452100
rect 441291 451620 441357 451621
rect 441291 451556 441292 451620
rect 441356 451556 441357 451620
rect 441291 451555 441357 451556
rect 440003 451348 440069 451349
rect 440003 451284 440004 451348
rect 440068 451284 440069 451348
rect 440003 451283 440069 451284
rect 440739 451348 440805 451349
rect 440739 451284 440740 451348
rect 440804 451284 440805 451348
rect 440739 451283 440805 451284
rect 439234 440378 439266 440614
rect 439502 440378 439586 440614
rect 439822 440378 439854 440614
rect 439234 421162 439854 440378
rect 441794 443294 442414 452000
rect 441794 443058 441826 443294
rect 442062 443058 442146 443294
rect 442382 443058 442414 443294
rect 441794 423294 442414 443058
rect 441794 423058 441826 423294
rect 442062 423058 442146 423294
rect 442382 423058 442414 423294
rect 441794 421162 442414 423058
rect 442954 444274 443574 452000
rect 444606 451349 444666 453190
rect 445894 453190 445972 453250
rect 446048 453250 446108 454106
rect 447000 453250 447060 454106
rect 446048 453190 446138 453250
rect 445894 452165 445954 453190
rect 446078 452165 446138 453190
rect 446998 453190 447060 453250
rect 448088 453250 448148 454106
rect 448496 453250 448556 454106
rect 449448 453250 449508 454106
rect 448088 453190 448162 453250
rect 445891 452164 445957 452165
rect 445891 452100 445892 452164
rect 445956 452100 445957 452164
rect 445891 452099 445957 452100
rect 446075 452164 446141 452165
rect 446075 452100 446076 452164
rect 446140 452100 446141 452164
rect 446075 452099 446141 452100
rect 444603 451348 444669 451349
rect 444603 451284 444604 451348
rect 444668 451284 444669 451348
rect 444603 451283 444669 451284
rect 442954 444038 442986 444274
rect 443222 444038 443306 444274
rect 443542 444038 443574 444274
rect 442954 424274 443574 444038
rect 442954 424038 442986 424274
rect 443222 424038 443306 424274
rect 443542 424038 443574 424274
rect 442954 421162 443574 424038
rect 445514 446954 446134 452000
rect 446998 451349 447058 453190
rect 448102 451349 448162 453190
rect 448470 453190 448556 453250
rect 449390 453190 449508 453250
rect 450672 453250 450732 454106
rect 451080 453250 451140 454106
rect 450672 453190 450738 453250
rect 448470 451349 448530 453190
rect 449390 452165 449450 453190
rect 450678 452573 450738 453190
rect 451046 453190 451140 453250
rect 451760 453250 451820 454106
rect 452848 453250 452908 454106
rect 453528 453250 453588 454106
rect 453936 453250 453996 454106
rect 455296 453250 455356 454106
rect 451760 453190 451842 453250
rect 452848 453190 452946 453250
rect 453528 453190 453682 453250
rect 453936 453190 454050 453250
rect 450675 452572 450741 452573
rect 450675 452508 450676 452572
rect 450740 452508 450741 452572
rect 450675 452507 450741 452508
rect 449387 452164 449453 452165
rect 449387 452100 449388 452164
rect 449452 452100 449453 452164
rect 449387 452099 449453 452100
rect 446995 451348 447061 451349
rect 446995 451284 446996 451348
rect 447060 451284 447061 451348
rect 446995 451283 447061 451284
rect 448099 451348 448165 451349
rect 448099 451284 448100 451348
rect 448164 451284 448165 451348
rect 448099 451283 448165 451284
rect 448467 451348 448533 451349
rect 448467 451284 448468 451348
rect 448532 451284 448533 451348
rect 448467 451283 448533 451284
rect 445514 446718 445546 446954
rect 445782 446718 445866 446954
rect 446102 446718 446134 446954
rect 445514 426954 446134 446718
rect 445514 426718 445546 426954
rect 445782 426718 445866 426954
rect 446102 426718 446134 426954
rect 445514 421162 446134 426718
rect 449234 450614 449854 452000
rect 451046 451349 451106 453190
rect 451782 452165 451842 453190
rect 452886 452573 452946 453190
rect 452883 452572 452949 452573
rect 452883 452508 452884 452572
rect 452948 452508 452949 452572
rect 452883 452507 452949 452508
rect 453622 452165 453682 453190
rect 451779 452164 451845 452165
rect 451779 452100 451780 452164
rect 451844 452100 451845 452164
rect 451779 452099 451845 452100
rect 453619 452164 453685 452165
rect 453619 452100 453620 452164
rect 453684 452100 453685 452164
rect 453619 452099 453685 452100
rect 451043 451348 451109 451349
rect 451043 451284 451044 451348
rect 451108 451284 451109 451348
rect 451043 451283 451109 451284
rect 449234 450378 449266 450614
rect 449502 450378 449586 450614
rect 449822 450378 449854 450614
rect 449234 430614 449854 450378
rect 449234 430378 449266 430614
rect 449502 430378 449586 430614
rect 449822 430378 449854 430614
rect 449234 421162 449854 430378
rect 451794 433294 452414 452000
rect 451794 433058 451826 433294
rect 452062 433058 452146 433294
rect 452382 433058 452414 433294
rect 451794 421162 452414 433058
rect 452954 434274 453574 452000
rect 453990 451349 454050 453190
rect 455278 453190 455356 453250
rect 455976 453250 456036 454106
rect 456384 453250 456444 454106
rect 455976 453190 456074 453250
rect 455278 452301 455338 453190
rect 455275 452300 455341 452301
rect 455275 452236 455276 452300
rect 455340 452236 455341 452300
rect 455275 452235 455341 452236
rect 456014 452165 456074 453190
rect 456382 453190 456444 453250
rect 457608 453250 457668 454106
rect 458288 453250 458348 454106
rect 458696 453250 458756 454106
rect 459784 453250 459844 454106
rect 461008 453250 461068 454106
rect 457608 453190 457730 453250
rect 458288 453190 458466 453250
rect 456011 452164 456077 452165
rect 456011 452100 456012 452164
rect 456076 452100 456077 452164
rect 456011 452099 456077 452100
rect 453987 451348 454053 451349
rect 453987 451284 453988 451348
rect 454052 451284 454053 451348
rect 453987 451283 454053 451284
rect 452954 434038 452986 434274
rect 453222 434038 453306 434274
rect 453542 434038 453574 434274
rect 452954 421162 453574 434038
rect 455514 436954 456134 452000
rect 456382 451349 456442 453190
rect 457670 451349 457730 453190
rect 458406 451621 458466 453190
rect 458590 453190 458756 453250
rect 459694 453190 459844 453250
rect 460982 453190 461068 453250
rect 461144 453250 461204 454106
rect 462232 453250 462292 454106
rect 463320 453250 463380 454106
rect 463592 453250 463652 454106
rect 464408 453250 464468 454106
rect 465768 454040 465828 454106
rect 461144 453190 461226 453250
rect 462232 453190 462330 453250
rect 463320 453190 463434 453250
rect 458403 451620 458469 451621
rect 458403 451556 458404 451620
rect 458468 451556 458469 451620
rect 458403 451555 458469 451556
rect 458590 451349 458650 453190
rect 459694 452165 459754 453190
rect 459691 452164 459757 452165
rect 459691 452100 459692 452164
rect 459756 452100 459757 452164
rect 459691 452099 459757 452100
rect 456379 451348 456445 451349
rect 456379 451284 456380 451348
rect 456444 451284 456445 451348
rect 456379 451283 456445 451284
rect 457667 451348 457733 451349
rect 457667 451284 457668 451348
rect 457732 451284 457733 451348
rect 457667 451283 457733 451284
rect 458587 451348 458653 451349
rect 458587 451284 458588 451348
rect 458652 451284 458653 451348
rect 458587 451283 458653 451284
rect 455514 436718 455546 436954
rect 455782 436718 455866 436954
rect 456102 436718 456134 436954
rect 455514 421162 456134 436718
rect 459234 440614 459854 452000
rect 460982 449173 461042 453190
rect 461166 449309 461226 453190
rect 462270 452165 462330 453190
rect 463374 452301 463434 453190
rect 463558 453190 463652 453250
rect 464294 453190 464468 453250
rect 465766 453980 465828 454040
rect 463371 452300 463437 452301
rect 463371 452236 463372 452300
rect 463436 452236 463437 452300
rect 463371 452235 463437 452236
rect 463558 452165 463618 453190
rect 462267 452164 462333 452165
rect 462267 452100 462268 452164
rect 462332 452100 462333 452164
rect 462267 452099 462333 452100
rect 463555 452164 463621 452165
rect 463555 452100 463556 452164
rect 463620 452100 463621 452164
rect 463555 452099 463621 452100
rect 461163 449308 461229 449309
rect 461163 449244 461164 449308
rect 461228 449244 461229 449308
rect 461163 449243 461229 449244
rect 460979 449172 461045 449173
rect 460979 449108 460980 449172
rect 461044 449108 461045 449172
rect 460979 449107 461045 449108
rect 459234 440378 459266 440614
rect 459502 440378 459586 440614
rect 459822 440378 459854 440614
rect 459234 421162 459854 440378
rect 461794 443294 462414 452000
rect 461794 443058 461826 443294
rect 462062 443058 462146 443294
rect 462382 443058 462414 443294
rect 461794 423294 462414 443058
rect 461794 423058 461826 423294
rect 462062 423058 462146 423294
rect 462382 423058 462414 423294
rect 461794 421162 462414 423058
rect 462954 444274 463574 452000
rect 464294 451349 464354 453190
rect 465766 452165 465826 453980
rect 466040 453250 466100 454106
rect 466992 453250 467052 454106
rect 468080 453250 468140 454106
rect 466040 453190 466194 453250
rect 466992 453190 467114 453250
rect 466134 452573 466194 453190
rect 467054 452573 467114 453190
rect 467974 453190 468140 453250
rect 468488 453250 468548 454106
rect 469168 453250 469228 454106
rect 470936 453250 470996 454106
rect 473520 453250 473580 454106
rect 468488 453190 468586 453250
rect 467974 452573 468034 453190
rect 468526 452573 468586 453190
rect 469078 453190 469228 453250
rect 470918 453190 470996 453250
rect 473494 453190 473580 453250
rect 475968 453250 476028 454106
rect 478280 453250 478340 454106
rect 475968 453190 476130 453250
rect 466131 452572 466197 452573
rect 466131 452508 466132 452572
rect 466196 452508 466197 452572
rect 466131 452507 466197 452508
rect 467051 452572 467117 452573
rect 467051 452508 467052 452572
rect 467116 452508 467117 452572
rect 467051 452507 467117 452508
rect 467971 452572 468037 452573
rect 467971 452508 467972 452572
rect 468036 452508 468037 452572
rect 467971 452507 468037 452508
rect 468523 452572 468589 452573
rect 468523 452508 468524 452572
rect 468588 452508 468589 452572
rect 468523 452507 468589 452508
rect 469078 452301 469138 453190
rect 470918 452573 470978 453190
rect 473494 452573 473554 453190
rect 476070 452573 476130 453190
rect 478278 453190 478340 453250
rect 481000 453250 481060 454106
rect 483448 453250 483508 454106
rect 481000 453190 481098 453250
rect 478278 452573 478338 453190
rect 481038 452573 481098 453190
rect 483430 453190 483508 453250
rect 485896 453250 485956 454106
rect 488480 453250 488540 454106
rect 485896 453190 486066 453250
rect 483430 452573 483490 453190
rect 486006 452573 486066 453190
rect 488398 453190 488540 453250
rect 490928 453250 490988 454106
rect 493512 453250 493572 454106
rect 495960 453250 496020 454106
rect 498544 453250 498604 454106
rect 490928 453190 491034 453250
rect 493512 453190 493610 453250
rect 488398 452573 488458 453190
rect 490974 452573 491034 453190
rect 493550 452573 493610 453190
rect 495942 453190 496020 453250
rect 498518 453190 498604 453250
rect 500992 453250 501052 454106
rect 503440 453250 503500 454106
rect 505888 453250 505948 454106
rect 508472 453250 508532 454106
rect 500992 453190 501154 453250
rect 503440 453190 503546 453250
rect 495942 452573 496002 453190
rect 498518 452573 498578 453190
rect 501094 452573 501154 453190
rect 503486 452573 503546 453190
rect 505878 453190 505948 453250
rect 508454 453190 508532 453250
rect 510920 453250 510980 454106
rect 513368 453250 513428 454106
rect 515952 453250 516012 454106
rect 533224 453661 533284 454106
rect 532739 453660 532805 453661
rect 532739 453596 532740 453660
rect 532804 453596 532805 453660
rect 532739 453595 532805 453596
rect 533221 453660 533287 453661
rect 533221 453596 533222 453660
rect 533286 453596 533287 453660
rect 533221 453595 533287 453596
rect 510920 453190 511090 453250
rect 513368 453190 513482 453250
rect 515952 453190 516058 453250
rect 505878 452573 505938 453190
rect 508454 452573 508514 453190
rect 511030 452573 511090 453190
rect 513422 452573 513482 453190
rect 515998 452573 516058 453190
rect 470915 452572 470981 452573
rect 470915 452508 470916 452572
rect 470980 452508 470981 452572
rect 470915 452507 470981 452508
rect 473491 452572 473557 452573
rect 473491 452508 473492 452572
rect 473556 452508 473557 452572
rect 473491 452507 473557 452508
rect 476067 452572 476133 452573
rect 476067 452508 476068 452572
rect 476132 452508 476133 452572
rect 476067 452507 476133 452508
rect 478275 452572 478341 452573
rect 478275 452508 478276 452572
rect 478340 452508 478341 452572
rect 478275 452507 478341 452508
rect 481035 452572 481101 452573
rect 481035 452508 481036 452572
rect 481100 452508 481101 452572
rect 481035 452507 481101 452508
rect 483427 452572 483493 452573
rect 483427 452508 483428 452572
rect 483492 452508 483493 452572
rect 483427 452507 483493 452508
rect 486003 452572 486069 452573
rect 486003 452508 486004 452572
rect 486068 452508 486069 452572
rect 486003 452507 486069 452508
rect 488395 452572 488461 452573
rect 488395 452508 488396 452572
rect 488460 452508 488461 452572
rect 488395 452507 488461 452508
rect 490971 452572 491037 452573
rect 490971 452508 490972 452572
rect 491036 452508 491037 452572
rect 490971 452507 491037 452508
rect 493547 452572 493613 452573
rect 493547 452508 493548 452572
rect 493612 452508 493613 452572
rect 493547 452507 493613 452508
rect 495939 452572 496005 452573
rect 495939 452508 495940 452572
rect 496004 452508 496005 452572
rect 495939 452507 496005 452508
rect 498515 452572 498581 452573
rect 498515 452508 498516 452572
rect 498580 452508 498581 452572
rect 498515 452507 498581 452508
rect 501091 452572 501157 452573
rect 501091 452508 501092 452572
rect 501156 452508 501157 452572
rect 501091 452507 501157 452508
rect 503483 452572 503549 452573
rect 503483 452508 503484 452572
rect 503548 452508 503549 452572
rect 503483 452507 503549 452508
rect 505875 452572 505941 452573
rect 505875 452508 505876 452572
rect 505940 452508 505941 452572
rect 505875 452507 505941 452508
rect 508451 452572 508517 452573
rect 508451 452508 508452 452572
rect 508516 452508 508517 452572
rect 508451 452507 508517 452508
rect 511027 452572 511093 452573
rect 511027 452508 511028 452572
rect 511092 452508 511093 452572
rect 511027 452507 511093 452508
rect 513419 452572 513485 452573
rect 513419 452508 513420 452572
rect 513484 452508 513485 452572
rect 513419 452507 513485 452508
rect 515995 452572 516061 452573
rect 515995 452508 515996 452572
rect 516060 452508 516061 452572
rect 515995 452507 516061 452508
rect 469075 452300 469141 452301
rect 469075 452236 469076 452300
rect 469140 452236 469141 452300
rect 469075 452235 469141 452236
rect 465763 452164 465829 452165
rect 465763 452100 465764 452164
rect 465828 452100 465829 452164
rect 465763 452099 465829 452100
rect 464291 451348 464357 451349
rect 464291 451284 464292 451348
rect 464356 451284 464357 451348
rect 464291 451283 464357 451284
rect 462954 444038 462986 444274
rect 463222 444038 463306 444274
rect 463542 444038 463574 444274
rect 462954 424274 463574 444038
rect 462954 424038 462986 424274
rect 463222 424038 463306 424274
rect 463542 424038 463574 424274
rect 462954 421162 463574 424038
rect 465514 446954 466134 452000
rect 465514 446718 465546 446954
rect 465782 446718 465866 446954
rect 466102 446718 466134 446954
rect 465514 426954 466134 446718
rect 465514 426718 465546 426954
rect 465782 426718 465866 426954
rect 466102 426718 466134 426954
rect 465514 421162 466134 426718
rect 469234 450614 469854 452000
rect 469234 450378 469266 450614
rect 469502 450378 469586 450614
rect 469822 450378 469854 450614
rect 469234 430614 469854 450378
rect 469234 430378 469266 430614
rect 469502 430378 469586 430614
rect 469822 430378 469854 430614
rect 469234 421162 469854 430378
rect 471794 433294 472414 452000
rect 471794 433058 471826 433294
rect 472062 433058 472146 433294
rect 472382 433058 472414 433294
rect 471794 421162 472414 433058
rect 472954 434274 473574 452000
rect 472954 434038 472986 434274
rect 473222 434038 473306 434274
rect 473542 434038 473574 434274
rect 472954 421162 473574 434038
rect 475514 436954 476134 452000
rect 475514 436718 475546 436954
rect 475782 436718 475866 436954
rect 476102 436718 476134 436954
rect 475514 421162 476134 436718
rect 479234 440614 479854 452000
rect 479234 440378 479266 440614
rect 479502 440378 479586 440614
rect 479822 440378 479854 440614
rect 479234 421162 479854 440378
rect 481794 443294 482414 452000
rect 481794 443058 481826 443294
rect 482062 443058 482146 443294
rect 482382 443058 482414 443294
rect 481794 423294 482414 443058
rect 481794 423058 481826 423294
rect 482062 423058 482146 423294
rect 482382 423058 482414 423294
rect 481794 421162 482414 423058
rect 482954 444274 483574 452000
rect 482954 444038 482986 444274
rect 483222 444038 483306 444274
rect 483542 444038 483574 444274
rect 482954 424274 483574 444038
rect 482954 424038 482986 424274
rect 483222 424038 483306 424274
rect 483542 424038 483574 424274
rect 482954 421162 483574 424038
rect 485514 446954 486134 452000
rect 485514 446718 485546 446954
rect 485782 446718 485866 446954
rect 486102 446718 486134 446954
rect 485514 426954 486134 446718
rect 485514 426718 485546 426954
rect 485782 426718 485866 426954
rect 486102 426718 486134 426954
rect 485514 421162 486134 426718
rect 489234 450614 489854 452000
rect 489234 450378 489266 450614
rect 489502 450378 489586 450614
rect 489822 450378 489854 450614
rect 489234 430614 489854 450378
rect 489234 430378 489266 430614
rect 489502 430378 489586 430614
rect 489822 430378 489854 430614
rect 489234 421162 489854 430378
rect 491794 433294 492414 452000
rect 491794 433058 491826 433294
rect 492062 433058 492146 433294
rect 492382 433058 492414 433294
rect 491794 421162 492414 433058
rect 492954 434274 493574 452000
rect 492954 434038 492986 434274
rect 493222 434038 493306 434274
rect 493542 434038 493574 434274
rect 492954 421162 493574 434038
rect 495514 436954 496134 452000
rect 495514 436718 495546 436954
rect 495782 436718 495866 436954
rect 496102 436718 496134 436954
rect 495514 421162 496134 436718
rect 499234 440614 499854 452000
rect 499234 440378 499266 440614
rect 499502 440378 499586 440614
rect 499822 440378 499854 440614
rect 499234 421162 499854 440378
rect 501794 443294 502414 452000
rect 501794 443058 501826 443294
rect 502062 443058 502146 443294
rect 502382 443058 502414 443294
rect 501794 423294 502414 443058
rect 501794 423058 501826 423294
rect 502062 423058 502146 423294
rect 502382 423058 502414 423294
rect 501794 421162 502414 423058
rect 502954 444274 503574 452000
rect 502954 444038 502986 444274
rect 503222 444038 503306 444274
rect 503542 444038 503574 444274
rect 502954 424274 503574 444038
rect 502954 424038 502986 424274
rect 503222 424038 503306 424274
rect 503542 424038 503574 424274
rect 502954 421162 503574 424038
rect 505514 446954 506134 452000
rect 505514 446718 505546 446954
rect 505782 446718 505866 446954
rect 506102 446718 506134 446954
rect 505514 426954 506134 446718
rect 505514 426718 505546 426954
rect 505782 426718 505866 426954
rect 506102 426718 506134 426954
rect 505514 421162 506134 426718
rect 509234 450614 509854 452000
rect 509234 450378 509266 450614
rect 509502 450378 509586 450614
rect 509822 450378 509854 450614
rect 509234 430614 509854 450378
rect 509234 430378 509266 430614
rect 509502 430378 509586 430614
rect 509822 430378 509854 430614
rect 509234 421162 509854 430378
rect 511794 433294 512414 452000
rect 511794 433058 511826 433294
rect 512062 433058 512146 433294
rect 512382 433058 512414 433294
rect 511794 421162 512414 433058
rect 512954 434274 513574 452000
rect 512954 434038 512986 434274
rect 513222 434038 513306 434274
rect 513542 434038 513574 434274
rect 512954 421162 513574 434038
rect 515514 436954 516134 452000
rect 515514 436718 515546 436954
rect 515782 436718 515866 436954
rect 516102 436718 516134 436954
rect 515514 421162 516134 436718
rect 519234 440614 519854 452000
rect 519234 440378 519266 440614
rect 519502 440378 519586 440614
rect 519822 440378 519854 440614
rect 519234 421162 519854 440378
rect 521794 443294 522414 452000
rect 521794 443058 521826 443294
rect 522062 443058 522146 443294
rect 522382 443058 522414 443294
rect 521794 423294 522414 443058
rect 521794 423058 521826 423294
rect 522062 423058 522146 423294
rect 522382 423058 522414 423294
rect 521794 421162 522414 423058
rect 522954 444274 523574 452000
rect 522954 444038 522986 444274
rect 523222 444038 523306 444274
rect 523542 444038 523574 444274
rect 522954 424274 523574 444038
rect 522954 424038 522986 424274
rect 523222 424038 523306 424274
rect 523542 424038 523574 424274
rect 522954 421162 523574 424038
rect 525514 446954 526134 452000
rect 525514 446718 525546 446954
rect 525782 446718 525866 446954
rect 526102 446718 526134 446954
rect 525514 426954 526134 446718
rect 525514 426718 525546 426954
rect 525782 426718 525866 426954
rect 526102 426718 526134 426954
rect 525514 421162 526134 426718
rect 529234 450614 529854 452000
rect 529234 450378 529266 450614
rect 529502 450378 529586 450614
rect 529822 450378 529854 450614
rect 529234 430614 529854 450378
rect 529234 430378 529266 430614
rect 529502 430378 529586 430614
rect 529822 430378 529854 430614
rect 529234 421162 529854 430378
rect 531794 433294 532414 452000
rect 532742 451485 532802 453595
rect 533360 453250 533420 454106
rect 533294 453190 533420 453250
rect 533294 452437 533354 453190
rect 533291 452436 533357 452437
rect 533291 452372 533292 452436
rect 533356 452372 533357 452436
rect 533291 452371 533357 452372
rect 532739 451484 532805 451485
rect 532739 451420 532740 451484
rect 532804 451420 532805 451484
rect 532739 451419 532805 451420
rect 531794 433058 531826 433294
rect 532062 433058 532146 433294
rect 532382 433058 532414 433294
rect 531794 421162 532414 433058
rect 532954 434274 533574 452000
rect 532954 434038 532986 434274
rect 533222 434038 533306 434274
rect 533542 434038 533574 434274
rect 532954 421162 533574 434038
rect 535514 436954 536134 452000
rect 535514 436718 535546 436954
rect 535782 436718 535866 436954
rect 536102 436718 536134 436954
rect 535514 421162 536134 436718
rect 539234 440614 539854 452000
rect 539234 440378 539266 440614
rect 539502 440378 539586 440614
rect 539822 440378 539854 440614
rect 539234 421162 539854 440378
rect 541794 443294 542414 452000
rect 541794 443058 541826 443294
rect 542062 443058 542146 443294
rect 542382 443058 542414 443294
rect 541794 423294 542414 443058
rect 541794 423058 541826 423294
rect 542062 423058 542146 423294
rect 542382 423058 542414 423294
rect 541794 421162 542414 423058
rect 542954 444274 543574 452000
rect 542954 444038 542986 444274
rect 543222 444038 543306 444274
rect 543542 444038 543574 444274
rect 542954 424274 543574 444038
rect 542954 424038 542986 424274
rect 543222 424038 543306 424274
rect 543542 424038 543574 424274
rect 542954 421162 543574 424038
rect 545514 446954 546134 452000
rect 545514 446718 545546 446954
rect 545782 446718 545866 446954
rect 546102 446718 546134 446954
rect 545514 426954 546134 446718
rect 545514 426718 545546 426954
rect 545782 426718 545866 426954
rect 546102 426718 546134 426954
rect 545514 421162 546134 426718
rect 549234 450614 549854 470378
rect 549234 450378 549266 450614
rect 549502 450378 549586 450614
rect 549822 450378 549854 450614
rect 549234 430614 549854 450378
rect 549234 430378 549266 430614
rect 549502 430378 549586 430614
rect 549822 430378 549854 430614
rect 549234 421162 549854 430378
rect 551794 705798 552414 705830
rect 551794 705562 551826 705798
rect 552062 705562 552146 705798
rect 552382 705562 552414 705798
rect 551794 705478 552414 705562
rect 551794 705242 551826 705478
rect 552062 705242 552146 705478
rect 552382 705242 552414 705478
rect 551794 693294 552414 705242
rect 551794 693058 551826 693294
rect 552062 693058 552146 693294
rect 552382 693058 552414 693294
rect 551794 673294 552414 693058
rect 551794 673058 551826 673294
rect 552062 673058 552146 673294
rect 552382 673058 552414 673294
rect 551794 653294 552414 673058
rect 551794 653058 551826 653294
rect 552062 653058 552146 653294
rect 552382 653058 552414 653294
rect 551794 633294 552414 653058
rect 551794 633058 551826 633294
rect 552062 633058 552146 633294
rect 552382 633058 552414 633294
rect 551794 613294 552414 633058
rect 551794 613058 551826 613294
rect 552062 613058 552146 613294
rect 552382 613058 552414 613294
rect 551794 593294 552414 613058
rect 551794 593058 551826 593294
rect 552062 593058 552146 593294
rect 552382 593058 552414 593294
rect 551794 573294 552414 593058
rect 551794 573058 551826 573294
rect 552062 573058 552146 573294
rect 552382 573058 552414 573294
rect 551794 553294 552414 573058
rect 551794 553058 551826 553294
rect 552062 553058 552146 553294
rect 552382 553058 552414 553294
rect 551794 533294 552414 553058
rect 551794 533058 551826 533294
rect 552062 533058 552146 533294
rect 552382 533058 552414 533294
rect 551794 513294 552414 533058
rect 551794 513058 551826 513294
rect 552062 513058 552146 513294
rect 552382 513058 552414 513294
rect 551794 493294 552414 513058
rect 551794 493058 551826 493294
rect 552062 493058 552146 493294
rect 552382 493058 552414 493294
rect 551794 473294 552414 493058
rect 551794 473058 551826 473294
rect 552062 473058 552146 473294
rect 552382 473058 552414 473294
rect 551794 453294 552414 473058
rect 551794 453058 551826 453294
rect 552062 453058 552146 453294
rect 552382 453058 552414 453294
rect 551794 433294 552414 453058
rect 551794 433058 551826 433294
rect 552062 433058 552146 433294
rect 552382 433058 552414 433294
rect 551794 421162 552414 433058
rect 552954 694274 553574 710042
rect 562954 711558 563574 711590
rect 562954 711322 562986 711558
rect 563222 711322 563306 711558
rect 563542 711322 563574 711558
rect 562954 711238 563574 711322
rect 562954 711002 562986 711238
rect 563222 711002 563306 711238
rect 563542 711002 563574 711238
rect 559234 709638 559854 709670
rect 559234 709402 559266 709638
rect 559502 709402 559586 709638
rect 559822 709402 559854 709638
rect 559234 709318 559854 709402
rect 559234 709082 559266 709318
rect 559502 709082 559586 709318
rect 559822 709082 559854 709318
rect 552954 694038 552986 694274
rect 553222 694038 553306 694274
rect 553542 694038 553574 694274
rect 552954 674274 553574 694038
rect 552954 674038 552986 674274
rect 553222 674038 553306 674274
rect 553542 674038 553574 674274
rect 552954 654274 553574 674038
rect 552954 654038 552986 654274
rect 553222 654038 553306 654274
rect 553542 654038 553574 654274
rect 552954 634274 553574 654038
rect 552954 634038 552986 634274
rect 553222 634038 553306 634274
rect 553542 634038 553574 634274
rect 552954 614274 553574 634038
rect 552954 614038 552986 614274
rect 553222 614038 553306 614274
rect 553542 614038 553574 614274
rect 552954 594274 553574 614038
rect 552954 594038 552986 594274
rect 553222 594038 553306 594274
rect 553542 594038 553574 594274
rect 552954 574274 553574 594038
rect 552954 574038 552986 574274
rect 553222 574038 553306 574274
rect 553542 574038 553574 574274
rect 552954 554274 553574 574038
rect 552954 554038 552986 554274
rect 553222 554038 553306 554274
rect 553542 554038 553574 554274
rect 552954 534274 553574 554038
rect 552954 534038 552986 534274
rect 553222 534038 553306 534274
rect 553542 534038 553574 534274
rect 552954 514274 553574 534038
rect 552954 514038 552986 514274
rect 553222 514038 553306 514274
rect 553542 514038 553574 514274
rect 552954 494274 553574 514038
rect 552954 494038 552986 494274
rect 553222 494038 553306 494274
rect 553542 494038 553574 494274
rect 552954 474274 553574 494038
rect 552954 474038 552986 474274
rect 553222 474038 553306 474274
rect 553542 474038 553574 474274
rect 552954 454274 553574 474038
rect 552954 454038 552986 454274
rect 553222 454038 553306 454274
rect 553542 454038 553574 454274
rect 552954 434274 553574 454038
rect 552954 434038 552986 434274
rect 553222 434038 553306 434274
rect 553542 434038 553574 434274
rect 552954 421162 553574 434038
rect 555514 707718 556134 707750
rect 555514 707482 555546 707718
rect 555782 707482 555866 707718
rect 556102 707482 556134 707718
rect 555514 707398 556134 707482
rect 555514 707162 555546 707398
rect 555782 707162 555866 707398
rect 556102 707162 556134 707398
rect 555514 696954 556134 707162
rect 555514 696718 555546 696954
rect 555782 696718 555866 696954
rect 556102 696718 556134 696954
rect 555514 676954 556134 696718
rect 555514 676718 555546 676954
rect 555782 676718 555866 676954
rect 556102 676718 556134 676954
rect 555514 656954 556134 676718
rect 555514 656718 555546 656954
rect 555782 656718 555866 656954
rect 556102 656718 556134 656954
rect 555514 636954 556134 656718
rect 555514 636718 555546 636954
rect 555782 636718 555866 636954
rect 556102 636718 556134 636954
rect 555514 616954 556134 636718
rect 555514 616718 555546 616954
rect 555782 616718 555866 616954
rect 556102 616718 556134 616954
rect 555514 596954 556134 616718
rect 555514 596718 555546 596954
rect 555782 596718 555866 596954
rect 556102 596718 556134 596954
rect 555514 576954 556134 596718
rect 555514 576718 555546 576954
rect 555782 576718 555866 576954
rect 556102 576718 556134 576954
rect 555514 556954 556134 576718
rect 555514 556718 555546 556954
rect 555782 556718 555866 556954
rect 556102 556718 556134 556954
rect 555514 536954 556134 556718
rect 555514 536718 555546 536954
rect 555782 536718 555866 536954
rect 556102 536718 556134 536954
rect 555514 516954 556134 536718
rect 555514 516718 555546 516954
rect 555782 516718 555866 516954
rect 556102 516718 556134 516954
rect 555514 496954 556134 516718
rect 555514 496718 555546 496954
rect 555782 496718 555866 496954
rect 556102 496718 556134 496954
rect 555514 476954 556134 496718
rect 555514 476718 555546 476954
rect 555782 476718 555866 476954
rect 556102 476718 556134 476954
rect 555514 456954 556134 476718
rect 555514 456718 555546 456954
rect 555782 456718 555866 456954
rect 556102 456718 556134 456954
rect 555514 436954 556134 456718
rect 555514 436718 555546 436954
rect 555782 436718 555866 436954
rect 556102 436718 556134 436954
rect 555514 421162 556134 436718
rect 559234 700614 559854 709082
rect 559234 700378 559266 700614
rect 559502 700378 559586 700614
rect 559822 700378 559854 700614
rect 559234 680614 559854 700378
rect 559234 680378 559266 680614
rect 559502 680378 559586 680614
rect 559822 680378 559854 680614
rect 559234 660614 559854 680378
rect 559234 660378 559266 660614
rect 559502 660378 559586 660614
rect 559822 660378 559854 660614
rect 559234 640614 559854 660378
rect 559234 640378 559266 640614
rect 559502 640378 559586 640614
rect 559822 640378 559854 640614
rect 559234 620614 559854 640378
rect 559234 620378 559266 620614
rect 559502 620378 559586 620614
rect 559822 620378 559854 620614
rect 559234 600614 559854 620378
rect 559234 600378 559266 600614
rect 559502 600378 559586 600614
rect 559822 600378 559854 600614
rect 559234 580614 559854 600378
rect 559234 580378 559266 580614
rect 559502 580378 559586 580614
rect 559822 580378 559854 580614
rect 559234 560614 559854 580378
rect 559234 560378 559266 560614
rect 559502 560378 559586 560614
rect 559822 560378 559854 560614
rect 559234 540614 559854 560378
rect 559234 540378 559266 540614
rect 559502 540378 559586 540614
rect 559822 540378 559854 540614
rect 559234 520614 559854 540378
rect 559234 520378 559266 520614
rect 559502 520378 559586 520614
rect 559822 520378 559854 520614
rect 559234 500614 559854 520378
rect 559234 500378 559266 500614
rect 559502 500378 559586 500614
rect 559822 500378 559854 500614
rect 559234 480614 559854 500378
rect 559234 480378 559266 480614
rect 559502 480378 559586 480614
rect 559822 480378 559854 480614
rect 559234 460614 559854 480378
rect 559234 460378 559266 460614
rect 559502 460378 559586 460614
rect 559822 460378 559854 460614
rect 559234 440614 559854 460378
rect 559234 440378 559266 440614
rect 559502 440378 559586 440614
rect 559822 440378 559854 440614
rect 559234 420614 559854 440378
rect 559234 420378 559266 420614
rect 559502 420378 559586 420614
rect 559822 420378 559854 420614
rect 219568 413294 219888 413456
rect 219568 413058 219610 413294
rect 219846 413058 219888 413294
rect 219568 412896 219888 413058
rect 250288 413294 250608 413456
rect 250288 413058 250330 413294
rect 250566 413058 250608 413294
rect 250288 412896 250608 413058
rect 281008 413294 281328 413456
rect 281008 413058 281050 413294
rect 281286 413058 281328 413294
rect 281008 412896 281328 413058
rect 311728 413294 312048 413456
rect 311728 413058 311770 413294
rect 312006 413058 312048 413294
rect 311728 412896 312048 413058
rect 342448 413294 342768 413456
rect 342448 413058 342490 413294
rect 342726 413058 342768 413294
rect 342448 412896 342768 413058
rect 373168 413294 373488 413456
rect 373168 413058 373210 413294
rect 373446 413058 373488 413294
rect 373168 412896 373488 413058
rect 403888 413294 404208 413456
rect 403888 413058 403930 413294
rect 404166 413058 404208 413294
rect 403888 412896 404208 413058
rect 434608 413294 434928 413456
rect 434608 413058 434650 413294
rect 434886 413058 434928 413294
rect 434608 412896 434928 413058
rect 465328 413294 465648 413456
rect 465328 413058 465370 413294
rect 465606 413058 465648 413294
rect 465328 412896 465648 413058
rect 496048 413294 496368 413456
rect 496048 413058 496090 413294
rect 496326 413058 496368 413294
rect 496048 412896 496368 413058
rect 526768 413294 527088 413456
rect 526768 413058 526810 413294
rect 527046 413058 527088 413294
rect 526768 412896 527088 413058
rect 204208 403294 204528 403456
rect 204208 403058 204250 403294
rect 204486 403058 204528 403294
rect 204208 402896 204528 403058
rect 234928 403294 235248 403456
rect 234928 403058 234970 403294
rect 235206 403058 235248 403294
rect 234928 402896 235248 403058
rect 265648 403294 265968 403456
rect 265648 403058 265690 403294
rect 265926 403058 265968 403294
rect 265648 402896 265968 403058
rect 296368 403294 296688 403456
rect 296368 403058 296410 403294
rect 296646 403058 296688 403294
rect 296368 402896 296688 403058
rect 327088 403294 327408 403456
rect 327088 403058 327130 403294
rect 327366 403058 327408 403294
rect 327088 402896 327408 403058
rect 357808 403294 358128 403456
rect 357808 403058 357850 403294
rect 358086 403058 358128 403294
rect 357808 402896 358128 403058
rect 388528 403294 388848 403456
rect 388528 403058 388570 403294
rect 388806 403058 388848 403294
rect 388528 402896 388848 403058
rect 419248 403294 419568 403456
rect 419248 403058 419290 403294
rect 419526 403058 419568 403294
rect 419248 402896 419568 403058
rect 449968 403294 450288 403456
rect 449968 403058 450010 403294
rect 450246 403058 450288 403294
rect 449968 402896 450288 403058
rect 480688 403294 481008 403456
rect 480688 403058 480730 403294
rect 480966 403058 481008 403294
rect 480688 402896 481008 403058
rect 511408 403294 511728 403456
rect 511408 403058 511450 403294
rect 511686 403058 511728 403294
rect 511408 402896 511728 403058
rect 542128 403294 542448 403456
rect 542128 403058 542170 403294
rect 542406 403058 542448 403294
rect 542128 402896 542448 403058
rect 559234 400614 559854 420378
rect 559234 400378 559266 400614
rect 559502 400378 559586 400614
rect 559822 400378 559854 400614
rect 219568 393294 219888 393456
rect 219568 393058 219610 393294
rect 219846 393058 219888 393294
rect 219568 392896 219888 393058
rect 250288 393294 250608 393456
rect 250288 393058 250330 393294
rect 250566 393058 250608 393294
rect 250288 392896 250608 393058
rect 281008 393294 281328 393456
rect 281008 393058 281050 393294
rect 281286 393058 281328 393294
rect 281008 392896 281328 393058
rect 311728 393294 312048 393456
rect 311728 393058 311770 393294
rect 312006 393058 312048 393294
rect 311728 392896 312048 393058
rect 342448 393294 342768 393456
rect 342448 393058 342490 393294
rect 342726 393058 342768 393294
rect 342448 392896 342768 393058
rect 373168 393294 373488 393456
rect 373168 393058 373210 393294
rect 373446 393058 373488 393294
rect 373168 392896 373488 393058
rect 403888 393294 404208 393456
rect 403888 393058 403930 393294
rect 404166 393058 404208 393294
rect 403888 392896 404208 393058
rect 434608 393294 434928 393456
rect 434608 393058 434650 393294
rect 434886 393058 434928 393294
rect 434608 392896 434928 393058
rect 465328 393294 465648 393456
rect 465328 393058 465370 393294
rect 465606 393058 465648 393294
rect 465328 392896 465648 393058
rect 496048 393294 496368 393456
rect 496048 393058 496090 393294
rect 496326 393058 496368 393294
rect 496048 392896 496368 393058
rect 526768 393294 527088 393456
rect 526768 393058 526810 393294
rect 527046 393058 527088 393294
rect 526768 392896 527088 393058
rect 204208 383294 204528 383456
rect 204208 383058 204250 383294
rect 204486 383058 204528 383294
rect 204208 382896 204528 383058
rect 234928 383294 235248 383456
rect 234928 383058 234970 383294
rect 235206 383058 235248 383294
rect 234928 382896 235248 383058
rect 265648 383294 265968 383456
rect 265648 383058 265690 383294
rect 265926 383058 265968 383294
rect 265648 382896 265968 383058
rect 296368 383294 296688 383456
rect 296368 383058 296410 383294
rect 296646 383058 296688 383294
rect 296368 382896 296688 383058
rect 327088 383294 327408 383456
rect 327088 383058 327130 383294
rect 327366 383058 327408 383294
rect 327088 382896 327408 383058
rect 357808 383294 358128 383456
rect 357808 383058 357850 383294
rect 358086 383058 358128 383294
rect 357808 382896 358128 383058
rect 388528 383294 388848 383456
rect 388528 383058 388570 383294
rect 388806 383058 388848 383294
rect 388528 382896 388848 383058
rect 419248 383294 419568 383456
rect 419248 383058 419290 383294
rect 419526 383058 419568 383294
rect 419248 382896 419568 383058
rect 449968 383294 450288 383456
rect 449968 383058 450010 383294
rect 450246 383058 450288 383294
rect 449968 382896 450288 383058
rect 480688 383294 481008 383456
rect 480688 383058 480730 383294
rect 480966 383058 481008 383294
rect 480688 382896 481008 383058
rect 511408 383294 511728 383456
rect 511408 383058 511450 383294
rect 511686 383058 511728 383294
rect 511408 382896 511728 383058
rect 542128 383294 542448 383456
rect 542128 383058 542170 383294
rect 542406 383058 542448 383294
rect 542128 382896 542448 383058
rect 559234 380614 559854 400378
rect 559234 380378 559266 380614
rect 559502 380378 559586 380614
rect 559822 380378 559854 380614
rect 219568 373294 219888 373456
rect 219568 373058 219610 373294
rect 219846 373058 219888 373294
rect 219568 372896 219888 373058
rect 250288 373294 250608 373456
rect 250288 373058 250330 373294
rect 250566 373058 250608 373294
rect 250288 372896 250608 373058
rect 281008 373294 281328 373456
rect 281008 373058 281050 373294
rect 281286 373058 281328 373294
rect 281008 372896 281328 373058
rect 311728 373294 312048 373456
rect 311728 373058 311770 373294
rect 312006 373058 312048 373294
rect 311728 372896 312048 373058
rect 342448 373294 342768 373456
rect 342448 373058 342490 373294
rect 342726 373058 342768 373294
rect 342448 372896 342768 373058
rect 373168 373294 373488 373456
rect 373168 373058 373210 373294
rect 373446 373058 373488 373294
rect 373168 372896 373488 373058
rect 403888 373294 404208 373456
rect 403888 373058 403930 373294
rect 404166 373058 404208 373294
rect 403888 372896 404208 373058
rect 434608 373294 434928 373456
rect 434608 373058 434650 373294
rect 434886 373058 434928 373294
rect 434608 372896 434928 373058
rect 465328 373294 465648 373456
rect 465328 373058 465370 373294
rect 465606 373058 465648 373294
rect 465328 372896 465648 373058
rect 496048 373294 496368 373456
rect 496048 373058 496090 373294
rect 496326 373058 496368 373294
rect 496048 372896 496368 373058
rect 526768 373294 527088 373456
rect 526768 373058 526810 373294
rect 527046 373058 527088 373294
rect 526768 372896 527088 373058
rect 204208 363294 204528 363456
rect 204208 363058 204250 363294
rect 204486 363058 204528 363294
rect 204208 362896 204528 363058
rect 234928 363294 235248 363456
rect 234928 363058 234970 363294
rect 235206 363058 235248 363294
rect 234928 362896 235248 363058
rect 265648 363294 265968 363456
rect 265648 363058 265690 363294
rect 265926 363058 265968 363294
rect 265648 362896 265968 363058
rect 296368 363294 296688 363456
rect 296368 363058 296410 363294
rect 296646 363058 296688 363294
rect 296368 362896 296688 363058
rect 327088 363294 327408 363456
rect 327088 363058 327130 363294
rect 327366 363058 327408 363294
rect 327088 362896 327408 363058
rect 357808 363294 358128 363456
rect 357808 363058 357850 363294
rect 358086 363058 358128 363294
rect 357808 362896 358128 363058
rect 388528 363294 388848 363456
rect 388528 363058 388570 363294
rect 388806 363058 388848 363294
rect 388528 362896 388848 363058
rect 419248 363294 419568 363456
rect 419248 363058 419290 363294
rect 419526 363058 419568 363294
rect 419248 362896 419568 363058
rect 449968 363294 450288 363456
rect 449968 363058 450010 363294
rect 450246 363058 450288 363294
rect 449968 362896 450288 363058
rect 480688 363294 481008 363456
rect 480688 363058 480730 363294
rect 480966 363058 481008 363294
rect 480688 362896 481008 363058
rect 511408 363294 511728 363456
rect 511408 363058 511450 363294
rect 511686 363058 511728 363294
rect 511408 362896 511728 363058
rect 542128 363294 542448 363456
rect 542128 363058 542170 363294
rect 542406 363058 542448 363294
rect 542128 362896 542448 363058
rect 559234 360614 559854 380378
rect 559234 360378 559266 360614
rect 559502 360378 559586 360614
rect 559822 360378 559854 360614
rect 219568 353294 219888 353456
rect 219568 353058 219610 353294
rect 219846 353058 219888 353294
rect 219568 352896 219888 353058
rect 250288 353294 250608 353456
rect 250288 353058 250330 353294
rect 250566 353058 250608 353294
rect 250288 352896 250608 353058
rect 281008 353294 281328 353456
rect 281008 353058 281050 353294
rect 281286 353058 281328 353294
rect 281008 352896 281328 353058
rect 311728 353294 312048 353456
rect 311728 353058 311770 353294
rect 312006 353058 312048 353294
rect 311728 352896 312048 353058
rect 342448 353294 342768 353456
rect 342448 353058 342490 353294
rect 342726 353058 342768 353294
rect 342448 352896 342768 353058
rect 373168 353294 373488 353456
rect 373168 353058 373210 353294
rect 373446 353058 373488 353294
rect 373168 352896 373488 353058
rect 403888 353294 404208 353456
rect 403888 353058 403930 353294
rect 404166 353058 404208 353294
rect 403888 352896 404208 353058
rect 434608 353294 434928 353456
rect 434608 353058 434650 353294
rect 434886 353058 434928 353294
rect 434608 352896 434928 353058
rect 465328 353294 465648 353456
rect 465328 353058 465370 353294
rect 465606 353058 465648 353294
rect 465328 352896 465648 353058
rect 496048 353294 496368 353456
rect 496048 353058 496090 353294
rect 496326 353058 496368 353294
rect 496048 352896 496368 353058
rect 526768 353294 527088 353456
rect 526768 353058 526810 353294
rect 527046 353058 527088 353294
rect 526768 352896 527088 353058
rect 204208 343294 204528 343456
rect 204208 343058 204250 343294
rect 204486 343058 204528 343294
rect 204208 342896 204528 343058
rect 234928 343294 235248 343456
rect 234928 343058 234970 343294
rect 235206 343058 235248 343294
rect 234928 342896 235248 343058
rect 265648 343294 265968 343456
rect 265648 343058 265690 343294
rect 265926 343058 265968 343294
rect 265648 342896 265968 343058
rect 296368 343294 296688 343456
rect 296368 343058 296410 343294
rect 296646 343058 296688 343294
rect 296368 342896 296688 343058
rect 327088 343294 327408 343456
rect 327088 343058 327130 343294
rect 327366 343058 327408 343294
rect 327088 342896 327408 343058
rect 357808 343294 358128 343456
rect 357808 343058 357850 343294
rect 358086 343058 358128 343294
rect 357808 342896 358128 343058
rect 388528 343294 388848 343456
rect 388528 343058 388570 343294
rect 388806 343058 388848 343294
rect 388528 342896 388848 343058
rect 419248 343294 419568 343456
rect 419248 343058 419290 343294
rect 419526 343058 419568 343294
rect 419248 342896 419568 343058
rect 449968 343294 450288 343456
rect 449968 343058 450010 343294
rect 450246 343058 450288 343294
rect 449968 342896 450288 343058
rect 480688 343294 481008 343456
rect 480688 343058 480730 343294
rect 480966 343058 481008 343294
rect 480688 342896 481008 343058
rect 511408 343294 511728 343456
rect 511408 343058 511450 343294
rect 511686 343058 511728 343294
rect 511408 342896 511728 343058
rect 542128 343294 542448 343456
rect 542128 343058 542170 343294
rect 542406 343058 542448 343294
rect 542128 342896 542448 343058
rect 559234 340614 559854 360378
rect 559234 340378 559266 340614
rect 559502 340378 559586 340614
rect 559822 340378 559854 340614
rect 219568 333294 219888 333456
rect 219568 333058 219610 333294
rect 219846 333058 219888 333294
rect 219568 332896 219888 333058
rect 250288 333294 250608 333456
rect 250288 333058 250330 333294
rect 250566 333058 250608 333294
rect 250288 332896 250608 333058
rect 281008 333294 281328 333456
rect 281008 333058 281050 333294
rect 281286 333058 281328 333294
rect 281008 332896 281328 333058
rect 311728 333294 312048 333456
rect 311728 333058 311770 333294
rect 312006 333058 312048 333294
rect 311728 332896 312048 333058
rect 342448 333294 342768 333456
rect 342448 333058 342490 333294
rect 342726 333058 342768 333294
rect 342448 332896 342768 333058
rect 373168 333294 373488 333456
rect 373168 333058 373210 333294
rect 373446 333058 373488 333294
rect 373168 332896 373488 333058
rect 403888 333294 404208 333456
rect 403888 333058 403930 333294
rect 404166 333058 404208 333294
rect 403888 332896 404208 333058
rect 434608 333294 434928 333456
rect 434608 333058 434650 333294
rect 434886 333058 434928 333294
rect 434608 332896 434928 333058
rect 465328 333294 465648 333456
rect 465328 333058 465370 333294
rect 465606 333058 465648 333294
rect 465328 332896 465648 333058
rect 496048 333294 496368 333456
rect 496048 333058 496090 333294
rect 496326 333058 496368 333294
rect 496048 332896 496368 333058
rect 526768 333294 527088 333456
rect 526768 333058 526810 333294
rect 527046 333058 527088 333294
rect 526768 332896 527088 333058
rect 204208 323294 204528 323456
rect 204208 323058 204250 323294
rect 204486 323058 204528 323294
rect 204208 322896 204528 323058
rect 234928 323294 235248 323456
rect 234928 323058 234970 323294
rect 235206 323058 235248 323294
rect 234928 322896 235248 323058
rect 265648 323294 265968 323456
rect 265648 323058 265690 323294
rect 265926 323058 265968 323294
rect 265648 322896 265968 323058
rect 296368 323294 296688 323456
rect 296368 323058 296410 323294
rect 296646 323058 296688 323294
rect 296368 322896 296688 323058
rect 327088 323294 327408 323456
rect 327088 323058 327130 323294
rect 327366 323058 327408 323294
rect 327088 322896 327408 323058
rect 357808 323294 358128 323456
rect 357808 323058 357850 323294
rect 358086 323058 358128 323294
rect 357808 322896 358128 323058
rect 388528 323294 388848 323456
rect 388528 323058 388570 323294
rect 388806 323058 388848 323294
rect 388528 322896 388848 323058
rect 419248 323294 419568 323456
rect 419248 323058 419290 323294
rect 419526 323058 419568 323294
rect 419248 322896 419568 323058
rect 449968 323294 450288 323456
rect 449968 323058 450010 323294
rect 450246 323058 450288 323294
rect 449968 322896 450288 323058
rect 480688 323294 481008 323456
rect 480688 323058 480730 323294
rect 480966 323058 481008 323294
rect 480688 322896 481008 323058
rect 511408 323294 511728 323456
rect 511408 323058 511450 323294
rect 511686 323058 511728 323294
rect 511408 322896 511728 323058
rect 542128 323294 542448 323456
rect 542128 323058 542170 323294
rect 542406 323058 542448 323294
rect 542128 322896 542448 323058
rect 559234 320614 559854 340378
rect 559234 320378 559266 320614
rect 559502 320378 559586 320614
rect 559822 320378 559854 320614
rect 219568 313294 219888 313456
rect 219568 313058 219610 313294
rect 219846 313058 219888 313294
rect 219568 312896 219888 313058
rect 250288 313294 250608 313456
rect 250288 313058 250330 313294
rect 250566 313058 250608 313294
rect 250288 312896 250608 313058
rect 281008 313294 281328 313456
rect 281008 313058 281050 313294
rect 281286 313058 281328 313294
rect 281008 312896 281328 313058
rect 311728 313294 312048 313456
rect 311728 313058 311770 313294
rect 312006 313058 312048 313294
rect 311728 312896 312048 313058
rect 342448 313294 342768 313456
rect 342448 313058 342490 313294
rect 342726 313058 342768 313294
rect 342448 312896 342768 313058
rect 373168 313294 373488 313456
rect 373168 313058 373210 313294
rect 373446 313058 373488 313294
rect 373168 312896 373488 313058
rect 403888 313294 404208 313456
rect 403888 313058 403930 313294
rect 404166 313058 404208 313294
rect 403888 312896 404208 313058
rect 434608 313294 434928 313456
rect 434608 313058 434650 313294
rect 434886 313058 434928 313294
rect 434608 312896 434928 313058
rect 465328 313294 465648 313456
rect 465328 313058 465370 313294
rect 465606 313058 465648 313294
rect 465328 312896 465648 313058
rect 496048 313294 496368 313456
rect 496048 313058 496090 313294
rect 496326 313058 496368 313294
rect 496048 312896 496368 313058
rect 526768 313294 527088 313456
rect 526768 313058 526810 313294
rect 527046 313058 527088 313294
rect 526768 312896 527088 313058
rect 204208 303294 204528 303456
rect 204208 303058 204250 303294
rect 204486 303058 204528 303294
rect 204208 302896 204528 303058
rect 234928 303294 235248 303456
rect 234928 303058 234970 303294
rect 235206 303058 235248 303294
rect 234928 302896 235248 303058
rect 265648 303294 265968 303456
rect 265648 303058 265690 303294
rect 265926 303058 265968 303294
rect 265648 302896 265968 303058
rect 296368 303294 296688 303456
rect 296368 303058 296410 303294
rect 296646 303058 296688 303294
rect 296368 302896 296688 303058
rect 327088 303294 327408 303456
rect 327088 303058 327130 303294
rect 327366 303058 327408 303294
rect 327088 302896 327408 303058
rect 357808 303294 358128 303456
rect 357808 303058 357850 303294
rect 358086 303058 358128 303294
rect 357808 302896 358128 303058
rect 388528 303294 388848 303456
rect 388528 303058 388570 303294
rect 388806 303058 388848 303294
rect 388528 302896 388848 303058
rect 419248 303294 419568 303456
rect 419248 303058 419290 303294
rect 419526 303058 419568 303294
rect 419248 302896 419568 303058
rect 449968 303294 450288 303456
rect 449968 303058 450010 303294
rect 450246 303058 450288 303294
rect 449968 302896 450288 303058
rect 480688 303294 481008 303456
rect 480688 303058 480730 303294
rect 480966 303058 481008 303294
rect 480688 302896 481008 303058
rect 511408 303294 511728 303456
rect 511408 303058 511450 303294
rect 511686 303058 511728 303294
rect 511408 302896 511728 303058
rect 542128 303294 542448 303456
rect 542128 303058 542170 303294
rect 542406 303058 542448 303294
rect 542128 302896 542448 303058
rect 559234 300614 559854 320378
rect 559234 300378 559266 300614
rect 559502 300378 559586 300614
rect 559822 300378 559854 300614
rect 219568 293294 219888 293456
rect 219568 293058 219610 293294
rect 219846 293058 219888 293294
rect 219568 292896 219888 293058
rect 250288 293294 250608 293456
rect 250288 293058 250330 293294
rect 250566 293058 250608 293294
rect 250288 292896 250608 293058
rect 281008 293294 281328 293456
rect 281008 293058 281050 293294
rect 281286 293058 281328 293294
rect 281008 292896 281328 293058
rect 311728 293294 312048 293456
rect 311728 293058 311770 293294
rect 312006 293058 312048 293294
rect 311728 292896 312048 293058
rect 342448 293294 342768 293456
rect 342448 293058 342490 293294
rect 342726 293058 342768 293294
rect 342448 292896 342768 293058
rect 373168 293294 373488 293456
rect 373168 293058 373210 293294
rect 373446 293058 373488 293294
rect 373168 292896 373488 293058
rect 403888 293294 404208 293456
rect 403888 293058 403930 293294
rect 404166 293058 404208 293294
rect 403888 292896 404208 293058
rect 434608 293294 434928 293456
rect 434608 293058 434650 293294
rect 434886 293058 434928 293294
rect 434608 292896 434928 293058
rect 465328 293294 465648 293456
rect 465328 293058 465370 293294
rect 465606 293058 465648 293294
rect 465328 292896 465648 293058
rect 496048 293294 496368 293456
rect 496048 293058 496090 293294
rect 496326 293058 496368 293294
rect 496048 292896 496368 293058
rect 526768 293294 527088 293456
rect 526768 293058 526810 293294
rect 527046 293058 527088 293294
rect 526768 292896 527088 293058
rect 204208 283294 204528 283456
rect 204208 283058 204250 283294
rect 204486 283058 204528 283294
rect 204208 282896 204528 283058
rect 234928 283294 235248 283456
rect 234928 283058 234970 283294
rect 235206 283058 235248 283294
rect 234928 282896 235248 283058
rect 265648 283294 265968 283456
rect 265648 283058 265690 283294
rect 265926 283058 265968 283294
rect 265648 282896 265968 283058
rect 296368 283294 296688 283456
rect 296368 283058 296410 283294
rect 296646 283058 296688 283294
rect 296368 282896 296688 283058
rect 327088 283294 327408 283456
rect 327088 283058 327130 283294
rect 327366 283058 327408 283294
rect 327088 282896 327408 283058
rect 357808 283294 358128 283456
rect 357808 283058 357850 283294
rect 358086 283058 358128 283294
rect 357808 282896 358128 283058
rect 388528 283294 388848 283456
rect 388528 283058 388570 283294
rect 388806 283058 388848 283294
rect 388528 282896 388848 283058
rect 419248 283294 419568 283456
rect 419248 283058 419290 283294
rect 419526 283058 419568 283294
rect 419248 282896 419568 283058
rect 449968 283294 450288 283456
rect 449968 283058 450010 283294
rect 450246 283058 450288 283294
rect 449968 282896 450288 283058
rect 480688 283294 481008 283456
rect 480688 283058 480730 283294
rect 480966 283058 481008 283294
rect 480688 282896 481008 283058
rect 511408 283294 511728 283456
rect 511408 283058 511450 283294
rect 511686 283058 511728 283294
rect 511408 282896 511728 283058
rect 542128 283294 542448 283456
rect 542128 283058 542170 283294
rect 542406 283058 542448 283294
rect 542128 282896 542448 283058
rect 559234 280614 559854 300378
rect 559234 280378 559266 280614
rect 559502 280378 559586 280614
rect 559822 280378 559854 280614
rect 219568 273294 219888 273456
rect 219568 273058 219610 273294
rect 219846 273058 219888 273294
rect 219568 272896 219888 273058
rect 250288 273294 250608 273456
rect 250288 273058 250330 273294
rect 250566 273058 250608 273294
rect 250288 272896 250608 273058
rect 281008 273294 281328 273456
rect 281008 273058 281050 273294
rect 281286 273058 281328 273294
rect 281008 272896 281328 273058
rect 311728 273294 312048 273456
rect 311728 273058 311770 273294
rect 312006 273058 312048 273294
rect 311728 272896 312048 273058
rect 342448 273294 342768 273456
rect 342448 273058 342490 273294
rect 342726 273058 342768 273294
rect 342448 272896 342768 273058
rect 373168 273294 373488 273456
rect 373168 273058 373210 273294
rect 373446 273058 373488 273294
rect 373168 272896 373488 273058
rect 403888 273294 404208 273456
rect 403888 273058 403930 273294
rect 404166 273058 404208 273294
rect 403888 272896 404208 273058
rect 434608 273294 434928 273456
rect 434608 273058 434650 273294
rect 434886 273058 434928 273294
rect 434608 272896 434928 273058
rect 465328 273294 465648 273456
rect 465328 273058 465370 273294
rect 465606 273058 465648 273294
rect 465328 272896 465648 273058
rect 496048 273294 496368 273456
rect 496048 273058 496090 273294
rect 496326 273058 496368 273294
rect 496048 272896 496368 273058
rect 526768 273294 527088 273456
rect 526768 273058 526810 273294
rect 527046 273058 527088 273294
rect 526768 272896 527088 273058
rect 204208 263294 204528 263456
rect 204208 263058 204250 263294
rect 204486 263058 204528 263294
rect 204208 262896 204528 263058
rect 234928 263294 235248 263456
rect 234928 263058 234970 263294
rect 235206 263058 235248 263294
rect 234928 262896 235248 263058
rect 265648 263294 265968 263456
rect 265648 263058 265690 263294
rect 265926 263058 265968 263294
rect 265648 262896 265968 263058
rect 296368 263294 296688 263456
rect 296368 263058 296410 263294
rect 296646 263058 296688 263294
rect 296368 262896 296688 263058
rect 327088 263294 327408 263456
rect 327088 263058 327130 263294
rect 327366 263058 327408 263294
rect 327088 262896 327408 263058
rect 357808 263294 358128 263456
rect 357808 263058 357850 263294
rect 358086 263058 358128 263294
rect 357808 262896 358128 263058
rect 388528 263294 388848 263456
rect 388528 263058 388570 263294
rect 388806 263058 388848 263294
rect 388528 262896 388848 263058
rect 419248 263294 419568 263456
rect 419248 263058 419290 263294
rect 419526 263058 419568 263294
rect 419248 262896 419568 263058
rect 449968 263294 450288 263456
rect 449968 263058 450010 263294
rect 450246 263058 450288 263294
rect 449968 262896 450288 263058
rect 480688 263294 481008 263456
rect 480688 263058 480730 263294
rect 480966 263058 481008 263294
rect 480688 262896 481008 263058
rect 511408 263294 511728 263456
rect 511408 263058 511450 263294
rect 511686 263058 511728 263294
rect 511408 262896 511728 263058
rect 542128 263294 542448 263456
rect 542128 263058 542170 263294
rect 542406 263058 542448 263294
rect 542128 262896 542448 263058
rect 559234 260614 559854 280378
rect 559234 260378 559266 260614
rect 559502 260378 559586 260614
rect 559822 260378 559854 260614
rect 219568 253294 219888 253456
rect 219568 253058 219610 253294
rect 219846 253058 219888 253294
rect 219568 252896 219888 253058
rect 250288 253294 250608 253456
rect 250288 253058 250330 253294
rect 250566 253058 250608 253294
rect 250288 252896 250608 253058
rect 281008 253294 281328 253456
rect 281008 253058 281050 253294
rect 281286 253058 281328 253294
rect 281008 252896 281328 253058
rect 311728 253294 312048 253456
rect 311728 253058 311770 253294
rect 312006 253058 312048 253294
rect 311728 252896 312048 253058
rect 342448 253294 342768 253456
rect 342448 253058 342490 253294
rect 342726 253058 342768 253294
rect 342448 252896 342768 253058
rect 373168 253294 373488 253456
rect 373168 253058 373210 253294
rect 373446 253058 373488 253294
rect 373168 252896 373488 253058
rect 403888 253294 404208 253456
rect 403888 253058 403930 253294
rect 404166 253058 404208 253294
rect 403888 252896 404208 253058
rect 434608 253294 434928 253456
rect 434608 253058 434650 253294
rect 434886 253058 434928 253294
rect 434608 252896 434928 253058
rect 465328 253294 465648 253456
rect 465328 253058 465370 253294
rect 465606 253058 465648 253294
rect 465328 252896 465648 253058
rect 496048 253294 496368 253456
rect 496048 253058 496090 253294
rect 496326 253058 496368 253294
rect 496048 252896 496368 253058
rect 526768 253294 527088 253456
rect 526768 253058 526810 253294
rect 527046 253058 527088 253294
rect 526768 252896 527088 253058
rect 198779 248028 198845 248029
rect 198779 247964 198780 248028
rect 198844 247964 198845 248028
rect 198779 247963 198845 247964
rect 204208 243294 204528 243456
rect 204208 243058 204250 243294
rect 204486 243058 204528 243294
rect 204208 242896 204528 243058
rect 234928 243294 235248 243456
rect 234928 243058 234970 243294
rect 235206 243058 235248 243294
rect 234928 242896 235248 243058
rect 265648 243294 265968 243456
rect 265648 243058 265690 243294
rect 265926 243058 265968 243294
rect 265648 242896 265968 243058
rect 296368 243294 296688 243456
rect 296368 243058 296410 243294
rect 296646 243058 296688 243294
rect 296368 242896 296688 243058
rect 327088 243294 327408 243456
rect 327088 243058 327130 243294
rect 327366 243058 327408 243294
rect 327088 242896 327408 243058
rect 357808 243294 358128 243456
rect 357808 243058 357850 243294
rect 358086 243058 358128 243294
rect 357808 242896 358128 243058
rect 388528 243294 388848 243456
rect 388528 243058 388570 243294
rect 388806 243058 388848 243294
rect 388528 242896 388848 243058
rect 419248 243294 419568 243456
rect 419248 243058 419290 243294
rect 419526 243058 419568 243294
rect 419248 242896 419568 243058
rect 449968 243294 450288 243456
rect 449968 243058 450010 243294
rect 450246 243058 450288 243294
rect 449968 242896 450288 243058
rect 480688 243294 481008 243456
rect 480688 243058 480730 243294
rect 480966 243058 481008 243294
rect 480688 242896 481008 243058
rect 511408 243294 511728 243456
rect 511408 243058 511450 243294
rect 511686 243058 511728 243294
rect 511408 242896 511728 243058
rect 542128 243294 542448 243456
rect 542128 243058 542170 243294
rect 542406 243058 542448 243294
rect 542128 242896 542448 243058
rect 195514 236718 195546 236954
rect 195782 236718 195866 236954
rect 196102 236718 196134 236954
rect 195514 216954 196134 236718
rect 559234 240614 559854 260378
rect 559234 240378 559266 240614
rect 559502 240378 559586 240614
rect 559822 240378 559854 240614
rect 219568 233294 219888 233456
rect 219568 233058 219610 233294
rect 219846 233058 219888 233294
rect 219568 232896 219888 233058
rect 250288 233294 250608 233456
rect 250288 233058 250330 233294
rect 250566 233058 250608 233294
rect 250288 232896 250608 233058
rect 281008 233294 281328 233456
rect 281008 233058 281050 233294
rect 281286 233058 281328 233294
rect 281008 232896 281328 233058
rect 311728 233294 312048 233456
rect 311728 233058 311770 233294
rect 312006 233058 312048 233294
rect 311728 232896 312048 233058
rect 342448 233294 342768 233456
rect 342448 233058 342490 233294
rect 342726 233058 342768 233294
rect 342448 232896 342768 233058
rect 373168 233294 373488 233456
rect 373168 233058 373210 233294
rect 373446 233058 373488 233294
rect 373168 232896 373488 233058
rect 403888 233294 404208 233456
rect 403888 233058 403930 233294
rect 404166 233058 404208 233294
rect 403888 232896 404208 233058
rect 434608 233294 434928 233456
rect 434608 233058 434650 233294
rect 434886 233058 434928 233294
rect 434608 232896 434928 233058
rect 465328 233294 465648 233456
rect 465328 233058 465370 233294
rect 465606 233058 465648 233294
rect 465328 232896 465648 233058
rect 496048 233294 496368 233456
rect 496048 233058 496090 233294
rect 496326 233058 496368 233294
rect 496048 232896 496368 233058
rect 526768 233294 527088 233456
rect 526768 233058 526810 233294
rect 527046 233058 527088 233294
rect 526768 232896 527088 233058
rect 204208 223294 204528 223456
rect 204208 223058 204250 223294
rect 204486 223058 204528 223294
rect 204208 222896 204528 223058
rect 234928 223294 235248 223456
rect 234928 223058 234970 223294
rect 235206 223058 235248 223294
rect 234928 222896 235248 223058
rect 265648 223294 265968 223456
rect 265648 223058 265690 223294
rect 265926 223058 265968 223294
rect 265648 222896 265968 223058
rect 296368 223294 296688 223456
rect 296368 223058 296410 223294
rect 296646 223058 296688 223294
rect 296368 222896 296688 223058
rect 327088 223294 327408 223456
rect 327088 223058 327130 223294
rect 327366 223058 327408 223294
rect 327088 222896 327408 223058
rect 357808 223294 358128 223456
rect 357808 223058 357850 223294
rect 358086 223058 358128 223294
rect 357808 222896 358128 223058
rect 388528 223294 388848 223456
rect 388528 223058 388570 223294
rect 388806 223058 388848 223294
rect 388528 222896 388848 223058
rect 419248 223294 419568 223456
rect 419248 223058 419290 223294
rect 419526 223058 419568 223294
rect 419248 222896 419568 223058
rect 449968 223294 450288 223456
rect 449968 223058 450010 223294
rect 450246 223058 450288 223294
rect 449968 222896 450288 223058
rect 480688 223294 481008 223456
rect 480688 223058 480730 223294
rect 480966 223058 481008 223294
rect 480688 222896 481008 223058
rect 511408 223294 511728 223456
rect 511408 223058 511450 223294
rect 511686 223058 511728 223294
rect 511408 222896 511728 223058
rect 542128 223294 542448 223456
rect 542128 223058 542170 223294
rect 542406 223058 542448 223294
rect 542128 222896 542448 223058
rect 195514 216718 195546 216954
rect 195782 216718 195866 216954
rect 196102 216718 196134 216954
rect 195514 196954 196134 216718
rect 559234 220614 559854 240378
rect 559234 220378 559266 220614
rect 559502 220378 559586 220614
rect 559822 220378 559854 220614
rect 219568 213294 219888 213456
rect 219568 213058 219610 213294
rect 219846 213058 219888 213294
rect 219568 212896 219888 213058
rect 250288 213294 250608 213456
rect 250288 213058 250330 213294
rect 250566 213058 250608 213294
rect 250288 212896 250608 213058
rect 281008 213294 281328 213456
rect 281008 213058 281050 213294
rect 281286 213058 281328 213294
rect 281008 212896 281328 213058
rect 311728 213294 312048 213456
rect 311728 213058 311770 213294
rect 312006 213058 312048 213294
rect 311728 212896 312048 213058
rect 342448 213294 342768 213456
rect 342448 213058 342490 213294
rect 342726 213058 342768 213294
rect 342448 212896 342768 213058
rect 373168 213294 373488 213456
rect 373168 213058 373210 213294
rect 373446 213058 373488 213294
rect 373168 212896 373488 213058
rect 403888 213294 404208 213456
rect 403888 213058 403930 213294
rect 404166 213058 404208 213294
rect 403888 212896 404208 213058
rect 434608 213294 434928 213456
rect 434608 213058 434650 213294
rect 434886 213058 434928 213294
rect 434608 212896 434928 213058
rect 465328 213294 465648 213456
rect 465328 213058 465370 213294
rect 465606 213058 465648 213294
rect 465328 212896 465648 213058
rect 496048 213294 496368 213456
rect 496048 213058 496090 213294
rect 496326 213058 496368 213294
rect 496048 212896 496368 213058
rect 526768 213294 527088 213456
rect 526768 213058 526810 213294
rect 527046 213058 527088 213294
rect 526768 212896 527088 213058
rect 204208 203294 204528 203456
rect 204208 203058 204250 203294
rect 204486 203058 204528 203294
rect 204208 202896 204528 203058
rect 234928 203294 235248 203456
rect 234928 203058 234970 203294
rect 235206 203058 235248 203294
rect 234928 202896 235248 203058
rect 265648 203294 265968 203456
rect 265648 203058 265690 203294
rect 265926 203058 265968 203294
rect 265648 202896 265968 203058
rect 296368 203294 296688 203456
rect 296368 203058 296410 203294
rect 296646 203058 296688 203294
rect 296368 202896 296688 203058
rect 327088 203294 327408 203456
rect 327088 203058 327130 203294
rect 327366 203058 327408 203294
rect 327088 202896 327408 203058
rect 357808 203294 358128 203456
rect 357808 203058 357850 203294
rect 358086 203058 358128 203294
rect 357808 202896 358128 203058
rect 388528 203294 388848 203456
rect 388528 203058 388570 203294
rect 388806 203058 388848 203294
rect 388528 202896 388848 203058
rect 419248 203294 419568 203456
rect 419248 203058 419290 203294
rect 419526 203058 419568 203294
rect 419248 202896 419568 203058
rect 449968 203294 450288 203456
rect 449968 203058 450010 203294
rect 450246 203058 450288 203294
rect 449968 202896 450288 203058
rect 480688 203294 481008 203456
rect 480688 203058 480730 203294
rect 480966 203058 481008 203294
rect 480688 202896 481008 203058
rect 511408 203294 511728 203456
rect 511408 203058 511450 203294
rect 511686 203058 511728 203294
rect 511408 202896 511728 203058
rect 542128 203294 542448 203456
rect 542128 203058 542170 203294
rect 542406 203058 542448 203294
rect 542128 202896 542448 203058
rect 195514 196718 195546 196954
rect 195782 196718 195866 196954
rect 196102 196718 196134 196954
rect 195514 176954 196134 196718
rect 559234 200614 559854 220378
rect 559234 200378 559266 200614
rect 559502 200378 559586 200614
rect 559822 200378 559854 200614
rect 219568 193294 219888 193456
rect 219568 193058 219610 193294
rect 219846 193058 219888 193294
rect 219568 192896 219888 193058
rect 250288 193294 250608 193456
rect 250288 193058 250330 193294
rect 250566 193058 250608 193294
rect 250288 192896 250608 193058
rect 281008 193294 281328 193456
rect 281008 193058 281050 193294
rect 281286 193058 281328 193294
rect 281008 192896 281328 193058
rect 311728 193294 312048 193456
rect 311728 193058 311770 193294
rect 312006 193058 312048 193294
rect 311728 192896 312048 193058
rect 342448 193294 342768 193456
rect 342448 193058 342490 193294
rect 342726 193058 342768 193294
rect 342448 192896 342768 193058
rect 373168 193294 373488 193456
rect 373168 193058 373210 193294
rect 373446 193058 373488 193294
rect 373168 192896 373488 193058
rect 403888 193294 404208 193456
rect 403888 193058 403930 193294
rect 404166 193058 404208 193294
rect 403888 192896 404208 193058
rect 434608 193294 434928 193456
rect 434608 193058 434650 193294
rect 434886 193058 434928 193294
rect 434608 192896 434928 193058
rect 465328 193294 465648 193456
rect 465328 193058 465370 193294
rect 465606 193058 465648 193294
rect 465328 192896 465648 193058
rect 496048 193294 496368 193456
rect 496048 193058 496090 193294
rect 496326 193058 496368 193294
rect 496048 192896 496368 193058
rect 526768 193294 527088 193456
rect 526768 193058 526810 193294
rect 527046 193058 527088 193294
rect 526768 192896 527088 193058
rect 204208 183294 204528 183456
rect 204208 183058 204250 183294
rect 204486 183058 204528 183294
rect 204208 182896 204528 183058
rect 234928 183294 235248 183456
rect 234928 183058 234970 183294
rect 235206 183058 235248 183294
rect 234928 182896 235248 183058
rect 265648 183294 265968 183456
rect 265648 183058 265690 183294
rect 265926 183058 265968 183294
rect 265648 182896 265968 183058
rect 296368 183294 296688 183456
rect 296368 183058 296410 183294
rect 296646 183058 296688 183294
rect 296368 182896 296688 183058
rect 327088 183294 327408 183456
rect 327088 183058 327130 183294
rect 327366 183058 327408 183294
rect 327088 182896 327408 183058
rect 357808 183294 358128 183456
rect 357808 183058 357850 183294
rect 358086 183058 358128 183294
rect 357808 182896 358128 183058
rect 388528 183294 388848 183456
rect 388528 183058 388570 183294
rect 388806 183058 388848 183294
rect 388528 182896 388848 183058
rect 419248 183294 419568 183456
rect 419248 183058 419290 183294
rect 419526 183058 419568 183294
rect 419248 182896 419568 183058
rect 449968 183294 450288 183456
rect 449968 183058 450010 183294
rect 450246 183058 450288 183294
rect 449968 182896 450288 183058
rect 480688 183294 481008 183456
rect 480688 183058 480730 183294
rect 480966 183058 481008 183294
rect 480688 182896 481008 183058
rect 511408 183294 511728 183456
rect 511408 183058 511450 183294
rect 511686 183058 511728 183294
rect 511408 182896 511728 183058
rect 542128 183294 542448 183456
rect 542128 183058 542170 183294
rect 542406 183058 542448 183294
rect 542128 182896 542448 183058
rect 195514 176718 195546 176954
rect 195782 176718 195866 176954
rect 196102 176718 196134 176954
rect 195514 156954 196134 176718
rect 559234 180614 559854 200378
rect 559234 180378 559266 180614
rect 559502 180378 559586 180614
rect 559822 180378 559854 180614
rect 219568 173294 219888 173456
rect 219568 173058 219610 173294
rect 219846 173058 219888 173294
rect 219568 172896 219888 173058
rect 250288 173294 250608 173456
rect 250288 173058 250330 173294
rect 250566 173058 250608 173294
rect 250288 172896 250608 173058
rect 281008 173294 281328 173456
rect 281008 173058 281050 173294
rect 281286 173058 281328 173294
rect 281008 172896 281328 173058
rect 311728 173294 312048 173456
rect 311728 173058 311770 173294
rect 312006 173058 312048 173294
rect 311728 172896 312048 173058
rect 342448 173294 342768 173456
rect 342448 173058 342490 173294
rect 342726 173058 342768 173294
rect 342448 172896 342768 173058
rect 373168 173294 373488 173456
rect 373168 173058 373210 173294
rect 373446 173058 373488 173294
rect 373168 172896 373488 173058
rect 403888 173294 404208 173456
rect 403888 173058 403930 173294
rect 404166 173058 404208 173294
rect 403888 172896 404208 173058
rect 434608 173294 434928 173456
rect 434608 173058 434650 173294
rect 434886 173058 434928 173294
rect 434608 172896 434928 173058
rect 465328 173294 465648 173456
rect 465328 173058 465370 173294
rect 465606 173058 465648 173294
rect 465328 172896 465648 173058
rect 496048 173294 496368 173456
rect 496048 173058 496090 173294
rect 496326 173058 496368 173294
rect 496048 172896 496368 173058
rect 526768 173294 527088 173456
rect 526768 173058 526810 173294
rect 527046 173058 527088 173294
rect 526768 172896 527088 173058
rect 204208 163294 204528 163456
rect 204208 163058 204250 163294
rect 204486 163058 204528 163294
rect 204208 162896 204528 163058
rect 234928 163294 235248 163456
rect 234928 163058 234970 163294
rect 235206 163058 235248 163294
rect 234928 162896 235248 163058
rect 265648 163294 265968 163456
rect 265648 163058 265690 163294
rect 265926 163058 265968 163294
rect 265648 162896 265968 163058
rect 296368 163294 296688 163456
rect 296368 163058 296410 163294
rect 296646 163058 296688 163294
rect 296368 162896 296688 163058
rect 327088 163294 327408 163456
rect 327088 163058 327130 163294
rect 327366 163058 327408 163294
rect 327088 162896 327408 163058
rect 357808 163294 358128 163456
rect 357808 163058 357850 163294
rect 358086 163058 358128 163294
rect 357808 162896 358128 163058
rect 388528 163294 388848 163456
rect 388528 163058 388570 163294
rect 388806 163058 388848 163294
rect 388528 162896 388848 163058
rect 419248 163294 419568 163456
rect 419248 163058 419290 163294
rect 419526 163058 419568 163294
rect 419248 162896 419568 163058
rect 449968 163294 450288 163456
rect 449968 163058 450010 163294
rect 450246 163058 450288 163294
rect 449968 162896 450288 163058
rect 480688 163294 481008 163456
rect 480688 163058 480730 163294
rect 480966 163058 481008 163294
rect 480688 162896 481008 163058
rect 511408 163294 511728 163456
rect 511408 163058 511450 163294
rect 511686 163058 511728 163294
rect 511408 162896 511728 163058
rect 542128 163294 542448 163456
rect 542128 163058 542170 163294
rect 542406 163058 542448 163294
rect 542128 162896 542448 163058
rect 195514 156718 195546 156954
rect 195782 156718 195866 156954
rect 196102 156718 196134 156954
rect 195514 136954 196134 156718
rect 559234 160614 559854 180378
rect 559234 160378 559266 160614
rect 559502 160378 559586 160614
rect 559822 160378 559854 160614
rect 219568 153294 219888 153456
rect 219568 153058 219610 153294
rect 219846 153058 219888 153294
rect 219568 152896 219888 153058
rect 250288 153294 250608 153456
rect 250288 153058 250330 153294
rect 250566 153058 250608 153294
rect 250288 152896 250608 153058
rect 281008 153294 281328 153456
rect 281008 153058 281050 153294
rect 281286 153058 281328 153294
rect 281008 152896 281328 153058
rect 311728 153294 312048 153456
rect 311728 153058 311770 153294
rect 312006 153058 312048 153294
rect 311728 152896 312048 153058
rect 342448 153294 342768 153456
rect 342448 153058 342490 153294
rect 342726 153058 342768 153294
rect 342448 152896 342768 153058
rect 373168 153294 373488 153456
rect 373168 153058 373210 153294
rect 373446 153058 373488 153294
rect 373168 152896 373488 153058
rect 403888 153294 404208 153456
rect 403888 153058 403930 153294
rect 404166 153058 404208 153294
rect 403888 152896 404208 153058
rect 434608 153294 434928 153456
rect 434608 153058 434650 153294
rect 434886 153058 434928 153294
rect 434608 152896 434928 153058
rect 465328 153294 465648 153456
rect 465328 153058 465370 153294
rect 465606 153058 465648 153294
rect 465328 152896 465648 153058
rect 496048 153294 496368 153456
rect 496048 153058 496090 153294
rect 496326 153058 496368 153294
rect 496048 152896 496368 153058
rect 526768 153294 527088 153456
rect 526768 153058 526810 153294
rect 527046 153058 527088 153294
rect 526768 152896 527088 153058
rect 204208 143294 204528 143456
rect 204208 143058 204250 143294
rect 204486 143058 204528 143294
rect 204208 142896 204528 143058
rect 234928 143294 235248 143456
rect 234928 143058 234970 143294
rect 235206 143058 235248 143294
rect 234928 142896 235248 143058
rect 265648 143294 265968 143456
rect 265648 143058 265690 143294
rect 265926 143058 265968 143294
rect 265648 142896 265968 143058
rect 296368 143294 296688 143456
rect 296368 143058 296410 143294
rect 296646 143058 296688 143294
rect 296368 142896 296688 143058
rect 327088 143294 327408 143456
rect 327088 143058 327130 143294
rect 327366 143058 327408 143294
rect 327088 142896 327408 143058
rect 357808 143294 358128 143456
rect 357808 143058 357850 143294
rect 358086 143058 358128 143294
rect 357808 142896 358128 143058
rect 388528 143294 388848 143456
rect 388528 143058 388570 143294
rect 388806 143058 388848 143294
rect 388528 142896 388848 143058
rect 419248 143294 419568 143456
rect 419248 143058 419290 143294
rect 419526 143058 419568 143294
rect 419248 142896 419568 143058
rect 449968 143294 450288 143456
rect 449968 143058 450010 143294
rect 450246 143058 450288 143294
rect 449968 142896 450288 143058
rect 480688 143294 481008 143456
rect 480688 143058 480730 143294
rect 480966 143058 481008 143294
rect 480688 142896 481008 143058
rect 511408 143294 511728 143456
rect 511408 143058 511450 143294
rect 511686 143058 511728 143294
rect 511408 142896 511728 143058
rect 542128 143294 542448 143456
rect 542128 143058 542170 143294
rect 542406 143058 542448 143294
rect 542128 142896 542448 143058
rect 195514 136718 195546 136954
rect 195782 136718 195866 136954
rect 196102 136718 196134 136954
rect 195514 116954 196134 136718
rect 559234 140614 559854 160378
rect 559234 140378 559266 140614
rect 559502 140378 559586 140614
rect 559822 140378 559854 140614
rect 219568 133294 219888 133456
rect 219568 133058 219610 133294
rect 219846 133058 219888 133294
rect 219568 132896 219888 133058
rect 250288 133294 250608 133456
rect 250288 133058 250330 133294
rect 250566 133058 250608 133294
rect 250288 132896 250608 133058
rect 281008 133294 281328 133456
rect 281008 133058 281050 133294
rect 281286 133058 281328 133294
rect 281008 132896 281328 133058
rect 311728 133294 312048 133456
rect 311728 133058 311770 133294
rect 312006 133058 312048 133294
rect 311728 132896 312048 133058
rect 342448 133294 342768 133456
rect 342448 133058 342490 133294
rect 342726 133058 342768 133294
rect 342448 132896 342768 133058
rect 373168 133294 373488 133456
rect 373168 133058 373210 133294
rect 373446 133058 373488 133294
rect 373168 132896 373488 133058
rect 403888 133294 404208 133456
rect 403888 133058 403930 133294
rect 404166 133058 404208 133294
rect 403888 132896 404208 133058
rect 434608 133294 434928 133456
rect 434608 133058 434650 133294
rect 434886 133058 434928 133294
rect 434608 132896 434928 133058
rect 465328 133294 465648 133456
rect 465328 133058 465370 133294
rect 465606 133058 465648 133294
rect 465328 132896 465648 133058
rect 496048 133294 496368 133456
rect 496048 133058 496090 133294
rect 496326 133058 496368 133294
rect 496048 132896 496368 133058
rect 526768 133294 527088 133456
rect 526768 133058 526810 133294
rect 527046 133058 527088 133294
rect 526768 132896 527088 133058
rect 204208 123294 204528 123456
rect 204208 123058 204250 123294
rect 204486 123058 204528 123294
rect 204208 122896 204528 123058
rect 234928 123294 235248 123456
rect 234928 123058 234970 123294
rect 235206 123058 235248 123294
rect 234928 122896 235248 123058
rect 265648 123294 265968 123456
rect 265648 123058 265690 123294
rect 265926 123058 265968 123294
rect 265648 122896 265968 123058
rect 296368 123294 296688 123456
rect 296368 123058 296410 123294
rect 296646 123058 296688 123294
rect 296368 122896 296688 123058
rect 327088 123294 327408 123456
rect 327088 123058 327130 123294
rect 327366 123058 327408 123294
rect 327088 122896 327408 123058
rect 357808 123294 358128 123456
rect 357808 123058 357850 123294
rect 358086 123058 358128 123294
rect 357808 122896 358128 123058
rect 388528 123294 388848 123456
rect 388528 123058 388570 123294
rect 388806 123058 388848 123294
rect 388528 122896 388848 123058
rect 419248 123294 419568 123456
rect 419248 123058 419290 123294
rect 419526 123058 419568 123294
rect 419248 122896 419568 123058
rect 449968 123294 450288 123456
rect 449968 123058 450010 123294
rect 450246 123058 450288 123294
rect 449968 122896 450288 123058
rect 480688 123294 481008 123456
rect 480688 123058 480730 123294
rect 480966 123058 481008 123294
rect 480688 122896 481008 123058
rect 511408 123294 511728 123456
rect 511408 123058 511450 123294
rect 511686 123058 511728 123294
rect 511408 122896 511728 123058
rect 542128 123294 542448 123456
rect 542128 123058 542170 123294
rect 542406 123058 542448 123294
rect 542128 122896 542448 123058
rect 195514 116718 195546 116954
rect 195782 116718 195866 116954
rect 196102 116718 196134 116954
rect 195514 96954 196134 116718
rect 559234 120614 559854 140378
rect 559234 120378 559266 120614
rect 559502 120378 559586 120614
rect 559822 120378 559854 120614
rect 219568 113294 219888 113456
rect 219568 113058 219610 113294
rect 219846 113058 219888 113294
rect 219568 112896 219888 113058
rect 250288 113294 250608 113456
rect 250288 113058 250330 113294
rect 250566 113058 250608 113294
rect 250288 112896 250608 113058
rect 281008 113294 281328 113456
rect 281008 113058 281050 113294
rect 281286 113058 281328 113294
rect 281008 112896 281328 113058
rect 311728 113294 312048 113456
rect 311728 113058 311770 113294
rect 312006 113058 312048 113294
rect 311728 112896 312048 113058
rect 342448 113294 342768 113456
rect 342448 113058 342490 113294
rect 342726 113058 342768 113294
rect 342448 112896 342768 113058
rect 373168 113294 373488 113456
rect 373168 113058 373210 113294
rect 373446 113058 373488 113294
rect 373168 112896 373488 113058
rect 403888 113294 404208 113456
rect 403888 113058 403930 113294
rect 404166 113058 404208 113294
rect 403888 112896 404208 113058
rect 434608 113294 434928 113456
rect 434608 113058 434650 113294
rect 434886 113058 434928 113294
rect 434608 112896 434928 113058
rect 465328 113294 465648 113456
rect 465328 113058 465370 113294
rect 465606 113058 465648 113294
rect 465328 112896 465648 113058
rect 496048 113294 496368 113456
rect 496048 113058 496090 113294
rect 496326 113058 496368 113294
rect 496048 112896 496368 113058
rect 526768 113294 527088 113456
rect 526768 113058 526810 113294
rect 527046 113058 527088 113294
rect 526768 112896 527088 113058
rect 204208 103294 204528 103456
rect 204208 103058 204250 103294
rect 204486 103058 204528 103294
rect 204208 102896 204528 103058
rect 234928 103294 235248 103456
rect 234928 103058 234970 103294
rect 235206 103058 235248 103294
rect 234928 102896 235248 103058
rect 265648 103294 265968 103456
rect 265648 103058 265690 103294
rect 265926 103058 265968 103294
rect 265648 102896 265968 103058
rect 296368 103294 296688 103456
rect 296368 103058 296410 103294
rect 296646 103058 296688 103294
rect 296368 102896 296688 103058
rect 327088 103294 327408 103456
rect 327088 103058 327130 103294
rect 327366 103058 327408 103294
rect 327088 102896 327408 103058
rect 357808 103294 358128 103456
rect 357808 103058 357850 103294
rect 358086 103058 358128 103294
rect 357808 102896 358128 103058
rect 388528 103294 388848 103456
rect 388528 103058 388570 103294
rect 388806 103058 388848 103294
rect 388528 102896 388848 103058
rect 419248 103294 419568 103456
rect 419248 103058 419290 103294
rect 419526 103058 419568 103294
rect 419248 102896 419568 103058
rect 449968 103294 450288 103456
rect 449968 103058 450010 103294
rect 450246 103058 450288 103294
rect 449968 102896 450288 103058
rect 480688 103294 481008 103456
rect 480688 103058 480730 103294
rect 480966 103058 481008 103294
rect 480688 102896 481008 103058
rect 511408 103294 511728 103456
rect 511408 103058 511450 103294
rect 511686 103058 511728 103294
rect 511408 102896 511728 103058
rect 542128 103294 542448 103456
rect 542128 103058 542170 103294
rect 542406 103058 542448 103294
rect 542128 102896 542448 103058
rect 195514 96718 195546 96954
rect 195782 96718 195866 96954
rect 196102 96718 196134 96954
rect 195514 76954 196134 96718
rect 559234 100614 559854 120378
rect 559234 100378 559266 100614
rect 559502 100378 559586 100614
rect 559822 100378 559854 100614
rect 219568 93294 219888 93456
rect 219568 93058 219610 93294
rect 219846 93058 219888 93294
rect 219568 92896 219888 93058
rect 250288 93294 250608 93456
rect 250288 93058 250330 93294
rect 250566 93058 250608 93294
rect 250288 92896 250608 93058
rect 281008 93294 281328 93456
rect 281008 93058 281050 93294
rect 281286 93058 281328 93294
rect 281008 92896 281328 93058
rect 311728 93294 312048 93456
rect 311728 93058 311770 93294
rect 312006 93058 312048 93294
rect 311728 92896 312048 93058
rect 342448 93294 342768 93456
rect 342448 93058 342490 93294
rect 342726 93058 342768 93294
rect 342448 92896 342768 93058
rect 373168 93294 373488 93456
rect 373168 93058 373210 93294
rect 373446 93058 373488 93294
rect 373168 92896 373488 93058
rect 403888 93294 404208 93456
rect 403888 93058 403930 93294
rect 404166 93058 404208 93294
rect 403888 92896 404208 93058
rect 434608 93294 434928 93456
rect 434608 93058 434650 93294
rect 434886 93058 434928 93294
rect 434608 92896 434928 93058
rect 465328 93294 465648 93456
rect 465328 93058 465370 93294
rect 465606 93058 465648 93294
rect 465328 92896 465648 93058
rect 496048 93294 496368 93456
rect 496048 93058 496090 93294
rect 496326 93058 496368 93294
rect 496048 92896 496368 93058
rect 526768 93294 527088 93456
rect 526768 93058 526810 93294
rect 527046 93058 527088 93294
rect 526768 92896 527088 93058
rect 204208 83294 204528 83456
rect 204208 83058 204250 83294
rect 204486 83058 204528 83294
rect 204208 82896 204528 83058
rect 234928 83294 235248 83456
rect 234928 83058 234970 83294
rect 235206 83058 235248 83294
rect 234928 82896 235248 83058
rect 265648 83294 265968 83456
rect 265648 83058 265690 83294
rect 265926 83058 265968 83294
rect 265648 82896 265968 83058
rect 296368 83294 296688 83456
rect 296368 83058 296410 83294
rect 296646 83058 296688 83294
rect 296368 82896 296688 83058
rect 327088 83294 327408 83456
rect 327088 83058 327130 83294
rect 327366 83058 327408 83294
rect 327088 82896 327408 83058
rect 357808 83294 358128 83456
rect 357808 83058 357850 83294
rect 358086 83058 358128 83294
rect 357808 82896 358128 83058
rect 388528 83294 388848 83456
rect 388528 83058 388570 83294
rect 388806 83058 388848 83294
rect 388528 82896 388848 83058
rect 419248 83294 419568 83456
rect 419248 83058 419290 83294
rect 419526 83058 419568 83294
rect 419248 82896 419568 83058
rect 449968 83294 450288 83456
rect 449968 83058 450010 83294
rect 450246 83058 450288 83294
rect 449968 82896 450288 83058
rect 480688 83294 481008 83456
rect 480688 83058 480730 83294
rect 480966 83058 481008 83294
rect 480688 82896 481008 83058
rect 511408 83294 511728 83456
rect 511408 83058 511450 83294
rect 511686 83058 511728 83294
rect 511408 82896 511728 83058
rect 542128 83294 542448 83456
rect 542128 83058 542170 83294
rect 542406 83058 542448 83294
rect 542128 82896 542448 83058
rect 195514 76718 195546 76954
rect 195782 76718 195866 76954
rect 196102 76718 196134 76954
rect 195514 56954 196134 76718
rect 559234 80614 559854 100378
rect 559234 80378 559266 80614
rect 559502 80378 559586 80614
rect 559822 80378 559854 80614
rect 219568 73294 219888 73456
rect 219568 73058 219610 73294
rect 219846 73058 219888 73294
rect 219568 72896 219888 73058
rect 250288 73294 250608 73456
rect 250288 73058 250330 73294
rect 250566 73058 250608 73294
rect 250288 72896 250608 73058
rect 281008 73294 281328 73456
rect 281008 73058 281050 73294
rect 281286 73058 281328 73294
rect 281008 72896 281328 73058
rect 311728 73294 312048 73456
rect 311728 73058 311770 73294
rect 312006 73058 312048 73294
rect 311728 72896 312048 73058
rect 342448 73294 342768 73456
rect 342448 73058 342490 73294
rect 342726 73058 342768 73294
rect 342448 72896 342768 73058
rect 373168 73294 373488 73456
rect 373168 73058 373210 73294
rect 373446 73058 373488 73294
rect 373168 72896 373488 73058
rect 403888 73294 404208 73456
rect 403888 73058 403930 73294
rect 404166 73058 404208 73294
rect 403888 72896 404208 73058
rect 434608 73294 434928 73456
rect 434608 73058 434650 73294
rect 434886 73058 434928 73294
rect 434608 72896 434928 73058
rect 465328 73294 465648 73456
rect 465328 73058 465370 73294
rect 465606 73058 465648 73294
rect 465328 72896 465648 73058
rect 496048 73294 496368 73456
rect 496048 73058 496090 73294
rect 496326 73058 496368 73294
rect 496048 72896 496368 73058
rect 526768 73294 527088 73456
rect 526768 73058 526810 73294
rect 527046 73058 527088 73294
rect 526768 72896 527088 73058
rect 204208 63294 204528 63456
rect 204208 63058 204250 63294
rect 204486 63058 204528 63294
rect 204208 62896 204528 63058
rect 234928 63294 235248 63456
rect 234928 63058 234970 63294
rect 235206 63058 235248 63294
rect 234928 62896 235248 63058
rect 265648 63294 265968 63456
rect 265648 63058 265690 63294
rect 265926 63058 265968 63294
rect 265648 62896 265968 63058
rect 296368 63294 296688 63456
rect 296368 63058 296410 63294
rect 296646 63058 296688 63294
rect 296368 62896 296688 63058
rect 327088 63294 327408 63456
rect 327088 63058 327130 63294
rect 327366 63058 327408 63294
rect 327088 62896 327408 63058
rect 357808 63294 358128 63456
rect 357808 63058 357850 63294
rect 358086 63058 358128 63294
rect 357808 62896 358128 63058
rect 388528 63294 388848 63456
rect 388528 63058 388570 63294
rect 388806 63058 388848 63294
rect 388528 62896 388848 63058
rect 419248 63294 419568 63456
rect 419248 63058 419290 63294
rect 419526 63058 419568 63294
rect 419248 62896 419568 63058
rect 449968 63294 450288 63456
rect 449968 63058 450010 63294
rect 450246 63058 450288 63294
rect 449968 62896 450288 63058
rect 480688 63294 481008 63456
rect 480688 63058 480730 63294
rect 480966 63058 481008 63294
rect 480688 62896 481008 63058
rect 511408 63294 511728 63456
rect 511408 63058 511450 63294
rect 511686 63058 511728 63294
rect 511408 62896 511728 63058
rect 542128 63294 542448 63456
rect 542128 63058 542170 63294
rect 542406 63058 542448 63294
rect 542128 62896 542448 63058
rect 559234 60614 559854 80378
rect 559234 60378 559266 60614
rect 559502 60378 559586 60614
rect 559822 60378 559854 60614
rect 195514 56718 195546 56954
rect 195782 56718 195866 56954
rect 196102 56718 196134 56954
rect 195514 36954 196134 56718
rect 195514 36718 195546 36954
rect 195782 36718 195866 36954
rect 196102 36718 196134 36954
rect 195514 16954 196134 36718
rect 195514 16718 195546 16954
rect 195782 16718 195866 16954
rect 196102 16718 196134 16954
rect 195514 -3226 196134 16718
rect 195514 -3462 195546 -3226
rect 195782 -3462 195866 -3226
rect 196102 -3462 196134 -3226
rect 195514 -3546 196134 -3462
rect 195514 -3782 195546 -3546
rect 195782 -3782 195866 -3546
rect 196102 -3782 196134 -3546
rect 195514 -3814 196134 -3782
rect 199234 40614 199854 58000
rect 199234 40378 199266 40614
rect 199502 40378 199586 40614
rect 199822 40378 199854 40614
rect 199234 20614 199854 40378
rect 199234 20378 199266 20614
rect 199502 20378 199586 20614
rect 199822 20378 199854 20614
rect 199234 -5146 199854 20378
rect 201794 43294 202414 58000
rect 201794 43058 201826 43294
rect 202062 43058 202146 43294
rect 202382 43058 202414 43294
rect 201794 23294 202414 43058
rect 201794 23058 201826 23294
rect 202062 23058 202146 23294
rect 202382 23058 202414 23294
rect 201794 3294 202414 23058
rect 201794 3058 201826 3294
rect 202062 3058 202146 3294
rect 202382 3058 202414 3294
rect 201794 -346 202414 3058
rect 201794 -582 201826 -346
rect 202062 -582 202146 -346
rect 202382 -582 202414 -346
rect 201794 -666 202414 -582
rect 201794 -902 201826 -666
rect 202062 -902 202146 -666
rect 202382 -902 202414 -666
rect 201794 -1894 202414 -902
rect 202954 44274 203574 58000
rect 202954 44038 202986 44274
rect 203222 44038 203306 44274
rect 203542 44038 203574 44274
rect 202954 24274 203574 44038
rect 202954 24038 202986 24274
rect 203222 24038 203306 24274
rect 203542 24038 203574 24274
rect 199234 -5382 199266 -5146
rect 199502 -5382 199586 -5146
rect 199822 -5382 199854 -5146
rect 199234 -5466 199854 -5382
rect 199234 -5702 199266 -5466
rect 199502 -5702 199586 -5466
rect 199822 -5702 199854 -5466
rect 199234 -5734 199854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 202954 -7066 203574 24038
rect 205514 46954 206134 58000
rect 205514 46718 205546 46954
rect 205782 46718 205866 46954
rect 206102 46718 206134 46954
rect 205514 26954 206134 46718
rect 205514 26718 205546 26954
rect 205782 26718 205866 26954
rect 206102 26718 206134 26954
rect 205514 6954 206134 26718
rect 205514 6718 205546 6954
rect 205782 6718 205866 6954
rect 206102 6718 206134 6954
rect 205514 -2266 206134 6718
rect 205514 -2502 205546 -2266
rect 205782 -2502 205866 -2266
rect 206102 -2502 206134 -2266
rect 205514 -2586 206134 -2502
rect 205514 -2822 205546 -2586
rect 205782 -2822 205866 -2586
rect 206102 -2822 206134 -2586
rect 205514 -3814 206134 -2822
rect 209234 50614 209854 58000
rect 209234 50378 209266 50614
rect 209502 50378 209586 50614
rect 209822 50378 209854 50614
rect 209234 30614 209854 50378
rect 209234 30378 209266 30614
rect 209502 30378 209586 30614
rect 209822 30378 209854 30614
rect 209234 10614 209854 30378
rect 209234 10378 209266 10614
rect 209502 10378 209586 10614
rect 209822 10378 209854 10614
rect 209234 -4186 209854 10378
rect 211794 53294 212414 58000
rect 211794 53058 211826 53294
rect 212062 53058 212146 53294
rect 212382 53058 212414 53294
rect 211794 33294 212414 53058
rect 211794 33058 211826 33294
rect 212062 33058 212146 33294
rect 212382 33058 212414 33294
rect 211794 13294 212414 33058
rect 211794 13058 211826 13294
rect 212062 13058 212146 13294
rect 212382 13058 212414 13294
rect 211794 -1306 212414 13058
rect 211794 -1542 211826 -1306
rect 212062 -1542 212146 -1306
rect 212382 -1542 212414 -1306
rect 211794 -1626 212414 -1542
rect 211794 -1862 211826 -1626
rect 212062 -1862 212146 -1626
rect 212382 -1862 212414 -1626
rect 211794 -1894 212414 -1862
rect 212954 54274 213574 58000
rect 212954 54038 212986 54274
rect 213222 54038 213306 54274
rect 213542 54038 213574 54274
rect 212954 34274 213574 54038
rect 212954 34038 212986 34274
rect 213222 34038 213306 34274
rect 213542 34038 213574 34274
rect 212954 14274 213574 34038
rect 212954 14038 212986 14274
rect 213222 14038 213306 14274
rect 213542 14038 213574 14274
rect 209234 -4422 209266 -4186
rect 209502 -4422 209586 -4186
rect 209822 -4422 209854 -4186
rect 209234 -4506 209854 -4422
rect 209234 -4742 209266 -4506
rect 209502 -4742 209586 -4506
rect 209822 -4742 209854 -4506
rect 209234 -5734 209854 -4742
rect 202954 -7302 202986 -7066
rect 203222 -7302 203306 -7066
rect 203542 -7302 203574 -7066
rect 202954 -7386 203574 -7302
rect 202954 -7622 202986 -7386
rect 203222 -7622 203306 -7386
rect 203542 -7622 203574 -7386
rect 202954 -7654 203574 -7622
rect 212954 -6106 213574 14038
rect 215514 56954 216134 58000
rect 215514 56718 215546 56954
rect 215782 56718 215866 56954
rect 216102 56718 216134 56954
rect 215514 36954 216134 56718
rect 215514 36718 215546 36954
rect 215782 36718 215866 36954
rect 216102 36718 216134 36954
rect 215514 16954 216134 36718
rect 215514 16718 215546 16954
rect 215782 16718 215866 16954
rect 216102 16718 216134 16954
rect 215514 -3226 216134 16718
rect 215514 -3462 215546 -3226
rect 215782 -3462 215866 -3226
rect 216102 -3462 216134 -3226
rect 215514 -3546 216134 -3462
rect 215514 -3782 215546 -3546
rect 215782 -3782 215866 -3546
rect 216102 -3782 216134 -3546
rect 215514 -3814 216134 -3782
rect 219234 40614 219854 58000
rect 219234 40378 219266 40614
rect 219502 40378 219586 40614
rect 219822 40378 219854 40614
rect 219234 20614 219854 40378
rect 219234 20378 219266 20614
rect 219502 20378 219586 20614
rect 219822 20378 219854 20614
rect 219234 -5146 219854 20378
rect 221794 43294 222414 58000
rect 221794 43058 221826 43294
rect 222062 43058 222146 43294
rect 222382 43058 222414 43294
rect 221794 23294 222414 43058
rect 221794 23058 221826 23294
rect 222062 23058 222146 23294
rect 222382 23058 222414 23294
rect 221794 3294 222414 23058
rect 221794 3058 221826 3294
rect 222062 3058 222146 3294
rect 222382 3058 222414 3294
rect 221794 -346 222414 3058
rect 221794 -582 221826 -346
rect 222062 -582 222146 -346
rect 222382 -582 222414 -346
rect 221794 -666 222414 -582
rect 221794 -902 221826 -666
rect 222062 -902 222146 -666
rect 222382 -902 222414 -666
rect 221794 -1894 222414 -902
rect 222954 44274 223574 58000
rect 222954 44038 222986 44274
rect 223222 44038 223306 44274
rect 223542 44038 223574 44274
rect 222954 24274 223574 44038
rect 222954 24038 222986 24274
rect 223222 24038 223306 24274
rect 223542 24038 223574 24274
rect 219234 -5382 219266 -5146
rect 219502 -5382 219586 -5146
rect 219822 -5382 219854 -5146
rect 219234 -5466 219854 -5382
rect 219234 -5702 219266 -5466
rect 219502 -5702 219586 -5466
rect 219822 -5702 219854 -5466
rect 219234 -5734 219854 -5702
rect 212954 -6342 212986 -6106
rect 213222 -6342 213306 -6106
rect 213542 -6342 213574 -6106
rect 212954 -6426 213574 -6342
rect 212954 -6662 212986 -6426
rect 213222 -6662 213306 -6426
rect 213542 -6662 213574 -6426
rect 212954 -7654 213574 -6662
rect 222954 -7066 223574 24038
rect 225514 46954 226134 58000
rect 225514 46718 225546 46954
rect 225782 46718 225866 46954
rect 226102 46718 226134 46954
rect 225514 26954 226134 46718
rect 225514 26718 225546 26954
rect 225782 26718 225866 26954
rect 226102 26718 226134 26954
rect 225514 6954 226134 26718
rect 225514 6718 225546 6954
rect 225782 6718 225866 6954
rect 226102 6718 226134 6954
rect 225514 -2266 226134 6718
rect 225514 -2502 225546 -2266
rect 225782 -2502 225866 -2266
rect 226102 -2502 226134 -2266
rect 225514 -2586 226134 -2502
rect 225514 -2822 225546 -2586
rect 225782 -2822 225866 -2586
rect 226102 -2822 226134 -2586
rect 225514 -3814 226134 -2822
rect 229234 50614 229854 58000
rect 229234 50378 229266 50614
rect 229502 50378 229586 50614
rect 229822 50378 229854 50614
rect 229234 30614 229854 50378
rect 229234 30378 229266 30614
rect 229502 30378 229586 30614
rect 229822 30378 229854 30614
rect 229234 10614 229854 30378
rect 229234 10378 229266 10614
rect 229502 10378 229586 10614
rect 229822 10378 229854 10614
rect 229234 -4186 229854 10378
rect 231794 53294 232414 58000
rect 231794 53058 231826 53294
rect 232062 53058 232146 53294
rect 232382 53058 232414 53294
rect 231794 33294 232414 53058
rect 231794 33058 231826 33294
rect 232062 33058 232146 33294
rect 232382 33058 232414 33294
rect 231794 13294 232414 33058
rect 231794 13058 231826 13294
rect 232062 13058 232146 13294
rect 232382 13058 232414 13294
rect 231794 -1306 232414 13058
rect 231794 -1542 231826 -1306
rect 232062 -1542 232146 -1306
rect 232382 -1542 232414 -1306
rect 231794 -1626 232414 -1542
rect 231794 -1862 231826 -1626
rect 232062 -1862 232146 -1626
rect 232382 -1862 232414 -1626
rect 231794 -1894 232414 -1862
rect 232954 54274 233574 58000
rect 232954 54038 232986 54274
rect 233222 54038 233306 54274
rect 233542 54038 233574 54274
rect 232954 34274 233574 54038
rect 232954 34038 232986 34274
rect 233222 34038 233306 34274
rect 233542 34038 233574 34274
rect 232954 14274 233574 34038
rect 232954 14038 232986 14274
rect 233222 14038 233306 14274
rect 233542 14038 233574 14274
rect 229234 -4422 229266 -4186
rect 229502 -4422 229586 -4186
rect 229822 -4422 229854 -4186
rect 229234 -4506 229854 -4422
rect 229234 -4742 229266 -4506
rect 229502 -4742 229586 -4506
rect 229822 -4742 229854 -4506
rect 229234 -5734 229854 -4742
rect 222954 -7302 222986 -7066
rect 223222 -7302 223306 -7066
rect 223542 -7302 223574 -7066
rect 222954 -7386 223574 -7302
rect 222954 -7622 222986 -7386
rect 223222 -7622 223306 -7386
rect 223542 -7622 223574 -7386
rect 222954 -7654 223574 -7622
rect 232954 -6106 233574 14038
rect 235514 56954 236134 58000
rect 235514 56718 235546 56954
rect 235782 56718 235866 56954
rect 236102 56718 236134 56954
rect 235514 36954 236134 56718
rect 235514 36718 235546 36954
rect 235782 36718 235866 36954
rect 236102 36718 236134 36954
rect 235514 16954 236134 36718
rect 235514 16718 235546 16954
rect 235782 16718 235866 16954
rect 236102 16718 236134 16954
rect 235514 -3226 236134 16718
rect 235514 -3462 235546 -3226
rect 235782 -3462 235866 -3226
rect 236102 -3462 236134 -3226
rect 235514 -3546 236134 -3462
rect 235514 -3782 235546 -3546
rect 235782 -3782 235866 -3546
rect 236102 -3782 236134 -3546
rect 235514 -3814 236134 -3782
rect 239234 40614 239854 58000
rect 239234 40378 239266 40614
rect 239502 40378 239586 40614
rect 239822 40378 239854 40614
rect 239234 20614 239854 40378
rect 239234 20378 239266 20614
rect 239502 20378 239586 20614
rect 239822 20378 239854 20614
rect 239234 -5146 239854 20378
rect 241794 43294 242414 58000
rect 241794 43058 241826 43294
rect 242062 43058 242146 43294
rect 242382 43058 242414 43294
rect 241794 23294 242414 43058
rect 241794 23058 241826 23294
rect 242062 23058 242146 23294
rect 242382 23058 242414 23294
rect 241794 3294 242414 23058
rect 241794 3058 241826 3294
rect 242062 3058 242146 3294
rect 242382 3058 242414 3294
rect 241794 -346 242414 3058
rect 241794 -582 241826 -346
rect 242062 -582 242146 -346
rect 242382 -582 242414 -346
rect 241794 -666 242414 -582
rect 241794 -902 241826 -666
rect 242062 -902 242146 -666
rect 242382 -902 242414 -666
rect 241794 -1894 242414 -902
rect 242954 44274 243574 58000
rect 242954 44038 242986 44274
rect 243222 44038 243306 44274
rect 243542 44038 243574 44274
rect 242954 24274 243574 44038
rect 242954 24038 242986 24274
rect 243222 24038 243306 24274
rect 243542 24038 243574 24274
rect 239234 -5382 239266 -5146
rect 239502 -5382 239586 -5146
rect 239822 -5382 239854 -5146
rect 239234 -5466 239854 -5382
rect 239234 -5702 239266 -5466
rect 239502 -5702 239586 -5466
rect 239822 -5702 239854 -5466
rect 239234 -5734 239854 -5702
rect 232954 -6342 232986 -6106
rect 233222 -6342 233306 -6106
rect 233542 -6342 233574 -6106
rect 232954 -6426 233574 -6342
rect 232954 -6662 232986 -6426
rect 233222 -6662 233306 -6426
rect 233542 -6662 233574 -6426
rect 232954 -7654 233574 -6662
rect 242954 -7066 243574 24038
rect 245514 46954 246134 58000
rect 245514 46718 245546 46954
rect 245782 46718 245866 46954
rect 246102 46718 246134 46954
rect 245514 26954 246134 46718
rect 245514 26718 245546 26954
rect 245782 26718 245866 26954
rect 246102 26718 246134 26954
rect 245514 6954 246134 26718
rect 245514 6718 245546 6954
rect 245782 6718 245866 6954
rect 246102 6718 246134 6954
rect 245514 -2266 246134 6718
rect 245514 -2502 245546 -2266
rect 245782 -2502 245866 -2266
rect 246102 -2502 246134 -2266
rect 245514 -2586 246134 -2502
rect 245514 -2822 245546 -2586
rect 245782 -2822 245866 -2586
rect 246102 -2822 246134 -2586
rect 245514 -3814 246134 -2822
rect 249234 50614 249854 58000
rect 249234 50378 249266 50614
rect 249502 50378 249586 50614
rect 249822 50378 249854 50614
rect 249234 30614 249854 50378
rect 249234 30378 249266 30614
rect 249502 30378 249586 30614
rect 249822 30378 249854 30614
rect 249234 10614 249854 30378
rect 249234 10378 249266 10614
rect 249502 10378 249586 10614
rect 249822 10378 249854 10614
rect 249234 -4186 249854 10378
rect 251794 53294 252414 58000
rect 251794 53058 251826 53294
rect 252062 53058 252146 53294
rect 252382 53058 252414 53294
rect 251794 33294 252414 53058
rect 251794 33058 251826 33294
rect 252062 33058 252146 33294
rect 252382 33058 252414 33294
rect 251794 13294 252414 33058
rect 251794 13058 251826 13294
rect 252062 13058 252146 13294
rect 252382 13058 252414 13294
rect 251794 -1306 252414 13058
rect 251794 -1542 251826 -1306
rect 252062 -1542 252146 -1306
rect 252382 -1542 252414 -1306
rect 251794 -1626 252414 -1542
rect 251794 -1862 251826 -1626
rect 252062 -1862 252146 -1626
rect 252382 -1862 252414 -1626
rect 251794 -1894 252414 -1862
rect 252954 54274 253574 58000
rect 252954 54038 252986 54274
rect 253222 54038 253306 54274
rect 253542 54038 253574 54274
rect 252954 34274 253574 54038
rect 252954 34038 252986 34274
rect 253222 34038 253306 34274
rect 253542 34038 253574 34274
rect 252954 14274 253574 34038
rect 252954 14038 252986 14274
rect 253222 14038 253306 14274
rect 253542 14038 253574 14274
rect 249234 -4422 249266 -4186
rect 249502 -4422 249586 -4186
rect 249822 -4422 249854 -4186
rect 249234 -4506 249854 -4422
rect 249234 -4742 249266 -4506
rect 249502 -4742 249586 -4506
rect 249822 -4742 249854 -4506
rect 249234 -5734 249854 -4742
rect 242954 -7302 242986 -7066
rect 243222 -7302 243306 -7066
rect 243542 -7302 243574 -7066
rect 242954 -7386 243574 -7302
rect 242954 -7622 242986 -7386
rect 243222 -7622 243306 -7386
rect 243542 -7622 243574 -7386
rect 242954 -7654 243574 -7622
rect 252954 -6106 253574 14038
rect 255514 56954 256134 58000
rect 255514 56718 255546 56954
rect 255782 56718 255866 56954
rect 256102 56718 256134 56954
rect 255514 36954 256134 56718
rect 255514 36718 255546 36954
rect 255782 36718 255866 36954
rect 256102 36718 256134 36954
rect 255514 16954 256134 36718
rect 255514 16718 255546 16954
rect 255782 16718 255866 16954
rect 256102 16718 256134 16954
rect 255514 -3226 256134 16718
rect 255514 -3462 255546 -3226
rect 255782 -3462 255866 -3226
rect 256102 -3462 256134 -3226
rect 255514 -3546 256134 -3462
rect 255514 -3782 255546 -3546
rect 255782 -3782 255866 -3546
rect 256102 -3782 256134 -3546
rect 255514 -3814 256134 -3782
rect 259234 40614 259854 58000
rect 259234 40378 259266 40614
rect 259502 40378 259586 40614
rect 259822 40378 259854 40614
rect 259234 20614 259854 40378
rect 259234 20378 259266 20614
rect 259502 20378 259586 20614
rect 259822 20378 259854 20614
rect 259234 -5146 259854 20378
rect 261794 43294 262414 58000
rect 261794 43058 261826 43294
rect 262062 43058 262146 43294
rect 262382 43058 262414 43294
rect 261794 23294 262414 43058
rect 261794 23058 261826 23294
rect 262062 23058 262146 23294
rect 262382 23058 262414 23294
rect 261794 3294 262414 23058
rect 261794 3058 261826 3294
rect 262062 3058 262146 3294
rect 262382 3058 262414 3294
rect 261794 -346 262414 3058
rect 261794 -582 261826 -346
rect 262062 -582 262146 -346
rect 262382 -582 262414 -346
rect 261794 -666 262414 -582
rect 261794 -902 261826 -666
rect 262062 -902 262146 -666
rect 262382 -902 262414 -666
rect 261794 -1894 262414 -902
rect 262954 44274 263574 58000
rect 262954 44038 262986 44274
rect 263222 44038 263306 44274
rect 263542 44038 263574 44274
rect 262954 24274 263574 44038
rect 262954 24038 262986 24274
rect 263222 24038 263306 24274
rect 263542 24038 263574 24274
rect 259234 -5382 259266 -5146
rect 259502 -5382 259586 -5146
rect 259822 -5382 259854 -5146
rect 259234 -5466 259854 -5382
rect 259234 -5702 259266 -5466
rect 259502 -5702 259586 -5466
rect 259822 -5702 259854 -5466
rect 259234 -5734 259854 -5702
rect 252954 -6342 252986 -6106
rect 253222 -6342 253306 -6106
rect 253542 -6342 253574 -6106
rect 252954 -6426 253574 -6342
rect 252954 -6662 252986 -6426
rect 253222 -6662 253306 -6426
rect 253542 -6662 253574 -6426
rect 252954 -7654 253574 -6662
rect 262954 -7066 263574 24038
rect 265514 46954 266134 58000
rect 265514 46718 265546 46954
rect 265782 46718 265866 46954
rect 266102 46718 266134 46954
rect 265514 26954 266134 46718
rect 265514 26718 265546 26954
rect 265782 26718 265866 26954
rect 266102 26718 266134 26954
rect 265514 6954 266134 26718
rect 265514 6718 265546 6954
rect 265782 6718 265866 6954
rect 266102 6718 266134 6954
rect 265514 -2266 266134 6718
rect 265514 -2502 265546 -2266
rect 265782 -2502 265866 -2266
rect 266102 -2502 266134 -2266
rect 265514 -2586 266134 -2502
rect 265514 -2822 265546 -2586
rect 265782 -2822 265866 -2586
rect 266102 -2822 266134 -2586
rect 265514 -3814 266134 -2822
rect 269234 50614 269854 58000
rect 269234 50378 269266 50614
rect 269502 50378 269586 50614
rect 269822 50378 269854 50614
rect 269234 30614 269854 50378
rect 269234 30378 269266 30614
rect 269502 30378 269586 30614
rect 269822 30378 269854 30614
rect 269234 10614 269854 30378
rect 269234 10378 269266 10614
rect 269502 10378 269586 10614
rect 269822 10378 269854 10614
rect 269234 -4186 269854 10378
rect 271794 53294 272414 58000
rect 271794 53058 271826 53294
rect 272062 53058 272146 53294
rect 272382 53058 272414 53294
rect 271794 33294 272414 53058
rect 271794 33058 271826 33294
rect 272062 33058 272146 33294
rect 272382 33058 272414 33294
rect 271794 13294 272414 33058
rect 271794 13058 271826 13294
rect 272062 13058 272146 13294
rect 272382 13058 272414 13294
rect 271794 -1306 272414 13058
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 272954 54274 273574 58000
rect 272954 54038 272986 54274
rect 273222 54038 273306 54274
rect 273542 54038 273574 54274
rect 272954 34274 273574 54038
rect 272954 34038 272986 34274
rect 273222 34038 273306 34274
rect 273542 34038 273574 34274
rect 272954 14274 273574 34038
rect 272954 14038 272986 14274
rect 273222 14038 273306 14274
rect 273542 14038 273574 14274
rect 269234 -4422 269266 -4186
rect 269502 -4422 269586 -4186
rect 269822 -4422 269854 -4186
rect 269234 -4506 269854 -4422
rect 269234 -4742 269266 -4506
rect 269502 -4742 269586 -4506
rect 269822 -4742 269854 -4506
rect 269234 -5734 269854 -4742
rect 262954 -7302 262986 -7066
rect 263222 -7302 263306 -7066
rect 263542 -7302 263574 -7066
rect 262954 -7386 263574 -7302
rect 262954 -7622 262986 -7386
rect 263222 -7622 263306 -7386
rect 263542 -7622 263574 -7386
rect 262954 -7654 263574 -7622
rect 272954 -6106 273574 14038
rect 275514 56954 276134 58000
rect 275514 56718 275546 56954
rect 275782 56718 275866 56954
rect 276102 56718 276134 56954
rect 275514 36954 276134 56718
rect 275514 36718 275546 36954
rect 275782 36718 275866 36954
rect 276102 36718 276134 36954
rect 275514 16954 276134 36718
rect 275514 16718 275546 16954
rect 275782 16718 275866 16954
rect 276102 16718 276134 16954
rect 275514 -3226 276134 16718
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 40614 279854 58000
rect 279234 40378 279266 40614
rect 279502 40378 279586 40614
rect 279822 40378 279854 40614
rect 279234 20614 279854 40378
rect 279234 20378 279266 20614
rect 279502 20378 279586 20614
rect 279822 20378 279854 20614
rect 279234 -5146 279854 20378
rect 281794 43294 282414 58000
rect 281794 43058 281826 43294
rect 282062 43058 282146 43294
rect 282382 43058 282414 43294
rect 281794 23294 282414 43058
rect 281794 23058 281826 23294
rect 282062 23058 282146 23294
rect 282382 23058 282414 23294
rect 281794 3294 282414 23058
rect 281794 3058 281826 3294
rect 282062 3058 282146 3294
rect 282382 3058 282414 3294
rect 281794 -346 282414 3058
rect 281794 -582 281826 -346
rect 282062 -582 282146 -346
rect 282382 -582 282414 -346
rect 281794 -666 282414 -582
rect 281794 -902 281826 -666
rect 282062 -902 282146 -666
rect 282382 -902 282414 -666
rect 281794 -1894 282414 -902
rect 282954 44274 283574 58000
rect 282954 44038 282986 44274
rect 283222 44038 283306 44274
rect 283542 44038 283574 44274
rect 282954 24274 283574 44038
rect 282954 24038 282986 24274
rect 283222 24038 283306 24274
rect 283542 24038 283574 24274
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 272954 -6342 272986 -6106
rect 273222 -6342 273306 -6106
rect 273542 -6342 273574 -6106
rect 272954 -6426 273574 -6342
rect 272954 -6662 272986 -6426
rect 273222 -6662 273306 -6426
rect 273542 -6662 273574 -6426
rect 272954 -7654 273574 -6662
rect 282954 -7066 283574 24038
rect 285514 46954 286134 58000
rect 285514 46718 285546 46954
rect 285782 46718 285866 46954
rect 286102 46718 286134 46954
rect 285514 26954 286134 46718
rect 285514 26718 285546 26954
rect 285782 26718 285866 26954
rect 286102 26718 286134 26954
rect 285514 6954 286134 26718
rect 285514 6718 285546 6954
rect 285782 6718 285866 6954
rect 286102 6718 286134 6954
rect 285514 -2266 286134 6718
rect 285514 -2502 285546 -2266
rect 285782 -2502 285866 -2266
rect 286102 -2502 286134 -2266
rect 285514 -2586 286134 -2502
rect 285514 -2822 285546 -2586
rect 285782 -2822 285866 -2586
rect 286102 -2822 286134 -2586
rect 285514 -3814 286134 -2822
rect 289234 50614 289854 58000
rect 289234 50378 289266 50614
rect 289502 50378 289586 50614
rect 289822 50378 289854 50614
rect 289234 30614 289854 50378
rect 289234 30378 289266 30614
rect 289502 30378 289586 30614
rect 289822 30378 289854 30614
rect 289234 10614 289854 30378
rect 289234 10378 289266 10614
rect 289502 10378 289586 10614
rect 289822 10378 289854 10614
rect 289234 -4186 289854 10378
rect 291794 53294 292414 58000
rect 291794 53058 291826 53294
rect 292062 53058 292146 53294
rect 292382 53058 292414 53294
rect 291794 33294 292414 53058
rect 291794 33058 291826 33294
rect 292062 33058 292146 33294
rect 292382 33058 292414 33294
rect 291794 13294 292414 33058
rect 291794 13058 291826 13294
rect 292062 13058 292146 13294
rect 292382 13058 292414 13294
rect 291794 -1306 292414 13058
rect 291794 -1542 291826 -1306
rect 292062 -1542 292146 -1306
rect 292382 -1542 292414 -1306
rect 291794 -1626 292414 -1542
rect 291794 -1862 291826 -1626
rect 292062 -1862 292146 -1626
rect 292382 -1862 292414 -1626
rect 291794 -1894 292414 -1862
rect 292954 54274 293574 58000
rect 292954 54038 292986 54274
rect 293222 54038 293306 54274
rect 293542 54038 293574 54274
rect 292954 34274 293574 54038
rect 292954 34038 292986 34274
rect 293222 34038 293306 34274
rect 293542 34038 293574 34274
rect 292954 14274 293574 34038
rect 292954 14038 292986 14274
rect 293222 14038 293306 14274
rect 293542 14038 293574 14274
rect 289234 -4422 289266 -4186
rect 289502 -4422 289586 -4186
rect 289822 -4422 289854 -4186
rect 289234 -4506 289854 -4422
rect 289234 -4742 289266 -4506
rect 289502 -4742 289586 -4506
rect 289822 -4742 289854 -4506
rect 289234 -5734 289854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 292954 -6106 293574 14038
rect 295514 56954 296134 58000
rect 295514 56718 295546 56954
rect 295782 56718 295866 56954
rect 296102 56718 296134 56954
rect 295514 36954 296134 56718
rect 295514 36718 295546 36954
rect 295782 36718 295866 36954
rect 296102 36718 296134 36954
rect 295514 16954 296134 36718
rect 295514 16718 295546 16954
rect 295782 16718 295866 16954
rect 296102 16718 296134 16954
rect 295514 -3226 296134 16718
rect 295514 -3462 295546 -3226
rect 295782 -3462 295866 -3226
rect 296102 -3462 296134 -3226
rect 295514 -3546 296134 -3462
rect 295514 -3782 295546 -3546
rect 295782 -3782 295866 -3546
rect 296102 -3782 296134 -3546
rect 295514 -3814 296134 -3782
rect 299234 40614 299854 58000
rect 299234 40378 299266 40614
rect 299502 40378 299586 40614
rect 299822 40378 299854 40614
rect 299234 20614 299854 40378
rect 299234 20378 299266 20614
rect 299502 20378 299586 20614
rect 299822 20378 299854 20614
rect 299234 -5146 299854 20378
rect 301794 43294 302414 58000
rect 301794 43058 301826 43294
rect 302062 43058 302146 43294
rect 302382 43058 302414 43294
rect 301794 23294 302414 43058
rect 301794 23058 301826 23294
rect 302062 23058 302146 23294
rect 302382 23058 302414 23294
rect 301794 3294 302414 23058
rect 301794 3058 301826 3294
rect 302062 3058 302146 3294
rect 302382 3058 302414 3294
rect 301794 -346 302414 3058
rect 301794 -582 301826 -346
rect 302062 -582 302146 -346
rect 302382 -582 302414 -346
rect 301794 -666 302414 -582
rect 301794 -902 301826 -666
rect 302062 -902 302146 -666
rect 302382 -902 302414 -666
rect 301794 -1894 302414 -902
rect 302954 44274 303574 58000
rect 302954 44038 302986 44274
rect 303222 44038 303306 44274
rect 303542 44038 303574 44274
rect 302954 24274 303574 44038
rect 302954 24038 302986 24274
rect 303222 24038 303306 24274
rect 303542 24038 303574 24274
rect 299234 -5382 299266 -5146
rect 299502 -5382 299586 -5146
rect 299822 -5382 299854 -5146
rect 299234 -5466 299854 -5382
rect 299234 -5702 299266 -5466
rect 299502 -5702 299586 -5466
rect 299822 -5702 299854 -5466
rect 299234 -5734 299854 -5702
rect 292954 -6342 292986 -6106
rect 293222 -6342 293306 -6106
rect 293542 -6342 293574 -6106
rect 292954 -6426 293574 -6342
rect 292954 -6662 292986 -6426
rect 293222 -6662 293306 -6426
rect 293542 -6662 293574 -6426
rect 292954 -7654 293574 -6662
rect 302954 -7066 303574 24038
rect 305514 46954 306134 58000
rect 305514 46718 305546 46954
rect 305782 46718 305866 46954
rect 306102 46718 306134 46954
rect 305514 26954 306134 46718
rect 305514 26718 305546 26954
rect 305782 26718 305866 26954
rect 306102 26718 306134 26954
rect 305514 6954 306134 26718
rect 305514 6718 305546 6954
rect 305782 6718 305866 6954
rect 306102 6718 306134 6954
rect 305514 -2266 306134 6718
rect 305514 -2502 305546 -2266
rect 305782 -2502 305866 -2266
rect 306102 -2502 306134 -2266
rect 305514 -2586 306134 -2502
rect 305514 -2822 305546 -2586
rect 305782 -2822 305866 -2586
rect 306102 -2822 306134 -2586
rect 305514 -3814 306134 -2822
rect 309234 50614 309854 58000
rect 309234 50378 309266 50614
rect 309502 50378 309586 50614
rect 309822 50378 309854 50614
rect 309234 30614 309854 50378
rect 309234 30378 309266 30614
rect 309502 30378 309586 30614
rect 309822 30378 309854 30614
rect 309234 10614 309854 30378
rect 309234 10378 309266 10614
rect 309502 10378 309586 10614
rect 309822 10378 309854 10614
rect 309234 -4186 309854 10378
rect 311794 53294 312414 58000
rect 311794 53058 311826 53294
rect 312062 53058 312146 53294
rect 312382 53058 312414 53294
rect 311794 33294 312414 53058
rect 311794 33058 311826 33294
rect 312062 33058 312146 33294
rect 312382 33058 312414 33294
rect 311794 13294 312414 33058
rect 311794 13058 311826 13294
rect 312062 13058 312146 13294
rect 312382 13058 312414 13294
rect 311794 -1306 312414 13058
rect 311794 -1542 311826 -1306
rect 312062 -1542 312146 -1306
rect 312382 -1542 312414 -1306
rect 311794 -1626 312414 -1542
rect 311794 -1862 311826 -1626
rect 312062 -1862 312146 -1626
rect 312382 -1862 312414 -1626
rect 311794 -1894 312414 -1862
rect 312954 54274 313574 58000
rect 312954 54038 312986 54274
rect 313222 54038 313306 54274
rect 313542 54038 313574 54274
rect 312954 34274 313574 54038
rect 312954 34038 312986 34274
rect 313222 34038 313306 34274
rect 313542 34038 313574 34274
rect 312954 14274 313574 34038
rect 312954 14038 312986 14274
rect 313222 14038 313306 14274
rect 313542 14038 313574 14274
rect 309234 -4422 309266 -4186
rect 309502 -4422 309586 -4186
rect 309822 -4422 309854 -4186
rect 309234 -4506 309854 -4422
rect 309234 -4742 309266 -4506
rect 309502 -4742 309586 -4506
rect 309822 -4742 309854 -4506
rect 309234 -5734 309854 -4742
rect 302954 -7302 302986 -7066
rect 303222 -7302 303306 -7066
rect 303542 -7302 303574 -7066
rect 302954 -7386 303574 -7302
rect 302954 -7622 302986 -7386
rect 303222 -7622 303306 -7386
rect 303542 -7622 303574 -7386
rect 302954 -7654 303574 -7622
rect 312954 -6106 313574 14038
rect 315514 56954 316134 58000
rect 315514 56718 315546 56954
rect 315782 56718 315866 56954
rect 316102 56718 316134 56954
rect 315514 36954 316134 56718
rect 315514 36718 315546 36954
rect 315782 36718 315866 36954
rect 316102 36718 316134 36954
rect 315514 16954 316134 36718
rect 315514 16718 315546 16954
rect 315782 16718 315866 16954
rect 316102 16718 316134 16954
rect 315514 -3226 316134 16718
rect 315514 -3462 315546 -3226
rect 315782 -3462 315866 -3226
rect 316102 -3462 316134 -3226
rect 315514 -3546 316134 -3462
rect 315514 -3782 315546 -3546
rect 315782 -3782 315866 -3546
rect 316102 -3782 316134 -3546
rect 315514 -3814 316134 -3782
rect 319234 40614 319854 58000
rect 319234 40378 319266 40614
rect 319502 40378 319586 40614
rect 319822 40378 319854 40614
rect 319234 20614 319854 40378
rect 319234 20378 319266 20614
rect 319502 20378 319586 20614
rect 319822 20378 319854 20614
rect 319234 -5146 319854 20378
rect 321794 43294 322414 58000
rect 321794 43058 321826 43294
rect 322062 43058 322146 43294
rect 322382 43058 322414 43294
rect 321794 23294 322414 43058
rect 321794 23058 321826 23294
rect 322062 23058 322146 23294
rect 322382 23058 322414 23294
rect 321794 3294 322414 23058
rect 321794 3058 321826 3294
rect 322062 3058 322146 3294
rect 322382 3058 322414 3294
rect 321794 -346 322414 3058
rect 321794 -582 321826 -346
rect 322062 -582 322146 -346
rect 322382 -582 322414 -346
rect 321794 -666 322414 -582
rect 321794 -902 321826 -666
rect 322062 -902 322146 -666
rect 322382 -902 322414 -666
rect 321794 -1894 322414 -902
rect 322954 44274 323574 58000
rect 322954 44038 322986 44274
rect 323222 44038 323306 44274
rect 323542 44038 323574 44274
rect 322954 24274 323574 44038
rect 322954 24038 322986 24274
rect 323222 24038 323306 24274
rect 323542 24038 323574 24274
rect 319234 -5382 319266 -5146
rect 319502 -5382 319586 -5146
rect 319822 -5382 319854 -5146
rect 319234 -5466 319854 -5382
rect 319234 -5702 319266 -5466
rect 319502 -5702 319586 -5466
rect 319822 -5702 319854 -5466
rect 319234 -5734 319854 -5702
rect 312954 -6342 312986 -6106
rect 313222 -6342 313306 -6106
rect 313542 -6342 313574 -6106
rect 312954 -6426 313574 -6342
rect 312954 -6662 312986 -6426
rect 313222 -6662 313306 -6426
rect 313542 -6662 313574 -6426
rect 312954 -7654 313574 -6662
rect 322954 -7066 323574 24038
rect 325514 46954 326134 58000
rect 325514 46718 325546 46954
rect 325782 46718 325866 46954
rect 326102 46718 326134 46954
rect 325514 26954 326134 46718
rect 325514 26718 325546 26954
rect 325782 26718 325866 26954
rect 326102 26718 326134 26954
rect 325514 6954 326134 26718
rect 325514 6718 325546 6954
rect 325782 6718 325866 6954
rect 326102 6718 326134 6954
rect 325514 -2266 326134 6718
rect 325514 -2502 325546 -2266
rect 325782 -2502 325866 -2266
rect 326102 -2502 326134 -2266
rect 325514 -2586 326134 -2502
rect 325514 -2822 325546 -2586
rect 325782 -2822 325866 -2586
rect 326102 -2822 326134 -2586
rect 325514 -3814 326134 -2822
rect 329234 50614 329854 58000
rect 329234 50378 329266 50614
rect 329502 50378 329586 50614
rect 329822 50378 329854 50614
rect 329234 30614 329854 50378
rect 329234 30378 329266 30614
rect 329502 30378 329586 30614
rect 329822 30378 329854 30614
rect 329234 10614 329854 30378
rect 329234 10378 329266 10614
rect 329502 10378 329586 10614
rect 329822 10378 329854 10614
rect 329234 -4186 329854 10378
rect 331794 53294 332414 58000
rect 331794 53058 331826 53294
rect 332062 53058 332146 53294
rect 332382 53058 332414 53294
rect 331794 33294 332414 53058
rect 331794 33058 331826 33294
rect 332062 33058 332146 33294
rect 332382 33058 332414 33294
rect 331794 13294 332414 33058
rect 331794 13058 331826 13294
rect 332062 13058 332146 13294
rect 332382 13058 332414 13294
rect 331794 -1306 332414 13058
rect 331794 -1542 331826 -1306
rect 332062 -1542 332146 -1306
rect 332382 -1542 332414 -1306
rect 331794 -1626 332414 -1542
rect 331794 -1862 331826 -1626
rect 332062 -1862 332146 -1626
rect 332382 -1862 332414 -1626
rect 331794 -1894 332414 -1862
rect 332954 54274 333574 58000
rect 332954 54038 332986 54274
rect 333222 54038 333306 54274
rect 333542 54038 333574 54274
rect 332954 34274 333574 54038
rect 332954 34038 332986 34274
rect 333222 34038 333306 34274
rect 333542 34038 333574 34274
rect 332954 14274 333574 34038
rect 332954 14038 332986 14274
rect 333222 14038 333306 14274
rect 333542 14038 333574 14274
rect 329234 -4422 329266 -4186
rect 329502 -4422 329586 -4186
rect 329822 -4422 329854 -4186
rect 329234 -4506 329854 -4422
rect 329234 -4742 329266 -4506
rect 329502 -4742 329586 -4506
rect 329822 -4742 329854 -4506
rect 329234 -5734 329854 -4742
rect 322954 -7302 322986 -7066
rect 323222 -7302 323306 -7066
rect 323542 -7302 323574 -7066
rect 322954 -7386 323574 -7302
rect 322954 -7622 322986 -7386
rect 323222 -7622 323306 -7386
rect 323542 -7622 323574 -7386
rect 322954 -7654 323574 -7622
rect 332954 -6106 333574 14038
rect 335514 56954 336134 58000
rect 335514 56718 335546 56954
rect 335782 56718 335866 56954
rect 336102 56718 336134 56954
rect 335514 36954 336134 56718
rect 335514 36718 335546 36954
rect 335782 36718 335866 36954
rect 336102 36718 336134 36954
rect 335514 16954 336134 36718
rect 335514 16718 335546 16954
rect 335782 16718 335866 16954
rect 336102 16718 336134 16954
rect 335514 -3226 336134 16718
rect 335514 -3462 335546 -3226
rect 335782 -3462 335866 -3226
rect 336102 -3462 336134 -3226
rect 335514 -3546 336134 -3462
rect 335514 -3782 335546 -3546
rect 335782 -3782 335866 -3546
rect 336102 -3782 336134 -3546
rect 335514 -3814 336134 -3782
rect 339234 40614 339854 58000
rect 339234 40378 339266 40614
rect 339502 40378 339586 40614
rect 339822 40378 339854 40614
rect 339234 20614 339854 40378
rect 339234 20378 339266 20614
rect 339502 20378 339586 20614
rect 339822 20378 339854 20614
rect 339234 -5146 339854 20378
rect 341794 43294 342414 58000
rect 341794 43058 341826 43294
rect 342062 43058 342146 43294
rect 342382 43058 342414 43294
rect 341794 23294 342414 43058
rect 341794 23058 341826 23294
rect 342062 23058 342146 23294
rect 342382 23058 342414 23294
rect 341794 3294 342414 23058
rect 341794 3058 341826 3294
rect 342062 3058 342146 3294
rect 342382 3058 342414 3294
rect 341794 -346 342414 3058
rect 341794 -582 341826 -346
rect 342062 -582 342146 -346
rect 342382 -582 342414 -346
rect 341794 -666 342414 -582
rect 341794 -902 341826 -666
rect 342062 -902 342146 -666
rect 342382 -902 342414 -666
rect 341794 -1894 342414 -902
rect 342954 44274 343574 58000
rect 342954 44038 342986 44274
rect 343222 44038 343306 44274
rect 343542 44038 343574 44274
rect 342954 24274 343574 44038
rect 342954 24038 342986 24274
rect 343222 24038 343306 24274
rect 343542 24038 343574 24274
rect 339234 -5382 339266 -5146
rect 339502 -5382 339586 -5146
rect 339822 -5382 339854 -5146
rect 339234 -5466 339854 -5382
rect 339234 -5702 339266 -5466
rect 339502 -5702 339586 -5466
rect 339822 -5702 339854 -5466
rect 339234 -5734 339854 -5702
rect 332954 -6342 332986 -6106
rect 333222 -6342 333306 -6106
rect 333542 -6342 333574 -6106
rect 332954 -6426 333574 -6342
rect 332954 -6662 332986 -6426
rect 333222 -6662 333306 -6426
rect 333542 -6662 333574 -6426
rect 332954 -7654 333574 -6662
rect 342954 -7066 343574 24038
rect 345514 46954 346134 58000
rect 345514 46718 345546 46954
rect 345782 46718 345866 46954
rect 346102 46718 346134 46954
rect 345514 26954 346134 46718
rect 345514 26718 345546 26954
rect 345782 26718 345866 26954
rect 346102 26718 346134 26954
rect 345514 6954 346134 26718
rect 345514 6718 345546 6954
rect 345782 6718 345866 6954
rect 346102 6718 346134 6954
rect 345514 -2266 346134 6718
rect 345514 -2502 345546 -2266
rect 345782 -2502 345866 -2266
rect 346102 -2502 346134 -2266
rect 345514 -2586 346134 -2502
rect 345514 -2822 345546 -2586
rect 345782 -2822 345866 -2586
rect 346102 -2822 346134 -2586
rect 345514 -3814 346134 -2822
rect 349234 50614 349854 58000
rect 349234 50378 349266 50614
rect 349502 50378 349586 50614
rect 349822 50378 349854 50614
rect 349234 30614 349854 50378
rect 349234 30378 349266 30614
rect 349502 30378 349586 30614
rect 349822 30378 349854 30614
rect 349234 10614 349854 30378
rect 349234 10378 349266 10614
rect 349502 10378 349586 10614
rect 349822 10378 349854 10614
rect 349234 -4186 349854 10378
rect 351794 53294 352414 58000
rect 351794 53058 351826 53294
rect 352062 53058 352146 53294
rect 352382 53058 352414 53294
rect 351794 33294 352414 53058
rect 351794 33058 351826 33294
rect 352062 33058 352146 33294
rect 352382 33058 352414 33294
rect 351794 13294 352414 33058
rect 351794 13058 351826 13294
rect 352062 13058 352146 13294
rect 352382 13058 352414 13294
rect 351794 -1306 352414 13058
rect 351794 -1542 351826 -1306
rect 352062 -1542 352146 -1306
rect 352382 -1542 352414 -1306
rect 351794 -1626 352414 -1542
rect 351794 -1862 351826 -1626
rect 352062 -1862 352146 -1626
rect 352382 -1862 352414 -1626
rect 351794 -1894 352414 -1862
rect 352954 54274 353574 58000
rect 352954 54038 352986 54274
rect 353222 54038 353306 54274
rect 353542 54038 353574 54274
rect 352954 34274 353574 54038
rect 352954 34038 352986 34274
rect 353222 34038 353306 34274
rect 353542 34038 353574 34274
rect 352954 14274 353574 34038
rect 352954 14038 352986 14274
rect 353222 14038 353306 14274
rect 353542 14038 353574 14274
rect 349234 -4422 349266 -4186
rect 349502 -4422 349586 -4186
rect 349822 -4422 349854 -4186
rect 349234 -4506 349854 -4422
rect 349234 -4742 349266 -4506
rect 349502 -4742 349586 -4506
rect 349822 -4742 349854 -4506
rect 349234 -5734 349854 -4742
rect 342954 -7302 342986 -7066
rect 343222 -7302 343306 -7066
rect 343542 -7302 343574 -7066
rect 342954 -7386 343574 -7302
rect 342954 -7622 342986 -7386
rect 343222 -7622 343306 -7386
rect 343542 -7622 343574 -7386
rect 342954 -7654 343574 -7622
rect 352954 -6106 353574 14038
rect 355514 56954 356134 58000
rect 355514 56718 355546 56954
rect 355782 56718 355866 56954
rect 356102 56718 356134 56954
rect 355514 36954 356134 56718
rect 355514 36718 355546 36954
rect 355782 36718 355866 36954
rect 356102 36718 356134 36954
rect 355514 16954 356134 36718
rect 355514 16718 355546 16954
rect 355782 16718 355866 16954
rect 356102 16718 356134 16954
rect 355514 -3226 356134 16718
rect 355514 -3462 355546 -3226
rect 355782 -3462 355866 -3226
rect 356102 -3462 356134 -3226
rect 355514 -3546 356134 -3462
rect 355514 -3782 355546 -3546
rect 355782 -3782 355866 -3546
rect 356102 -3782 356134 -3546
rect 355514 -3814 356134 -3782
rect 359234 40614 359854 58000
rect 359234 40378 359266 40614
rect 359502 40378 359586 40614
rect 359822 40378 359854 40614
rect 359234 20614 359854 40378
rect 359234 20378 359266 20614
rect 359502 20378 359586 20614
rect 359822 20378 359854 20614
rect 359234 -5146 359854 20378
rect 361794 43294 362414 58000
rect 361794 43058 361826 43294
rect 362062 43058 362146 43294
rect 362382 43058 362414 43294
rect 361794 23294 362414 43058
rect 361794 23058 361826 23294
rect 362062 23058 362146 23294
rect 362382 23058 362414 23294
rect 361794 3294 362414 23058
rect 361794 3058 361826 3294
rect 362062 3058 362146 3294
rect 362382 3058 362414 3294
rect 361794 -346 362414 3058
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 362954 44274 363574 58000
rect 362954 44038 362986 44274
rect 363222 44038 363306 44274
rect 363542 44038 363574 44274
rect 362954 24274 363574 44038
rect 362954 24038 362986 24274
rect 363222 24038 363306 24274
rect 363542 24038 363574 24274
rect 359234 -5382 359266 -5146
rect 359502 -5382 359586 -5146
rect 359822 -5382 359854 -5146
rect 359234 -5466 359854 -5382
rect 359234 -5702 359266 -5466
rect 359502 -5702 359586 -5466
rect 359822 -5702 359854 -5466
rect 359234 -5734 359854 -5702
rect 352954 -6342 352986 -6106
rect 353222 -6342 353306 -6106
rect 353542 -6342 353574 -6106
rect 352954 -6426 353574 -6342
rect 352954 -6662 352986 -6426
rect 353222 -6662 353306 -6426
rect 353542 -6662 353574 -6426
rect 352954 -7654 353574 -6662
rect 362954 -7066 363574 24038
rect 365514 46954 366134 58000
rect 365514 46718 365546 46954
rect 365782 46718 365866 46954
rect 366102 46718 366134 46954
rect 365514 26954 366134 46718
rect 365514 26718 365546 26954
rect 365782 26718 365866 26954
rect 366102 26718 366134 26954
rect 365514 6954 366134 26718
rect 365514 6718 365546 6954
rect 365782 6718 365866 6954
rect 366102 6718 366134 6954
rect 365514 -2266 366134 6718
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 50614 369854 58000
rect 369234 50378 369266 50614
rect 369502 50378 369586 50614
rect 369822 50378 369854 50614
rect 369234 30614 369854 50378
rect 369234 30378 369266 30614
rect 369502 30378 369586 30614
rect 369822 30378 369854 30614
rect 369234 10614 369854 30378
rect 369234 10378 369266 10614
rect 369502 10378 369586 10614
rect 369822 10378 369854 10614
rect 369234 -4186 369854 10378
rect 371794 53294 372414 58000
rect 371794 53058 371826 53294
rect 372062 53058 372146 53294
rect 372382 53058 372414 53294
rect 371794 33294 372414 53058
rect 371794 33058 371826 33294
rect 372062 33058 372146 33294
rect 372382 33058 372414 33294
rect 371794 13294 372414 33058
rect 371794 13058 371826 13294
rect 372062 13058 372146 13294
rect 372382 13058 372414 13294
rect 371794 -1306 372414 13058
rect 371794 -1542 371826 -1306
rect 372062 -1542 372146 -1306
rect 372382 -1542 372414 -1306
rect 371794 -1626 372414 -1542
rect 371794 -1862 371826 -1626
rect 372062 -1862 372146 -1626
rect 372382 -1862 372414 -1626
rect 371794 -1894 372414 -1862
rect 372954 54274 373574 58000
rect 372954 54038 372986 54274
rect 373222 54038 373306 54274
rect 373542 54038 373574 54274
rect 372954 34274 373574 54038
rect 372954 34038 372986 34274
rect 373222 34038 373306 34274
rect 373542 34038 373574 34274
rect 372954 14274 373574 34038
rect 372954 14038 372986 14274
rect 373222 14038 373306 14274
rect 373542 14038 373574 14274
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 362954 -7302 362986 -7066
rect 363222 -7302 363306 -7066
rect 363542 -7302 363574 -7066
rect 362954 -7386 363574 -7302
rect 362954 -7622 362986 -7386
rect 363222 -7622 363306 -7386
rect 363542 -7622 363574 -7386
rect 362954 -7654 363574 -7622
rect 372954 -6106 373574 14038
rect 375514 56954 376134 58000
rect 375514 56718 375546 56954
rect 375782 56718 375866 56954
rect 376102 56718 376134 56954
rect 375514 36954 376134 56718
rect 375514 36718 375546 36954
rect 375782 36718 375866 36954
rect 376102 36718 376134 36954
rect 375514 16954 376134 36718
rect 375514 16718 375546 16954
rect 375782 16718 375866 16954
rect 376102 16718 376134 16954
rect 375514 -3226 376134 16718
rect 375514 -3462 375546 -3226
rect 375782 -3462 375866 -3226
rect 376102 -3462 376134 -3226
rect 375514 -3546 376134 -3462
rect 375514 -3782 375546 -3546
rect 375782 -3782 375866 -3546
rect 376102 -3782 376134 -3546
rect 375514 -3814 376134 -3782
rect 379234 40614 379854 58000
rect 379234 40378 379266 40614
rect 379502 40378 379586 40614
rect 379822 40378 379854 40614
rect 379234 20614 379854 40378
rect 379234 20378 379266 20614
rect 379502 20378 379586 20614
rect 379822 20378 379854 20614
rect 379234 -5146 379854 20378
rect 381794 43294 382414 58000
rect 381794 43058 381826 43294
rect 382062 43058 382146 43294
rect 382382 43058 382414 43294
rect 381794 23294 382414 43058
rect 381794 23058 381826 23294
rect 382062 23058 382146 23294
rect 382382 23058 382414 23294
rect 381794 3294 382414 23058
rect 381794 3058 381826 3294
rect 382062 3058 382146 3294
rect 382382 3058 382414 3294
rect 381794 -346 382414 3058
rect 381794 -582 381826 -346
rect 382062 -582 382146 -346
rect 382382 -582 382414 -346
rect 381794 -666 382414 -582
rect 381794 -902 381826 -666
rect 382062 -902 382146 -666
rect 382382 -902 382414 -666
rect 381794 -1894 382414 -902
rect 382954 44274 383574 58000
rect 382954 44038 382986 44274
rect 383222 44038 383306 44274
rect 383542 44038 383574 44274
rect 382954 24274 383574 44038
rect 382954 24038 382986 24274
rect 383222 24038 383306 24274
rect 383542 24038 383574 24274
rect 379234 -5382 379266 -5146
rect 379502 -5382 379586 -5146
rect 379822 -5382 379854 -5146
rect 379234 -5466 379854 -5382
rect 379234 -5702 379266 -5466
rect 379502 -5702 379586 -5466
rect 379822 -5702 379854 -5466
rect 379234 -5734 379854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 382954 -7066 383574 24038
rect 385514 46954 386134 58000
rect 385514 46718 385546 46954
rect 385782 46718 385866 46954
rect 386102 46718 386134 46954
rect 385514 26954 386134 46718
rect 385514 26718 385546 26954
rect 385782 26718 385866 26954
rect 386102 26718 386134 26954
rect 385514 6954 386134 26718
rect 385514 6718 385546 6954
rect 385782 6718 385866 6954
rect 386102 6718 386134 6954
rect 385514 -2266 386134 6718
rect 385514 -2502 385546 -2266
rect 385782 -2502 385866 -2266
rect 386102 -2502 386134 -2266
rect 385514 -2586 386134 -2502
rect 385514 -2822 385546 -2586
rect 385782 -2822 385866 -2586
rect 386102 -2822 386134 -2586
rect 385514 -3814 386134 -2822
rect 389234 50614 389854 58000
rect 389234 50378 389266 50614
rect 389502 50378 389586 50614
rect 389822 50378 389854 50614
rect 389234 30614 389854 50378
rect 389234 30378 389266 30614
rect 389502 30378 389586 30614
rect 389822 30378 389854 30614
rect 389234 10614 389854 30378
rect 389234 10378 389266 10614
rect 389502 10378 389586 10614
rect 389822 10378 389854 10614
rect 389234 -4186 389854 10378
rect 391794 53294 392414 58000
rect 391794 53058 391826 53294
rect 392062 53058 392146 53294
rect 392382 53058 392414 53294
rect 391794 33294 392414 53058
rect 391794 33058 391826 33294
rect 392062 33058 392146 33294
rect 392382 33058 392414 33294
rect 391794 13294 392414 33058
rect 391794 13058 391826 13294
rect 392062 13058 392146 13294
rect 392382 13058 392414 13294
rect 391794 -1306 392414 13058
rect 391794 -1542 391826 -1306
rect 392062 -1542 392146 -1306
rect 392382 -1542 392414 -1306
rect 391794 -1626 392414 -1542
rect 391794 -1862 391826 -1626
rect 392062 -1862 392146 -1626
rect 392382 -1862 392414 -1626
rect 391794 -1894 392414 -1862
rect 392954 54274 393574 58000
rect 392954 54038 392986 54274
rect 393222 54038 393306 54274
rect 393542 54038 393574 54274
rect 392954 34274 393574 54038
rect 392954 34038 392986 34274
rect 393222 34038 393306 34274
rect 393542 34038 393574 34274
rect 392954 14274 393574 34038
rect 392954 14038 392986 14274
rect 393222 14038 393306 14274
rect 393542 14038 393574 14274
rect 389234 -4422 389266 -4186
rect 389502 -4422 389586 -4186
rect 389822 -4422 389854 -4186
rect 389234 -4506 389854 -4422
rect 389234 -4742 389266 -4506
rect 389502 -4742 389586 -4506
rect 389822 -4742 389854 -4506
rect 389234 -5734 389854 -4742
rect 382954 -7302 382986 -7066
rect 383222 -7302 383306 -7066
rect 383542 -7302 383574 -7066
rect 382954 -7386 383574 -7302
rect 382954 -7622 382986 -7386
rect 383222 -7622 383306 -7386
rect 383542 -7622 383574 -7386
rect 382954 -7654 383574 -7622
rect 392954 -6106 393574 14038
rect 395514 56954 396134 58000
rect 395514 56718 395546 56954
rect 395782 56718 395866 56954
rect 396102 56718 396134 56954
rect 395514 36954 396134 56718
rect 395514 36718 395546 36954
rect 395782 36718 395866 36954
rect 396102 36718 396134 36954
rect 395514 16954 396134 36718
rect 395514 16718 395546 16954
rect 395782 16718 395866 16954
rect 396102 16718 396134 16954
rect 395514 -3226 396134 16718
rect 395514 -3462 395546 -3226
rect 395782 -3462 395866 -3226
rect 396102 -3462 396134 -3226
rect 395514 -3546 396134 -3462
rect 395514 -3782 395546 -3546
rect 395782 -3782 395866 -3546
rect 396102 -3782 396134 -3546
rect 395514 -3814 396134 -3782
rect 399234 40614 399854 58000
rect 399234 40378 399266 40614
rect 399502 40378 399586 40614
rect 399822 40378 399854 40614
rect 399234 20614 399854 40378
rect 399234 20378 399266 20614
rect 399502 20378 399586 20614
rect 399822 20378 399854 20614
rect 399234 -5146 399854 20378
rect 401794 43294 402414 58000
rect 401794 43058 401826 43294
rect 402062 43058 402146 43294
rect 402382 43058 402414 43294
rect 401794 23294 402414 43058
rect 401794 23058 401826 23294
rect 402062 23058 402146 23294
rect 402382 23058 402414 23294
rect 401794 3294 402414 23058
rect 401794 3058 401826 3294
rect 402062 3058 402146 3294
rect 402382 3058 402414 3294
rect 401794 -346 402414 3058
rect 401794 -582 401826 -346
rect 402062 -582 402146 -346
rect 402382 -582 402414 -346
rect 401794 -666 402414 -582
rect 401794 -902 401826 -666
rect 402062 -902 402146 -666
rect 402382 -902 402414 -666
rect 401794 -1894 402414 -902
rect 402954 44274 403574 58000
rect 402954 44038 402986 44274
rect 403222 44038 403306 44274
rect 403542 44038 403574 44274
rect 402954 24274 403574 44038
rect 402954 24038 402986 24274
rect 403222 24038 403306 24274
rect 403542 24038 403574 24274
rect 399234 -5382 399266 -5146
rect 399502 -5382 399586 -5146
rect 399822 -5382 399854 -5146
rect 399234 -5466 399854 -5382
rect 399234 -5702 399266 -5466
rect 399502 -5702 399586 -5466
rect 399822 -5702 399854 -5466
rect 399234 -5734 399854 -5702
rect 392954 -6342 392986 -6106
rect 393222 -6342 393306 -6106
rect 393542 -6342 393574 -6106
rect 392954 -6426 393574 -6342
rect 392954 -6662 392986 -6426
rect 393222 -6662 393306 -6426
rect 393542 -6662 393574 -6426
rect 392954 -7654 393574 -6662
rect 402954 -7066 403574 24038
rect 405514 46954 406134 58000
rect 405514 46718 405546 46954
rect 405782 46718 405866 46954
rect 406102 46718 406134 46954
rect 405514 26954 406134 46718
rect 405514 26718 405546 26954
rect 405782 26718 405866 26954
rect 406102 26718 406134 26954
rect 405514 6954 406134 26718
rect 405514 6718 405546 6954
rect 405782 6718 405866 6954
rect 406102 6718 406134 6954
rect 405514 -2266 406134 6718
rect 405514 -2502 405546 -2266
rect 405782 -2502 405866 -2266
rect 406102 -2502 406134 -2266
rect 405514 -2586 406134 -2502
rect 405514 -2822 405546 -2586
rect 405782 -2822 405866 -2586
rect 406102 -2822 406134 -2586
rect 405514 -3814 406134 -2822
rect 409234 50614 409854 58000
rect 409234 50378 409266 50614
rect 409502 50378 409586 50614
rect 409822 50378 409854 50614
rect 409234 30614 409854 50378
rect 409234 30378 409266 30614
rect 409502 30378 409586 30614
rect 409822 30378 409854 30614
rect 409234 10614 409854 30378
rect 409234 10378 409266 10614
rect 409502 10378 409586 10614
rect 409822 10378 409854 10614
rect 409234 -4186 409854 10378
rect 411794 53294 412414 58000
rect 411794 53058 411826 53294
rect 412062 53058 412146 53294
rect 412382 53058 412414 53294
rect 411794 33294 412414 53058
rect 411794 33058 411826 33294
rect 412062 33058 412146 33294
rect 412382 33058 412414 33294
rect 411794 13294 412414 33058
rect 411794 13058 411826 13294
rect 412062 13058 412146 13294
rect 412382 13058 412414 13294
rect 411794 -1306 412414 13058
rect 411794 -1542 411826 -1306
rect 412062 -1542 412146 -1306
rect 412382 -1542 412414 -1306
rect 411794 -1626 412414 -1542
rect 411794 -1862 411826 -1626
rect 412062 -1862 412146 -1626
rect 412382 -1862 412414 -1626
rect 411794 -1894 412414 -1862
rect 412954 54274 413574 58000
rect 412954 54038 412986 54274
rect 413222 54038 413306 54274
rect 413542 54038 413574 54274
rect 412954 34274 413574 54038
rect 412954 34038 412986 34274
rect 413222 34038 413306 34274
rect 413542 34038 413574 34274
rect 412954 14274 413574 34038
rect 412954 14038 412986 14274
rect 413222 14038 413306 14274
rect 413542 14038 413574 14274
rect 409234 -4422 409266 -4186
rect 409502 -4422 409586 -4186
rect 409822 -4422 409854 -4186
rect 409234 -4506 409854 -4422
rect 409234 -4742 409266 -4506
rect 409502 -4742 409586 -4506
rect 409822 -4742 409854 -4506
rect 409234 -5734 409854 -4742
rect 402954 -7302 402986 -7066
rect 403222 -7302 403306 -7066
rect 403542 -7302 403574 -7066
rect 402954 -7386 403574 -7302
rect 402954 -7622 402986 -7386
rect 403222 -7622 403306 -7386
rect 403542 -7622 403574 -7386
rect 402954 -7654 403574 -7622
rect 412954 -6106 413574 14038
rect 415514 56954 416134 58000
rect 415514 56718 415546 56954
rect 415782 56718 415866 56954
rect 416102 56718 416134 56954
rect 415514 36954 416134 56718
rect 415514 36718 415546 36954
rect 415782 36718 415866 36954
rect 416102 36718 416134 36954
rect 415514 16954 416134 36718
rect 415514 16718 415546 16954
rect 415782 16718 415866 16954
rect 416102 16718 416134 16954
rect 415514 -3226 416134 16718
rect 415514 -3462 415546 -3226
rect 415782 -3462 415866 -3226
rect 416102 -3462 416134 -3226
rect 415514 -3546 416134 -3462
rect 415514 -3782 415546 -3546
rect 415782 -3782 415866 -3546
rect 416102 -3782 416134 -3546
rect 415514 -3814 416134 -3782
rect 419234 40614 419854 58000
rect 419234 40378 419266 40614
rect 419502 40378 419586 40614
rect 419822 40378 419854 40614
rect 419234 20614 419854 40378
rect 419234 20378 419266 20614
rect 419502 20378 419586 20614
rect 419822 20378 419854 20614
rect 419234 -5146 419854 20378
rect 421794 43294 422414 58000
rect 421794 43058 421826 43294
rect 422062 43058 422146 43294
rect 422382 43058 422414 43294
rect 421794 23294 422414 43058
rect 421794 23058 421826 23294
rect 422062 23058 422146 23294
rect 422382 23058 422414 23294
rect 421794 3294 422414 23058
rect 421794 3058 421826 3294
rect 422062 3058 422146 3294
rect 422382 3058 422414 3294
rect 421794 -346 422414 3058
rect 421794 -582 421826 -346
rect 422062 -582 422146 -346
rect 422382 -582 422414 -346
rect 421794 -666 422414 -582
rect 421794 -902 421826 -666
rect 422062 -902 422146 -666
rect 422382 -902 422414 -666
rect 421794 -1894 422414 -902
rect 422954 44274 423574 58000
rect 422954 44038 422986 44274
rect 423222 44038 423306 44274
rect 423542 44038 423574 44274
rect 422954 24274 423574 44038
rect 422954 24038 422986 24274
rect 423222 24038 423306 24274
rect 423542 24038 423574 24274
rect 419234 -5382 419266 -5146
rect 419502 -5382 419586 -5146
rect 419822 -5382 419854 -5146
rect 419234 -5466 419854 -5382
rect 419234 -5702 419266 -5466
rect 419502 -5702 419586 -5466
rect 419822 -5702 419854 -5466
rect 419234 -5734 419854 -5702
rect 412954 -6342 412986 -6106
rect 413222 -6342 413306 -6106
rect 413542 -6342 413574 -6106
rect 412954 -6426 413574 -6342
rect 412954 -6662 412986 -6426
rect 413222 -6662 413306 -6426
rect 413542 -6662 413574 -6426
rect 412954 -7654 413574 -6662
rect 422954 -7066 423574 24038
rect 425514 46954 426134 58000
rect 425514 46718 425546 46954
rect 425782 46718 425866 46954
rect 426102 46718 426134 46954
rect 425514 26954 426134 46718
rect 425514 26718 425546 26954
rect 425782 26718 425866 26954
rect 426102 26718 426134 26954
rect 425514 6954 426134 26718
rect 425514 6718 425546 6954
rect 425782 6718 425866 6954
rect 426102 6718 426134 6954
rect 425514 -2266 426134 6718
rect 425514 -2502 425546 -2266
rect 425782 -2502 425866 -2266
rect 426102 -2502 426134 -2266
rect 425514 -2586 426134 -2502
rect 425514 -2822 425546 -2586
rect 425782 -2822 425866 -2586
rect 426102 -2822 426134 -2586
rect 425514 -3814 426134 -2822
rect 429234 50614 429854 58000
rect 429234 50378 429266 50614
rect 429502 50378 429586 50614
rect 429822 50378 429854 50614
rect 429234 30614 429854 50378
rect 429234 30378 429266 30614
rect 429502 30378 429586 30614
rect 429822 30378 429854 30614
rect 429234 10614 429854 30378
rect 429234 10378 429266 10614
rect 429502 10378 429586 10614
rect 429822 10378 429854 10614
rect 429234 -4186 429854 10378
rect 431794 53294 432414 58000
rect 431794 53058 431826 53294
rect 432062 53058 432146 53294
rect 432382 53058 432414 53294
rect 431794 33294 432414 53058
rect 431794 33058 431826 33294
rect 432062 33058 432146 33294
rect 432382 33058 432414 33294
rect 431794 13294 432414 33058
rect 431794 13058 431826 13294
rect 432062 13058 432146 13294
rect 432382 13058 432414 13294
rect 431794 -1306 432414 13058
rect 431794 -1542 431826 -1306
rect 432062 -1542 432146 -1306
rect 432382 -1542 432414 -1306
rect 431794 -1626 432414 -1542
rect 431794 -1862 431826 -1626
rect 432062 -1862 432146 -1626
rect 432382 -1862 432414 -1626
rect 431794 -1894 432414 -1862
rect 432954 54274 433574 58000
rect 432954 54038 432986 54274
rect 433222 54038 433306 54274
rect 433542 54038 433574 54274
rect 432954 34274 433574 54038
rect 432954 34038 432986 34274
rect 433222 34038 433306 34274
rect 433542 34038 433574 34274
rect 432954 14274 433574 34038
rect 432954 14038 432986 14274
rect 433222 14038 433306 14274
rect 433542 14038 433574 14274
rect 429234 -4422 429266 -4186
rect 429502 -4422 429586 -4186
rect 429822 -4422 429854 -4186
rect 429234 -4506 429854 -4422
rect 429234 -4742 429266 -4506
rect 429502 -4742 429586 -4506
rect 429822 -4742 429854 -4506
rect 429234 -5734 429854 -4742
rect 422954 -7302 422986 -7066
rect 423222 -7302 423306 -7066
rect 423542 -7302 423574 -7066
rect 422954 -7386 423574 -7302
rect 422954 -7622 422986 -7386
rect 423222 -7622 423306 -7386
rect 423542 -7622 423574 -7386
rect 422954 -7654 423574 -7622
rect 432954 -6106 433574 14038
rect 435514 56954 436134 58000
rect 435514 56718 435546 56954
rect 435782 56718 435866 56954
rect 436102 56718 436134 56954
rect 435514 36954 436134 56718
rect 435514 36718 435546 36954
rect 435782 36718 435866 36954
rect 436102 36718 436134 36954
rect 435514 16954 436134 36718
rect 435514 16718 435546 16954
rect 435782 16718 435866 16954
rect 436102 16718 436134 16954
rect 435514 -3226 436134 16718
rect 435514 -3462 435546 -3226
rect 435782 -3462 435866 -3226
rect 436102 -3462 436134 -3226
rect 435514 -3546 436134 -3462
rect 435514 -3782 435546 -3546
rect 435782 -3782 435866 -3546
rect 436102 -3782 436134 -3546
rect 435514 -3814 436134 -3782
rect 439234 40614 439854 58000
rect 439234 40378 439266 40614
rect 439502 40378 439586 40614
rect 439822 40378 439854 40614
rect 439234 20614 439854 40378
rect 439234 20378 439266 20614
rect 439502 20378 439586 20614
rect 439822 20378 439854 20614
rect 439234 -5146 439854 20378
rect 441794 43294 442414 58000
rect 441794 43058 441826 43294
rect 442062 43058 442146 43294
rect 442382 43058 442414 43294
rect 441794 23294 442414 43058
rect 441794 23058 441826 23294
rect 442062 23058 442146 23294
rect 442382 23058 442414 23294
rect 441794 3294 442414 23058
rect 441794 3058 441826 3294
rect 442062 3058 442146 3294
rect 442382 3058 442414 3294
rect 441794 -346 442414 3058
rect 441794 -582 441826 -346
rect 442062 -582 442146 -346
rect 442382 -582 442414 -346
rect 441794 -666 442414 -582
rect 441794 -902 441826 -666
rect 442062 -902 442146 -666
rect 442382 -902 442414 -666
rect 441794 -1894 442414 -902
rect 442954 44274 443574 58000
rect 442954 44038 442986 44274
rect 443222 44038 443306 44274
rect 443542 44038 443574 44274
rect 442954 24274 443574 44038
rect 442954 24038 442986 24274
rect 443222 24038 443306 24274
rect 443542 24038 443574 24274
rect 439234 -5382 439266 -5146
rect 439502 -5382 439586 -5146
rect 439822 -5382 439854 -5146
rect 439234 -5466 439854 -5382
rect 439234 -5702 439266 -5466
rect 439502 -5702 439586 -5466
rect 439822 -5702 439854 -5466
rect 439234 -5734 439854 -5702
rect 432954 -6342 432986 -6106
rect 433222 -6342 433306 -6106
rect 433542 -6342 433574 -6106
rect 432954 -6426 433574 -6342
rect 432954 -6662 432986 -6426
rect 433222 -6662 433306 -6426
rect 433542 -6662 433574 -6426
rect 432954 -7654 433574 -6662
rect 442954 -7066 443574 24038
rect 445514 46954 446134 58000
rect 445514 46718 445546 46954
rect 445782 46718 445866 46954
rect 446102 46718 446134 46954
rect 445514 26954 446134 46718
rect 445514 26718 445546 26954
rect 445782 26718 445866 26954
rect 446102 26718 446134 26954
rect 445514 6954 446134 26718
rect 445514 6718 445546 6954
rect 445782 6718 445866 6954
rect 446102 6718 446134 6954
rect 445514 -2266 446134 6718
rect 445514 -2502 445546 -2266
rect 445782 -2502 445866 -2266
rect 446102 -2502 446134 -2266
rect 445514 -2586 446134 -2502
rect 445514 -2822 445546 -2586
rect 445782 -2822 445866 -2586
rect 446102 -2822 446134 -2586
rect 445514 -3814 446134 -2822
rect 449234 50614 449854 58000
rect 449234 50378 449266 50614
rect 449502 50378 449586 50614
rect 449822 50378 449854 50614
rect 449234 30614 449854 50378
rect 449234 30378 449266 30614
rect 449502 30378 449586 30614
rect 449822 30378 449854 30614
rect 449234 10614 449854 30378
rect 449234 10378 449266 10614
rect 449502 10378 449586 10614
rect 449822 10378 449854 10614
rect 449234 -4186 449854 10378
rect 451794 53294 452414 58000
rect 451794 53058 451826 53294
rect 452062 53058 452146 53294
rect 452382 53058 452414 53294
rect 451794 33294 452414 53058
rect 451794 33058 451826 33294
rect 452062 33058 452146 33294
rect 452382 33058 452414 33294
rect 451794 13294 452414 33058
rect 451794 13058 451826 13294
rect 452062 13058 452146 13294
rect 452382 13058 452414 13294
rect 451794 -1306 452414 13058
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 452954 54274 453574 58000
rect 452954 54038 452986 54274
rect 453222 54038 453306 54274
rect 453542 54038 453574 54274
rect 452954 34274 453574 54038
rect 452954 34038 452986 34274
rect 453222 34038 453306 34274
rect 453542 34038 453574 34274
rect 452954 14274 453574 34038
rect 452954 14038 452986 14274
rect 453222 14038 453306 14274
rect 453542 14038 453574 14274
rect 449234 -4422 449266 -4186
rect 449502 -4422 449586 -4186
rect 449822 -4422 449854 -4186
rect 449234 -4506 449854 -4422
rect 449234 -4742 449266 -4506
rect 449502 -4742 449586 -4506
rect 449822 -4742 449854 -4506
rect 449234 -5734 449854 -4742
rect 442954 -7302 442986 -7066
rect 443222 -7302 443306 -7066
rect 443542 -7302 443574 -7066
rect 442954 -7386 443574 -7302
rect 442954 -7622 442986 -7386
rect 443222 -7622 443306 -7386
rect 443542 -7622 443574 -7386
rect 442954 -7654 443574 -7622
rect 452954 -6106 453574 14038
rect 455514 56954 456134 58000
rect 455514 56718 455546 56954
rect 455782 56718 455866 56954
rect 456102 56718 456134 56954
rect 455514 36954 456134 56718
rect 455514 36718 455546 36954
rect 455782 36718 455866 36954
rect 456102 36718 456134 36954
rect 455514 16954 456134 36718
rect 455514 16718 455546 16954
rect 455782 16718 455866 16954
rect 456102 16718 456134 16954
rect 455514 -3226 456134 16718
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 40614 459854 58000
rect 459234 40378 459266 40614
rect 459502 40378 459586 40614
rect 459822 40378 459854 40614
rect 459234 20614 459854 40378
rect 459234 20378 459266 20614
rect 459502 20378 459586 20614
rect 459822 20378 459854 20614
rect 459234 -5146 459854 20378
rect 461794 43294 462414 58000
rect 461794 43058 461826 43294
rect 462062 43058 462146 43294
rect 462382 43058 462414 43294
rect 461794 23294 462414 43058
rect 461794 23058 461826 23294
rect 462062 23058 462146 23294
rect 462382 23058 462414 23294
rect 461794 3294 462414 23058
rect 461794 3058 461826 3294
rect 462062 3058 462146 3294
rect 462382 3058 462414 3294
rect 461794 -346 462414 3058
rect 461794 -582 461826 -346
rect 462062 -582 462146 -346
rect 462382 -582 462414 -346
rect 461794 -666 462414 -582
rect 461794 -902 461826 -666
rect 462062 -902 462146 -666
rect 462382 -902 462414 -666
rect 461794 -1894 462414 -902
rect 462954 44274 463574 58000
rect 462954 44038 462986 44274
rect 463222 44038 463306 44274
rect 463542 44038 463574 44274
rect 462954 24274 463574 44038
rect 462954 24038 462986 24274
rect 463222 24038 463306 24274
rect 463542 24038 463574 24274
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 452954 -6342 452986 -6106
rect 453222 -6342 453306 -6106
rect 453542 -6342 453574 -6106
rect 452954 -6426 453574 -6342
rect 452954 -6662 452986 -6426
rect 453222 -6662 453306 -6426
rect 453542 -6662 453574 -6426
rect 452954 -7654 453574 -6662
rect 462954 -7066 463574 24038
rect 465514 46954 466134 58000
rect 465514 46718 465546 46954
rect 465782 46718 465866 46954
rect 466102 46718 466134 46954
rect 465514 26954 466134 46718
rect 465514 26718 465546 26954
rect 465782 26718 465866 26954
rect 466102 26718 466134 26954
rect 465514 6954 466134 26718
rect 465514 6718 465546 6954
rect 465782 6718 465866 6954
rect 466102 6718 466134 6954
rect 465514 -2266 466134 6718
rect 465514 -2502 465546 -2266
rect 465782 -2502 465866 -2266
rect 466102 -2502 466134 -2266
rect 465514 -2586 466134 -2502
rect 465514 -2822 465546 -2586
rect 465782 -2822 465866 -2586
rect 466102 -2822 466134 -2586
rect 465514 -3814 466134 -2822
rect 469234 50614 469854 58000
rect 469234 50378 469266 50614
rect 469502 50378 469586 50614
rect 469822 50378 469854 50614
rect 469234 30614 469854 50378
rect 469234 30378 469266 30614
rect 469502 30378 469586 30614
rect 469822 30378 469854 30614
rect 469234 10614 469854 30378
rect 469234 10378 469266 10614
rect 469502 10378 469586 10614
rect 469822 10378 469854 10614
rect 469234 -4186 469854 10378
rect 471794 53294 472414 58000
rect 471794 53058 471826 53294
rect 472062 53058 472146 53294
rect 472382 53058 472414 53294
rect 471794 33294 472414 53058
rect 471794 33058 471826 33294
rect 472062 33058 472146 33294
rect 472382 33058 472414 33294
rect 471794 13294 472414 33058
rect 471794 13058 471826 13294
rect 472062 13058 472146 13294
rect 472382 13058 472414 13294
rect 471794 -1306 472414 13058
rect 471794 -1542 471826 -1306
rect 472062 -1542 472146 -1306
rect 472382 -1542 472414 -1306
rect 471794 -1626 472414 -1542
rect 471794 -1862 471826 -1626
rect 472062 -1862 472146 -1626
rect 472382 -1862 472414 -1626
rect 471794 -1894 472414 -1862
rect 472954 54274 473574 58000
rect 472954 54038 472986 54274
rect 473222 54038 473306 54274
rect 473542 54038 473574 54274
rect 472954 34274 473574 54038
rect 472954 34038 472986 34274
rect 473222 34038 473306 34274
rect 473542 34038 473574 34274
rect 472954 14274 473574 34038
rect 472954 14038 472986 14274
rect 473222 14038 473306 14274
rect 473542 14038 473574 14274
rect 469234 -4422 469266 -4186
rect 469502 -4422 469586 -4186
rect 469822 -4422 469854 -4186
rect 469234 -4506 469854 -4422
rect 469234 -4742 469266 -4506
rect 469502 -4742 469586 -4506
rect 469822 -4742 469854 -4506
rect 469234 -5734 469854 -4742
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 472954 -6106 473574 14038
rect 475514 56954 476134 58000
rect 475514 56718 475546 56954
rect 475782 56718 475866 56954
rect 476102 56718 476134 56954
rect 475514 36954 476134 56718
rect 475514 36718 475546 36954
rect 475782 36718 475866 36954
rect 476102 36718 476134 36954
rect 475514 16954 476134 36718
rect 475514 16718 475546 16954
rect 475782 16718 475866 16954
rect 476102 16718 476134 16954
rect 475514 -3226 476134 16718
rect 475514 -3462 475546 -3226
rect 475782 -3462 475866 -3226
rect 476102 -3462 476134 -3226
rect 475514 -3546 476134 -3462
rect 475514 -3782 475546 -3546
rect 475782 -3782 475866 -3546
rect 476102 -3782 476134 -3546
rect 475514 -3814 476134 -3782
rect 479234 40614 479854 58000
rect 479234 40378 479266 40614
rect 479502 40378 479586 40614
rect 479822 40378 479854 40614
rect 479234 20614 479854 40378
rect 479234 20378 479266 20614
rect 479502 20378 479586 20614
rect 479822 20378 479854 20614
rect 479234 -5146 479854 20378
rect 481794 43294 482414 58000
rect 481794 43058 481826 43294
rect 482062 43058 482146 43294
rect 482382 43058 482414 43294
rect 481794 23294 482414 43058
rect 481794 23058 481826 23294
rect 482062 23058 482146 23294
rect 482382 23058 482414 23294
rect 481794 3294 482414 23058
rect 481794 3058 481826 3294
rect 482062 3058 482146 3294
rect 482382 3058 482414 3294
rect 481794 -346 482414 3058
rect 481794 -582 481826 -346
rect 482062 -582 482146 -346
rect 482382 -582 482414 -346
rect 481794 -666 482414 -582
rect 481794 -902 481826 -666
rect 482062 -902 482146 -666
rect 482382 -902 482414 -666
rect 481794 -1894 482414 -902
rect 482954 44274 483574 58000
rect 482954 44038 482986 44274
rect 483222 44038 483306 44274
rect 483542 44038 483574 44274
rect 482954 24274 483574 44038
rect 482954 24038 482986 24274
rect 483222 24038 483306 24274
rect 483542 24038 483574 24274
rect 479234 -5382 479266 -5146
rect 479502 -5382 479586 -5146
rect 479822 -5382 479854 -5146
rect 479234 -5466 479854 -5382
rect 479234 -5702 479266 -5466
rect 479502 -5702 479586 -5466
rect 479822 -5702 479854 -5466
rect 479234 -5734 479854 -5702
rect 472954 -6342 472986 -6106
rect 473222 -6342 473306 -6106
rect 473542 -6342 473574 -6106
rect 472954 -6426 473574 -6342
rect 472954 -6662 472986 -6426
rect 473222 -6662 473306 -6426
rect 473542 -6662 473574 -6426
rect 472954 -7654 473574 -6662
rect 482954 -7066 483574 24038
rect 485514 46954 486134 58000
rect 485514 46718 485546 46954
rect 485782 46718 485866 46954
rect 486102 46718 486134 46954
rect 485514 26954 486134 46718
rect 485514 26718 485546 26954
rect 485782 26718 485866 26954
rect 486102 26718 486134 26954
rect 485514 6954 486134 26718
rect 485514 6718 485546 6954
rect 485782 6718 485866 6954
rect 486102 6718 486134 6954
rect 485514 -2266 486134 6718
rect 485514 -2502 485546 -2266
rect 485782 -2502 485866 -2266
rect 486102 -2502 486134 -2266
rect 485514 -2586 486134 -2502
rect 485514 -2822 485546 -2586
rect 485782 -2822 485866 -2586
rect 486102 -2822 486134 -2586
rect 485514 -3814 486134 -2822
rect 489234 50614 489854 58000
rect 489234 50378 489266 50614
rect 489502 50378 489586 50614
rect 489822 50378 489854 50614
rect 489234 30614 489854 50378
rect 489234 30378 489266 30614
rect 489502 30378 489586 30614
rect 489822 30378 489854 30614
rect 489234 10614 489854 30378
rect 489234 10378 489266 10614
rect 489502 10378 489586 10614
rect 489822 10378 489854 10614
rect 489234 -4186 489854 10378
rect 491794 53294 492414 58000
rect 491794 53058 491826 53294
rect 492062 53058 492146 53294
rect 492382 53058 492414 53294
rect 491794 33294 492414 53058
rect 491794 33058 491826 33294
rect 492062 33058 492146 33294
rect 492382 33058 492414 33294
rect 491794 13294 492414 33058
rect 491794 13058 491826 13294
rect 492062 13058 492146 13294
rect 492382 13058 492414 13294
rect 491794 -1306 492414 13058
rect 491794 -1542 491826 -1306
rect 492062 -1542 492146 -1306
rect 492382 -1542 492414 -1306
rect 491794 -1626 492414 -1542
rect 491794 -1862 491826 -1626
rect 492062 -1862 492146 -1626
rect 492382 -1862 492414 -1626
rect 491794 -1894 492414 -1862
rect 492954 54274 493574 58000
rect 492954 54038 492986 54274
rect 493222 54038 493306 54274
rect 493542 54038 493574 54274
rect 492954 34274 493574 54038
rect 492954 34038 492986 34274
rect 493222 34038 493306 34274
rect 493542 34038 493574 34274
rect 492954 14274 493574 34038
rect 492954 14038 492986 14274
rect 493222 14038 493306 14274
rect 493542 14038 493574 14274
rect 489234 -4422 489266 -4186
rect 489502 -4422 489586 -4186
rect 489822 -4422 489854 -4186
rect 489234 -4506 489854 -4422
rect 489234 -4742 489266 -4506
rect 489502 -4742 489586 -4506
rect 489822 -4742 489854 -4506
rect 489234 -5734 489854 -4742
rect 482954 -7302 482986 -7066
rect 483222 -7302 483306 -7066
rect 483542 -7302 483574 -7066
rect 482954 -7386 483574 -7302
rect 482954 -7622 482986 -7386
rect 483222 -7622 483306 -7386
rect 483542 -7622 483574 -7386
rect 482954 -7654 483574 -7622
rect 492954 -6106 493574 14038
rect 495514 56954 496134 58000
rect 495514 56718 495546 56954
rect 495782 56718 495866 56954
rect 496102 56718 496134 56954
rect 495514 36954 496134 56718
rect 495514 36718 495546 36954
rect 495782 36718 495866 36954
rect 496102 36718 496134 36954
rect 495514 16954 496134 36718
rect 495514 16718 495546 16954
rect 495782 16718 495866 16954
rect 496102 16718 496134 16954
rect 495514 -3226 496134 16718
rect 495514 -3462 495546 -3226
rect 495782 -3462 495866 -3226
rect 496102 -3462 496134 -3226
rect 495514 -3546 496134 -3462
rect 495514 -3782 495546 -3546
rect 495782 -3782 495866 -3546
rect 496102 -3782 496134 -3546
rect 495514 -3814 496134 -3782
rect 499234 40614 499854 58000
rect 499234 40378 499266 40614
rect 499502 40378 499586 40614
rect 499822 40378 499854 40614
rect 499234 20614 499854 40378
rect 499234 20378 499266 20614
rect 499502 20378 499586 20614
rect 499822 20378 499854 20614
rect 499234 -5146 499854 20378
rect 501794 43294 502414 58000
rect 501794 43058 501826 43294
rect 502062 43058 502146 43294
rect 502382 43058 502414 43294
rect 501794 23294 502414 43058
rect 501794 23058 501826 23294
rect 502062 23058 502146 23294
rect 502382 23058 502414 23294
rect 501794 3294 502414 23058
rect 501794 3058 501826 3294
rect 502062 3058 502146 3294
rect 502382 3058 502414 3294
rect 501794 -346 502414 3058
rect 501794 -582 501826 -346
rect 502062 -582 502146 -346
rect 502382 -582 502414 -346
rect 501794 -666 502414 -582
rect 501794 -902 501826 -666
rect 502062 -902 502146 -666
rect 502382 -902 502414 -666
rect 501794 -1894 502414 -902
rect 502954 44274 503574 58000
rect 502954 44038 502986 44274
rect 503222 44038 503306 44274
rect 503542 44038 503574 44274
rect 502954 24274 503574 44038
rect 502954 24038 502986 24274
rect 503222 24038 503306 24274
rect 503542 24038 503574 24274
rect 499234 -5382 499266 -5146
rect 499502 -5382 499586 -5146
rect 499822 -5382 499854 -5146
rect 499234 -5466 499854 -5382
rect 499234 -5702 499266 -5466
rect 499502 -5702 499586 -5466
rect 499822 -5702 499854 -5466
rect 499234 -5734 499854 -5702
rect 492954 -6342 492986 -6106
rect 493222 -6342 493306 -6106
rect 493542 -6342 493574 -6106
rect 492954 -6426 493574 -6342
rect 492954 -6662 492986 -6426
rect 493222 -6662 493306 -6426
rect 493542 -6662 493574 -6426
rect 492954 -7654 493574 -6662
rect 502954 -7066 503574 24038
rect 505514 46954 506134 58000
rect 505514 46718 505546 46954
rect 505782 46718 505866 46954
rect 506102 46718 506134 46954
rect 505514 26954 506134 46718
rect 505514 26718 505546 26954
rect 505782 26718 505866 26954
rect 506102 26718 506134 26954
rect 505514 6954 506134 26718
rect 505514 6718 505546 6954
rect 505782 6718 505866 6954
rect 506102 6718 506134 6954
rect 505514 -2266 506134 6718
rect 505514 -2502 505546 -2266
rect 505782 -2502 505866 -2266
rect 506102 -2502 506134 -2266
rect 505514 -2586 506134 -2502
rect 505514 -2822 505546 -2586
rect 505782 -2822 505866 -2586
rect 506102 -2822 506134 -2586
rect 505514 -3814 506134 -2822
rect 509234 50614 509854 58000
rect 509234 50378 509266 50614
rect 509502 50378 509586 50614
rect 509822 50378 509854 50614
rect 509234 30614 509854 50378
rect 509234 30378 509266 30614
rect 509502 30378 509586 30614
rect 509822 30378 509854 30614
rect 509234 10614 509854 30378
rect 509234 10378 509266 10614
rect 509502 10378 509586 10614
rect 509822 10378 509854 10614
rect 509234 -4186 509854 10378
rect 511794 53294 512414 58000
rect 511794 53058 511826 53294
rect 512062 53058 512146 53294
rect 512382 53058 512414 53294
rect 511794 33294 512414 53058
rect 511794 33058 511826 33294
rect 512062 33058 512146 33294
rect 512382 33058 512414 33294
rect 511794 13294 512414 33058
rect 511794 13058 511826 13294
rect 512062 13058 512146 13294
rect 512382 13058 512414 13294
rect 511794 -1306 512414 13058
rect 511794 -1542 511826 -1306
rect 512062 -1542 512146 -1306
rect 512382 -1542 512414 -1306
rect 511794 -1626 512414 -1542
rect 511794 -1862 511826 -1626
rect 512062 -1862 512146 -1626
rect 512382 -1862 512414 -1626
rect 511794 -1894 512414 -1862
rect 512954 54274 513574 58000
rect 512954 54038 512986 54274
rect 513222 54038 513306 54274
rect 513542 54038 513574 54274
rect 512954 34274 513574 54038
rect 512954 34038 512986 34274
rect 513222 34038 513306 34274
rect 513542 34038 513574 34274
rect 512954 14274 513574 34038
rect 512954 14038 512986 14274
rect 513222 14038 513306 14274
rect 513542 14038 513574 14274
rect 509234 -4422 509266 -4186
rect 509502 -4422 509586 -4186
rect 509822 -4422 509854 -4186
rect 509234 -4506 509854 -4422
rect 509234 -4742 509266 -4506
rect 509502 -4742 509586 -4506
rect 509822 -4742 509854 -4506
rect 509234 -5734 509854 -4742
rect 502954 -7302 502986 -7066
rect 503222 -7302 503306 -7066
rect 503542 -7302 503574 -7066
rect 502954 -7386 503574 -7302
rect 502954 -7622 502986 -7386
rect 503222 -7622 503306 -7386
rect 503542 -7622 503574 -7386
rect 502954 -7654 503574 -7622
rect 512954 -6106 513574 14038
rect 515514 56954 516134 58000
rect 515514 56718 515546 56954
rect 515782 56718 515866 56954
rect 516102 56718 516134 56954
rect 515514 36954 516134 56718
rect 515514 36718 515546 36954
rect 515782 36718 515866 36954
rect 516102 36718 516134 36954
rect 515514 16954 516134 36718
rect 515514 16718 515546 16954
rect 515782 16718 515866 16954
rect 516102 16718 516134 16954
rect 515514 -3226 516134 16718
rect 515514 -3462 515546 -3226
rect 515782 -3462 515866 -3226
rect 516102 -3462 516134 -3226
rect 515514 -3546 516134 -3462
rect 515514 -3782 515546 -3546
rect 515782 -3782 515866 -3546
rect 516102 -3782 516134 -3546
rect 515514 -3814 516134 -3782
rect 519234 40614 519854 58000
rect 519234 40378 519266 40614
rect 519502 40378 519586 40614
rect 519822 40378 519854 40614
rect 519234 20614 519854 40378
rect 519234 20378 519266 20614
rect 519502 20378 519586 20614
rect 519822 20378 519854 20614
rect 519234 -5146 519854 20378
rect 521794 43294 522414 58000
rect 521794 43058 521826 43294
rect 522062 43058 522146 43294
rect 522382 43058 522414 43294
rect 521794 23294 522414 43058
rect 521794 23058 521826 23294
rect 522062 23058 522146 23294
rect 522382 23058 522414 23294
rect 521794 3294 522414 23058
rect 521794 3058 521826 3294
rect 522062 3058 522146 3294
rect 522382 3058 522414 3294
rect 521794 -346 522414 3058
rect 521794 -582 521826 -346
rect 522062 -582 522146 -346
rect 522382 -582 522414 -346
rect 521794 -666 522414 -582
rect 521794 -902 521826 -666
rect 522062 -902 522146 -666
rect 522382 -902 522414 -666
rect 521794 -1894 522414 -902
rect 522954 44274 523574 58000
rect 522954 44038 522986 44274
rect 523222 44038 523306 44274
rect 523542 44038 523574 44274
rect 522954 24274 523574 44038
rect 522954 24038 522986 24274
rect 523222 24038 523306 24274
rect 523542 24038 523574 24274
rect 519234 -5382 519266 -5146
rect 519502 -5382 519586 -5146
rect 519822 -5382 519854 -5146
rect 519234 -5466 519854 -5382
rect 519234 -5702 519266 -5466
rect 519502 -5702 519586 -5466
rect 519822 -5702 519854 -5466
rect 519234 -5734 519854 -5702
rect 512954 -6342 512986 -6106
rect 513222 -6342 513306 -6106
rect 513542 -6342 513574 -6106
rect 512954 -6426 513574 -6342
rect 512954 -6662 512986 -6426
rect 513222 -6662 513306 -6426
rect 513542 -6662 513574 -6426
rect 512954 -7654 513574 -6662
rect 522954 -7066 523574 24038
rect 525514 46954 526134 58000
rect 525514 46718 525546 46954
rect 525782 46718 525866 46954
rect 526102 46718 526134 46954
rect 525514 26954 526134 46718
rect 525514 26718 525546 26954
rect 525782 26718 525866 26954
rect 526102 26718 526134 26954
rect 525514 6954 526134 26718
rect 525514 6718 525546 6954
rect 525782 6718 525866 6954
rect 526102 6718 526134 6954
rect 525514 -2266 526134 6718
rect 525514 -2502 525546 -2266
rect 525782 -2502 525866 -2266
rect 526102 -2502 526134 -2266
rect 525514 -2586 526134 -2502
rect 525514 -2822 525546 -2586
rect 525782 -2822 525866 -2586
rect 526102 -2822 526134 -2586
rect 525514 -3814 526134 -2822
rect 529234 50614 529854 58000
rect 529234 50378 529266 50614
rect 529502 50378 529586 50614
rect 529822 50378 529854 50614
rect 529234 30614 529854 50378
rect 529234 30378 529266 30614
rect 529502 30378 529586 30614
rect 529822 30378 529854 30614
rect 529234 10614 529854 30378
rect 529234 10378 529266 10614
rect 529502 10378 529586 10614
rect 529822 10378 529854 10614
rect 529234 -4186 529854 10378
rect 531794 53294 532414 58000
rect 531794 53058 531826 53294
rect 532062 53058 532146 53294
rect 532382 53058 532414 53294
rect 531794 33294 532414 53058
rect 531794 33058 531826 33294
rect 532062 33058 532146 33294
rect 532382 33058 532414 33294
rect 531794 13294 532414 33058
rect 531794 13058 531826 13294
rect 532062 13058 532146 13294
rect 532382 13058 532414 13294
rect 531794 -1306 532414 13058
rect 531794 -1542 531826 -1306
rect 532062 -1542 532146 -1306
rect 532382 -1542 532414 -1306
rect 531794 -1626 532414 -1542
rect 531794 -1862 531826 -1626
rect 532062 -1862 532146 -1626
rect 532382 -1862 532414 -1626
rect 531794 -1894 532414 -1862
rect 532954 54274 533574 58000
rect 532954 54038 532986 54274
rect 533222 54038 533306 54274
rect 533542 54038 533574 54274
rect 532954 34274 533574 54038
rect 532954 34038 532986 34274
rect 533222 34038 533306 34274
rect 533542 34038 533574 34274
rect 532954 14274 533574 34038
rect 532954 14038 532986 14274
rect 533222 14038 533306 14274
rect 533542 14038 533574 14274
rect 529234 -4422 529266 -4186
rect 529502 -4422 529586 -4186
rect 529822 -4422 529854 -4186
rect 529234 -4506 529854 -4422
rect 529234 -4742 529266 -4506
rect 529502 -4742 529586 -4506
rect 529822 -4742 529854 -4506
rect 529234 -5734 529854 -4742
rect 522954 -7302 522986 -7066
rect 523222 -7302 523306 -7066
rect 523542 -7302 523574 -7066
rect 522954 -7386 523574 -7302
rect 522954 -7622 522986 -7386
rect 523222 -7622 523306 -7386
rect 523542 -7622 523574 -7386
rect 522954 -7654 523574 -7622
rect 532954 -6106 533574 14038
rect 535514 56954 536134 58000
rect 535514 56718 535546 56954
rect 535782 56718 535866 56954
rect 536102 56718 536134 56954
rect 535514 36954 536134 56718
rect 535514 36718 535546 36954
rect 535782 36718 535866 36954
rect 536102 36718 536134 36954
rect 535514 16954 536134 36718
rect 535514 16718 535546 16954
rect 535782 16718 535866 16954
rect 536102 16718 536134 16954
rect 535514 -3226 536134 16718
rect 535514 -3462 535546 -3226
rect 535782 -3462 535866 -3226
rect 536102 -3462 536134 -3226
rect 535514 -3546 536134 -3462
rect 535514 -3782 535546 -3546
rect 535782 -3782 535866 -3546
rect 536102 -3782 536134 -3546
rect 535514 -3814 536134 -3782
rect 539234 40614 539854 58000
rect 539234 40378 539266 40614
rect 539502 40378 539586 40614
rect 539822 40378 539854 40614
rect 539234 20614 539854 40378
rect 539234 20378 539266 20614
rect 539502 20378 539586 20614
rect 539822 20378 539854 20614
rect 539234 -5146 539854 20378
rect 541794 43294 542414 58000
rect 541794 43058 541826 43294
rect 542062 43058 542146 43294
rect 542382 43058 542414 43294
rect 541794 23294 542414 43058
rect 541794 23058 541826 23294
rect 542062 23058 542146 23294
rect 542382 23058 542414 23294
rect 541794 3294 542414 23058
rect 541794 3058 541826 3294
rect 542062 3058 542146 3294
rect 542382 3058 542414 3294
rect 541794 -346 542414 3058
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 542954 44274 543574 58000
rect 542954 44038 542986 44274
rect 543222 44038 543306 44274
rect 543542 44038 543574 44274
rect 542954 24274 543574 44038
rect 542954 24038 542986 24274
rect 543222 24038 543306 24274
rect 543542 24038 543574 24274
rect 539234 -5382 539266 -5146
rect 539502 -5382 539586 -5146
rect 539822 -5382 539854 -5146
rect 539234 -5466 539854 -5382
rect 539234 -5702 539266 -5466
rect 539502 -5702 539586 -5466
rect 539822 -5702 539854 -5466
rect 539234 -5734 539854 -5702
rect 532954 -6342 532986 -6106
rect 533222 -6342 533306 -6106
rect 533542 -6342 533574 -6106
rect 532954 -6426 533574 -6342
rect 532954 -6662 532986 -6426
rect 533222 -6662 533306 -6426
rect 533542 -6662 533574 -6426
rect 532954 -7654 533574 -6662
rect 542954 -7066 543574 24038
rect 545514 46954 546134 58000
rect 545514 46718 545546 46954
rect 545782 46718 545866 46954
rect 546102 46718 546134 46954
rect 545514 26954 546134 46718
rect 545514 26718 545546 26954
rect 545782 26718 545866 26954
rect 546102 26718 546134 26954
rect 545514 6954 546134 26718
rect 545514 6718 545546 6954
rect 545782 6718 545866 6954
rect 546102 6718 546134 6954
rect 545514 -2266 546134 6718
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 50614 549854 58000
rect 549234 50378 549266 50614
rect 549502 50378 549586 50614
rect 549822 50378 549854 50614
rect 549234 30614 549854 50378
rect 549234 30378 549266 30614
rect 549502 30378 549586 30614
rect 549822 30378 549854 30614
rect 549234 10614 549854 30378
rect 549234 10378 549266 10614
rect 549502 10378 549586 10614
rect 549822 10378 549854 10614
rect 549234 -4186 549854 10378
rect 551794 53294 552414 58000
rect 551794 53058 551826 53294
rect 552062 53058 552146 53294
rect 552382 53058 552414 53294
rect 551794 33294 552414 53058
rect 551794 33058 551826 33294
rect 552062 33058 552146 33294
rect 552382 33058 552414 33294
rect 551794 13294 552414 33058
rect 551794 13058 551826 13294
rect 552062 13058 552146 13294
rect 552382 13058 552414 13294
rect 551794 -1306 552414 13058
rect 551794 -1542 551826 -1306
rect 552062 -1542 552146 -1306
rect 552382 -1542 552414 -1306
rect 551794 -1626 552414 -1542
rect 551794 -1862 551826 -1626
rect 552062 -1862 552146 -1626
rect 552382 -1862 552414 -1626
rect 551794 -1894 552414 -1862
rect 552954 54274 553574 58000
rect 552954 54038 552986 54274
rect 553222 54038 553306 54274
rect 553542 54038 553574 54274
rect 552954 34274 553574 54038
rect 552954 34038 552986 34274
rect 553222 34038 553306 34274
rect 553542 34038 553574 34274
rect 552954 14274 553574 34038
rect 552954 14038 552986 14274
rect 553222 14038 553306 14274
rect 553542 14038 553574 14274
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 542954 -7302 542986 -7066
rect 543222 -7302 543306 -7066
rect 543542 -7302 543574 -7066
rect 542954 -7386 543574 -7302
rect 542954 -7622 542986 -7386
rect 543222 -7622 543306 -7386
rect 543542 -7622 543574 -7386
rect 542954 -7654 543574 -7622
rect 552954 -6106 553574 14038
rect 555514 56954 556134 58000
rect 555514 56718 555546 56954
rect 555782 56718 555866 56954
rect 556102 56718 556134 56954
rect 555514 36954 556134 56718
rect 555514 36718 555546 36954
rect 555782 36718 555866 36954
rect 556102 36718 556134 36954
rect 555514 16954 556134 36718
rect 555514 16718 555546 16954
rect 555782 16718 555866 16954
rect 556102 16718 556134 16954
rect 555514 -3226 556134 16718
rect 555514 -3462 555546 -3226
rect 555782 -3462 555866 -3226
rect 556102 -3462 556134 -3226
rect 555514 -3546 556134 -3462
rect 555514 -3782 555546 -3546
rect 555782 -3782 555866 -3546
rect 556102 -3782 556134 -3546
rect 555514 -3814 556134 -3782
rect 559234 40614 559854 60378
rect 559234 40378 559266 40614
rect 559502 40378 559586 40614
rect 559822 40378 559854 40614
rect 559234 20614 559854 40378
rect 559234 20378 559266 20614
rect 559502 20378 559586 20614
rect 559822 20378 559854 20614
rect 559234 -5146 559854 20378
rect 561794 704838 562414 705830
rect 561794 704602 561826 704838
rect 562062 704602 562146 704838
rect 562382 704602 562414 704838
rect 561794 704518 562414 704602
rect 561794 704282 561826 704518
rect 562062 704282 562146 704518
rect 562382 704282 562414 704518
rect 561794 683294 562414 704282
rect 561794 683058 561826 683294
rect 562062 683058 562146 683294
rect 562382 683058 562414 683294
rect 561794 663294 562414 683058
rect 561794 663058 561826 663294
rect 562062 663058 562146 663294
rect 562382 663058 562414 663294
rect 561794 643294 562414 663058
rect 561794 643058 561826 643294
rect 562062 643058 562146 643294
rect 562382 643058 562414 643294
rect 561794 623294 562414 643058
rect 561794 623058 561826 623294
rect 562062 623058 562146 623294
rect 562382 623058 562414 623294
rect 561794 603294 562414 623058
rect 561794 603058 561826 603294
rect 562062 603058 562146 603294
rect 562382 603058 562414 603294
rect 561794 583294 562414 603058
rect 561794 583058 561826 583294
rect 562062 583058 562146 583294
rect 562382 583058 562414 583294
rect 561794 563294 562414 583058
rect 561794 563058 561826 563294
rect 562062 563058 562146 563294
rect 562382 563058 562414 563294
rect 561794 543294 562414 563058
rect 561794 543058 561826 543294
rect 562062 543058 562146 543294
rect 562382 543058 562414 543294
rect 561794 523294 562414 543058
rect 561794 523058 561826 523294
rect 562062 523058 562146 523294
rect 562382 523058 562414 523294
rect 561794 503294 562414 523058
rect 561794 503058 561826 503294
rect 562062 503058 562146 503294
rect 562382 503058 562414 503294
rect 561794 483294 562414 503058
rect 561794 483058 561826 483294
rect 562062 483058 562146 483294
rect 562382 483058 562414 483294
rect 561794 463294 562414 483058
rect 561794 463058 561826 463294
rect 562062 463058 562146 463294
rect 562382 463058 562414 463294
rect 561794 443294 562414 463058
rect 561794 443058 561826 443294
rect 562062 443058 562146 443294
rect 562382 443058 562414 443294
rect 561794 423294 562414 443058
rect 561794 423058 561826 423294
rect 562062 423058 562146 423294
rect 562382 423058 562414 423294
rect 561794 403294 562414 423058
rect 561794 403058 561826 403294
rect 562062 403058 562146 403294
rect 562382 403058 562414 403294
rect 561794 383294 562414 403058
rect 561794 383058 561826 383294
rect 562062 383058 562146 383294
rect 562382 383058 562414 383294
rect 561794 363294 562414 383058
rect 561794 363058 561826 363294
rect 562062 363058 562146 363294
rect 562382 363058 562414 363294
rect 561794 343294 562414 363058
rect 561794 343058 561826 343294
rect 562062 343058 562146 343294
rect 562382 343058 562414 343294
rect 561794 323294 562414 343058
rect 561794 323058 561826 323294
rect 562062 323058 562146 323294
rect 562382 323058 562414 323294
rect 561794 303294 562414 323058
rect 561794 303058 561826 303294
rect 562062 303058 562146 303294
rect 562382 303058 562414 303294
rect 561794 283294 562414 303058
rect 561794 283058 561826 283294
rect 562062 283058 562146 283294
rect 562382 283058 562414 283294
rect 561794 263294 562414 283058
rect 561794 263058 561826 263294
rect 562062 263058 562146 263294
rect 562382 263058 562414 263294
rect 561794 243294 562414 263058
rect 561794 243058 561826 243294
rect 562062 243058 562146 243294
rect 562382 243058 562414 243294
rect 561794 223294 562414 243058
rect 561794 223058 561826 223294
rect 562062 223058 562146 223294
rect 562382 223058 562414 223294
rect 561794 203294 562414 223058
rect 561794 203058 561826 203294
rect 562062 203058 562146 203294
rect 562382 203058 562414 203294
rect 561794 183294 562414 203058
rect 561794 183058 561826 183294
rect 562062 183058 562146 183294
rect 562382 183058 562414 183294
rect 561794 163294 562414 183058
rect 561794 163058 561826 163294
rect 562062 163058 562146 163294
rect 562382 163058 562414 163294
rect 561794 143294 562414 163058
rect 561794 143058 561826 143294
rect 562062 143058 562146 143294
rect 562382 143058 562414 143294
rect 561794 123294 562414 143058
rect 561794 123058 561826 123294
rect 562062 123058 562146 123294
rect 562382 123058 562414 123294
rect 561794 103294 562414 123058
rect 561794 103058 561826 103294
rect 562062 103058 562146 103294
rect 562382 103058 562414 103294
rect 561794 83294 562414 103058
rect 561794 83058 561826 83294
rect 562062 83058 562146 83294
rect 562382 83058 562414 83294
rect 561794 63294 562414 83058
rect 561794 63058 561826 63294
rect 562062 63058 562146 63294
rect 562382 63058 562414 63294
rect 561794 43294 562414 63058
rect 561794 43058 561826 43294
rect 562062 43058 562146 43294
rect 562382 43058 562414 43294
rect 561794 23294 562414 43058
rect 561794 23058 561826 23294
rect 562062 23058 562146 23294
rect 562382 23058 562414 23294
rect 561794 3294 562414 23058
rect 561794 3058 561826 3294
rect 562062 3058 562146 3294
rect 562382 3058 562414 3294
rect 561794 -346 562414 3058
rect 561794 -582 561826 -346
rect 562062 -582 562146 -346
rect 562382 -582 562414 -346
rect 561794 -666 562414 -582
rect 561794 -902 561826 -666
rect 562062 -902 562146 -666
rect 562382 -902 562414 -666
rect 561794 -1894 562414 -902
rect 562954 684274 563574 711002
rect 572954 710598 573574 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 572954 710362 572986 710598
rect 573222 710362 573306 710598
rect 573542 710362 573574 710598
rect 572954 710278 573574 710362
rect 572954 710042 572986 710278
rect 573222 710042 573306 710278
rect 573542 710042 573574 710278
rect 569234 708678 569854 709670
rect 569234 708442 569266 708678
rect 569502 708442 569586 708678
rect 569822 708442 569854 708678
rect 569234 708358 569854 708442
rect 569234 708122 569266 708358
rect 569502 708122 569586 708358
rect 569822 708122 569854 708358
rect 562954 684038 562986 684274
rect 563222 684038 563306 684274
rect 563542 684038 563574 684274
rect 562954 664274 563574 684038
rect 562954 664038 562986 664274
rect 563222 664038 563306 664274
rect 563542 664038 563574 664274
rect 562954 644274 563574 664038
rect 562954 644038 562986 644274
rect 563222 644038 563306 644274
rect 563542 644038 563574 644274
rect 562954 624274 563574 644038
rect 562954 624038 562986 624274
rect 563222 624038 563306 624274
rect 563542 624038 563574 624274
rect 562954 604274 563574 624038
rect 562954 604038 562986 604274
rect 563222 604038 563306 604274
rect 563542 604038 563574 604274
rect 562954 584274 563574 604038
rect 562954 584038 562986 584274
rect 563222 584038 563306 584274
rect 563542 584038 563574 584274
rect 562954 564274 563574 584038
rect 562954 564038 562986 564274
rect 563222 564038 563306 564274
rect 563542 564038 563574 564274
rect 562954 544274 563574 564038
rect 562954 544038 562986 544274
rect 563222 544038 563306 544274
rect 563542 544038 563574 544274
rect 562954 524274 563574 544038
rect 562954 524038 562986 524274
rect 563222 524038 563306 524274
rect 563542 524038 563574 524274
rect 562954 504274 563574 524038
rect 562954 504038 562986 504274
rect 563222 504038 563306 504274
rect 563542 504038 563574 504274
rect 562954 484274 563574 504038
rect 562954 484038 562986 484274
rect 563222 484038 563306 484274
rect 563542 484038 563574 484274
rect 562954 464274 563574 484038
rect 562954 464038 562986 464274
rect 563222 464038 563306 464274
rect 563542 464038 563574 464274
rect 562954 444274 563574 464038
rect 562954 444038 562986 444274
rect 563222 444038 563306 444274
rect 563542 444038 563574 444274
rect 562954 424274 563574 444038
rect 562954 424038 562986 424274
rect 563222 424038 563306 424274
rect 563542 424038 563574 424274
rect 562954 404274 563574 424038
rect 562954 404038 562986 404274
rect 563222 404038 563306 404274
rect 563542 404038 563574 404274
rect 562954 384274 563574 404038
rect 562954 384038 562986 384274
rect 563222 384038 563306 384274
rect 563542 384038 563574 384274
rect 562954 364274 563574 384038
rect 562954 364038 562986 364274
rect 563222 364038 563306 364274
rect 563542 364038 563574 364274
rect 562954 344274 563574 364038
rect 562954 344038 562986 344274
rect 563222 344038 563306 344274
rect 563542 344038 563574 344274
rect 562954 324274 563574 344038
rect 562954 324038 562986 324274
rect 563222 324038 563306 324274
rect 563542 324038 563574 324274
rect 562954 304274 563574 324038
rect 562954 304038 562986 304274
rect 563222 304038 563306 304274
rect 563542 304038 563574 304274
rect 562954 284274 563574 304038
rect 562954 284038 562986 284274
rect 563222 284038 563306 284274
rect 563542 284038 563574 284274
rect 562954 264274 563574 284038
rect 562954 264038 562986 264274
rect 563222 264038 563306 264274
rect 563542 264038 563574 264274
rect 562954 244274 563574 264038
rect 562954 244038 562986 244274
rect 563222 244038 563306 244274
rect 563542 244038 563574 244274
rect 562954 224274 563574 244038
rect 562954 224038 562986 224274
rect 563222 224038 563306 224274
rect 563542 224038 563574 224274
rect 562954 204274 563574 224038
rect 562954 204038 562986 204274
rect 563222 204038 563306 204274
rect 563542 204038 563574 204274
rect 562954 184274 563574 204038
rect 562954 184038 562986 184274
rect 563222 184038 563306 184274
rect 563542 184038 563574 184274
rect 562954 164274 563574 184038
rect 562954 164038 562986 164274
rect 563222 164038 563306 164274
rect 563542 164038 563574 164274
rect 562954 144274 563574 164038
rect 562954 144038 562986 144274
rect 563222 144038 563306 144274
rect 563542 144038 563574 144274
rect 562954 124274 563574 144038
rect 562954 124038 562986 124274
rect 563222 124038 563306 124274
rect 563542 124038 563574 124274
rect 562954 104274 563574 124038
rect 562954 104038 562986 104274
rect 563222 104038 563306 104274
rect 563542 104038 563574 104274
rect 562954 84274 563574 104038
rect 562954 84038 562986 84274
rect 563222 84038 563306 84274
rect 563542 84038 563574 84274
rect 562954 64274 563574 84038
rect 562954 64038 562986 64274
rect 563222 64038 563306 64274
rect 563542 64038 563574 64274
rect 562954 44274 563574 64038
rect 562954 44038 562986 44274
rect 563222 44038 563306 44274
rect 563542 44038 563574 44274
rect 562954 24274 563574 44038
rect 562954 24038 562986 24274
rect 563222 24038 563306 24274
rect 563542 24038 563574 24274
rect 559234 -5382 559266 -5146
rect 559502 -5382 559586 -5146
rect 559822 -5382 559854 -5146
rect 559234 -5466 559854 -5382
rect 559234 -5702 559266 -5466
rect 559502 -5702 559586 -5466
rect 559822 -5702 559854 -5466
rect 559234 -5734 559854 -5702
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 562954 -7066 563574 24038
rect 565514 706758 566134 707750
rect 565514 706522 565546 706758
rect 565782 706522 565866 706758
rect 566102 706522 566134 706758
rect 565514 706438 566134 706522
rect 565514 706202 565546 706438
rect 565782 706202 565866 706438
rect 566102 706202 566134 706438
rect 565514 686954 566134 706202
rect 565514 686718 565546 686954
rect 565782 686718 565866 686954
rect 566102 686718 566134 686954
rect 565514 666954 566134 686718
rect 565514 666718 565546 666954
rect 565782 666718 565866 666954
rect 566102 666718 566134 666954
rect 565514 646954 566134 666718
rect 565514 646718 565546 646954
rect 565782 646718 565866 646954
rect 566102 646718 566134 646954
rect 565514 626954 566134 646718
rect 565514 626718 565546 626954
rect 565782 626718 565866 626954
rect 566102 626718 566134 626954
rect 565514 606954 566134 626718
rect 565514 606718 565546 606954
rect 565782 606718 565866 606954
rect 566102 606718 566134 606954
rect 565514 586954 566134 606718
rect 565514 586718 565546 586954
rect 565782 586718 565866 586954
rect 566102 586718 566134 586954
rect 565514 566954 566134 586718
rect 565514 566718 565546 566954
rect 565782 566718 565866 566954
rect 566102 566718 566134 566954
rect 565514 546954 566134 566718
rect 565514 546718 565546 546954
rect 565782 546718 565866 546954
rect 566102 546718 566134 546954
rect 565514 526954 566134 546718
rect 565514 526718 565546 526954
rect 565782 526718 565866 526954
rect 566102 526718 566134 526954
rect 565514 506954 566134 526718
rect 565514 506718 565546 506954
rect 565782 506718 565866 506954
rect 566102 506718 566134 506954
rect 565514 486954 566134 506718
rect 565514 486718 565546 486954
rect 565782 486718 565866 486954
rect 566102 486718 566134 486954
rect 565514 466954 566134 486718
rect 565514 466718 565546 466954
rect 565782 466718 565866 466954
rect 566102 466718 566134 466954
rect 565514 446954 566134 466718
rect 565514 446718 565546 446954
rect 565782 446718 565866 446954
rect 566102 446718 566134 446954
rect 565514 426954 566134 446718
rect 565514 426718 565546 426954
rect 565782 426718 565866 426954
rect 566102 426718 566134 426954
rect 565514 406954 566134 426718
rect 565514 406718 565546 406954
rect 565782 406718 565866 406954
rect 566102 406718 566134 406954
rect 565514 386954 566134 406718
rect 565514 386718 565546 386954
rect 565782 386718 565866 386954
rect 566102 386718 566134 386954
rect 565514 366954 566134 386718
rect 565514 366718 565546 366954
rect 565782 366718 565866 366954
rect 566102 366718 566134 366954
rect 565514 346954 566134 366718
rect 565514 346718 565546 346954
rect 565782 346718 565866 346954
rect 566102 346718 566134 346954
rect 565514 326954 566134 346718
rect 565514 326718 565546 326954
rect 565782 326718 565866 326954
rect 566102 326718 566134 326954
rect 565514 306954 566134 326718
rect 565514 306718 565546 306954
rect 565782 306718 565866 306954
rect 566102 306718 566134 306954
rect 565514 286954 566134 306718
rect 565514 286718 565546 286954
rect 565782 286718 565866 286954
rect 566102 286718 566134 286954
rect 565514 266954 566134 286718
rect 565514 266718 565546 266954
rect 565782 266718 565866 266954
rect 566102 266718 566134 266954
rect 565514 246954 566134 266718
rect 565514 246718 565546 246954
rect 565782 246718 565866 246954
rect 566102 246718 566134 246954
rect 565514 226954 566134 246718
rect 565514 226718 565546 226954
rect 565782 226718 565866 226954
rect 566102 226718 566134 226954
rect 565514 206954 566134 226718
rect 565514 206718 565546 206954
rect 565782 206718 565866 206954
rect 566102 206718 566134 206954
rect 565514 186954 566134 206718
rect 565514 186718 565546 186954
rect 565782 186718 565866 186954
rect 566102 186718 566134 186954
rect 565514 166954 566134 186718
rect 565514 166718 565546 166954
rect 565782 166718 565866 166954
rect 566102 166718 566134 166954
rect 565514 146954 566134 166718
rect 565514 146718 565546 146954
rect 565782 146718 565866 146954
rect 566102 146718 566134 146954
rect 565514 126954 566134 146718
rect 565514 126718 565546 126954
rect 565782 126718 565866 126954
rect 566102 126718 566134 126954
rect 565514 106954 566134 126718
rect 565514 106718 565546 106954
rect 565782 106718 565866 106954
rect 566102 106718 566134 106954
rect 565514 86954 566134 106718
rect 565514 86718 565546 86954
rect 565782 86718 565866 86954
rect 566102 86718 566134 86954
rect 565514 66954 566134 86718
rect 565514 66718 565546 66954
rect 565782 66718 565866 66954
rect 566102 66718 566134 66954
rect 565514 46954 566134 66718
rect 565514 46718 565546 46954
rect 565782 46718 565866 46954
rect 566102 46718 566134 46954
rect 565514 26954 566134 46718
rect 565514 26718 565546 26954
rect 565782 26718 565866 26954
rect 566102 26718 566134 26954
rect 565514 6954 566134 26718
rect 565514 6718 565546 6954
rect 565782 6718 565866 6954
rect 566102 6718 566134 6954
rect 565514 -2266 566134 6718
rect 565514 -2502 565546 -2266
rect 565782 -2502 565866 -2266
rect 566102 -2502 566134 -2266
rect 565514 -2586 566134 -2502
rect 565514 -2822 565546 -2586
rect 565782 -2822 565866 -2586
rect 566102 -2822 566134 -2586
rect 565514 -3814 566134 -2822
rect 569234 690614 569854 708122
rect 569234 690378 569266 690614
rect 569502 690378 569586 690614
rect 569822 690378 569854 690614
rect 569234 670614 569854 690378
rect 569234 670378 569266 670614
rect 569502 670378 569586 670614
rect 569822 670378 569854 670614
rect 569234 650614 569854 670378
rect 569234 650378 569266 650614
rect 569502 650378 569586 650614
rect 569822 650378 569854 650614
rect 569234 630614 569854 650378
rect 569234 630378 569266 630614
rect 569502 630378 569586 630614
rect 569822 630378 569854 630614
rect 569234 610614 569854 630378
rect 569234 610378 569266 610614
rect 569502 610378 569586 610614
rect 569822 610378 569854 610614
rect 569234 590614 569854 610378
rect 569234 590378 569266 590614
rect 569502 590378 569586 590614
rect 569822 590378 569854 590614
rect 569234 570614 569854 590378
rect 569234 570378 569266 570614
rect 569502 570378 569586 570614
rect 569822 570378 569854 570614
rect 569234 550614 569854 570378
rect 569234 550378 569266 550614
rect 569502 550378 569586 550614
rect 569822 550378 569854 550614
rect 569234 530614 569854 550378
rect 569234 530378 569266 530614
rect 569502 530378 569586 530614
rect 569822 530378 569854 530614
rect 569234 510614 569854 530378
rect 569234 510378 569266 510614
rect 569502 510378 569586 510614
rect 569822 510378 569854 510614
rect 569234 490614 569854 510378
rect 569234 490378 569266 490614
rect 569502 490378 569586 490614
rect 569822 490378 569854 490614
rect 569234 470614 569854 490378
rect 569234 470378 569266 470614
rect 569502 470378 569586 470614
rect 569822 470378 569854 470614
rect 569234 450614 569854 470378
rect 569234 450378 569266 450614
rect 569502 450378 569586 450614
rect 569822 450378 569854 450614
rect 569234 430614 569854 450378
rect 569234 430378 569266 430614
rect 569502 430378 569586 430614
rect 569822 430378 569854 430614
rect 569234 410614 569854 430378
rect 569234 410378 569266 410614
rect 569502 410378 569586 410614
rect 569822 410378 569854 410614
rect 569234 390614 569854 410378
rect 569234 390378 569266 390614
rect 569502 390378 569586 390614
rect 569822 390378 569854 390614
rect 569234 370614 569854 390378
rect 569234 370378 569266 370614
rect 569502 370378 569586 370614
rect 569822 370378 569854 370614
rect 569234 350614 569854 370378
rect 569234 350378 569266 350614
rect 569502 350378 569586 350614
rect 569822 350378 569854 350614
rect 569234 330614 569854 350378
rect 569234 330378 569266 330614
rect 569502 330378 569586 330614
rect 569822 330378 569854 330614
rect 569234 310614 569854 330378
rect 569234 310378 569266 310614
rect 569502 310378 569586 310614
rect 569822 310378 569854 310614
rect 569234 290614 569854 310378
rect 569234 290378 569266 290614
rect 569502 290378 569586 290614
rect 569822 290378 569854 290614
rect 569234 270614 569854 290378
rect 569234 270378 569266 270614
rect 569502 270378 569586 270614
rect 569822 270378 569854 270614
rect 569234 250614 569854 270378
rect 569234 250378 569266 250614
rect 569502 250378 569586 250614
rect 569822 250378 569854 250614
rect 569234 230614 569854 250378
rect 569234 230378 569266 230614
rect 569502 230378 569586 230614
rect 569822 230378 569854 230614
rect 569234 210614 569854 230378
rect 569234 210378 569266 210614
rect 569502 210378 569586 210614
rect 569822 210378 569854 210614
rect 569234 190614 569854 210378
rect 569234 190378 569266 190614
rect 569502 190378 569586 190614
rect 569822 190378 569854 190614
rect 569234 170614 569854 190378
rect 569234 170378 569266 170614
rect 569502 170378 569586 170614
rect 569822 170378 569854 170614
rect 569234 150614 569854 170378
rect 569234 150378 569266 150614
rect 569502 150378 569586 150614
rect 569822 150378 569854 150614
rect 569234 130614 569854 150378
rect 569234 130378 569266 130614
rect 569502 130378 569586 130614
rect 569822 130378 569854 130614
rect 569234 110614 569854 130378
rect 569234 110378 569266 110614
rect 569502 110378 569586 110614
rect 569822 110378 569854 110614
rect 569234 90614 569854 110378
rect 569234 90378 569266 90614
rect 569502 90378 569586 90614
rect 569822 90378 569854 90614
rect 569234 70614 569854 90378
rect 569234 70378 569266 70614
rect 569502 70378 569586 70614
rect 569822 70378 569854 70614
rect 569234 50614 569854 70378
rect 569234 50378 569266 50614
rect 569502 50378 569586 50614
rect 569822 50378 569854 50614
rect 569234 30614 569854 50378
rect 569234 30378 569266 30614
rect 569502 30378 569586 30614
rect 569822 30378 569854 30614
rect 569234 10614 569854 30378
rect 569234 10378 569266 10614
rect 569502 10378 569586 10614
rect 569822 10378 569854 10614
rect 569234 -4186 569854 10378
rect 571794 705798 572414 705830
rect 571794 705562 571826 705798
rect 572062 705562 572146 705798
rect 572382 705562 572414 705798
rect 571794 705478 572414 705562
rect 571794 705242 571826 705478
rect 572062 705242 572146 705478
rect 572382 705242 572414 705478
rect 571794 693294 572414 705242
rect 571794 693058 571826 693294
rect 572062 693058 572146 693294
rect 572382 693058 572414 693294
rect 571794 673294 572414 693058
rect 571794 673058 571826 673294
rect 572062 673058 572146 673294
rect 572382 673058 572414 673294
rect 571794 653294 572414 673058
rect 571794 653058 571826 653294
rect 572062 653058 572146 653294
rect 572382 653058 572414 653294
rect 571794 633294 572414 653058
rect 571794 633058 571826 633294
rect 572062 633058 572146 633294
rect 572382 633058 572414 633294
rect 571794 613294 572414 633058
rect 571794 613058 571826 613294
rect 572062 613058 572146 613294
rect 572382 613058 572414 613294
rect 571794 593294 572414 613058
rect 571794 593058 571826 593294
rect 572062 593058 572146 593294
rect 572382 593058 572414 593294
rect 571794 573294 572414 593058
rect 571794 573058 571826 573294
rect 572062 573058 572146 573294
rect 572382 573058 572414 573294
rect 571794 553294 572414 573058
rect 571794 553058 571826 553294
rect 572062 553058 572146 553294
rect 572382 553058 572414 553294
rect 571794 533294 572414 553058
rect 571794 533058 571826 533294
rect 572062 533058 572146 533294
rect 572382 533058 572414 533294
rect 571794 513294 572414 533058
rect 571794 513058 571826 513294
rect 572062 513058 572146 513294
rect 572382 513058 572414 513294
rect 571794 493294 572414 513058
rect 571794 493058 571826 493294
rect 572062 493058 572146 493294
rect 572382 493058 572414 493294
rect 571794 473294 572414 493058
rect 571794 473058 571826 473294
rect 572062 473058 572146 473294
rect 572382 473058 572414 473294
rect 571794 453294 572414 473058
rect 571794 453058 571826 453294
rect 572062 453058 572146 453294
rect 572382 453058 572414 453294
rect 571794 433294 572414 453058
rect 571794 433058 571826 433294
rect 572062 433058 572146 433294
rect 572382 433058 572414 433294
rect 571794 413294 572414 433058
rect 571794 413058 571826 413294
rect 572062 413058 572146 413294
rect 572382 413058 572414 413294
rect 571794 393294 572414 413058
rect 571794 393058 571826 393294
rect 572062 393058 572146 393294
rect 572382 393058 572414 393294
rect 571794 373294 572414 393058
rect 571794 373058 571826 373294
rect 572062 373058 572146 373294
rect 572382 373058 572414 373294
rect 571794 353294 572414 373058
rect 571794 353058 571826 353294
rect 572062 353058 572146 353294
rect 572382 353058 572414 353294
rect 571794 333294 572414 353058
rect 571794 333058 571826 333294
rect 572062 333058 572146 333294
rect 572382 333058 572414 333294
rect 571794 313294 572414 333058
rect 571794 313058 571826 313294
rect 572062 313058 572146 313294
rect 572382 313058 572414 313294
rect 571794 293294 572414 313058
rect 571794 293058 571826 293294
rect 572062 293058 572146 293294
rect 572382 293058 572414 293294
rect 571794 273294 572414 293058
rect 571794 273058 571826 273294
rect 572062 273058 572146 273294
rect 572382 273058 572414 273294
rect 571794 253294 572414 273058
rect 571794 253058 571826 253294
rect 572062 253058 572146 253294
rect 572382 253058 572414 253294
rect 571794 233294 572414 253058
rect 571794 233058 571826 233294
rect 572062 233058 572146 233294
rect 572382 233058 572414 233294
rect 571794 213294 572414 233058
rect 571794 213058 571826 213294
rect 572062 213058 572146 213294
rect 572382 213058 572414 213294
rect 571794 193294 572414 213058
rect 571794 193058 571826 193294
rect 572062 193058 572146 193294
rect 572382 193058 572414 193294
rect 571794 173294 572414 193058
rect 571794 173058 571826 173294
rect 572062 173058 572146 173294
rect 572382 173058 572414 173294
rect 571794 153294 572414 173058
rect 571794 153058 571826 153294
rect 572062 153058 572146 153294
rect 572382 153058 572414 153294
rect 571794 133294 572414 153058
rect 571794 133058 571826 133294
rect 572062 133058 572146 133294
rect 572382 133058 572414 133294
rect 571794 113294 572414 133058
rect 571794 113058 571826 113294
rect 572062 113058 572146 113294
rect 572382 113058 572414 113294
rect 571794 93294 572414 113058
rect 571794 93058 571826 93294
rect 572062 93058 572146 93294
rect 572382 93058 572414 93294
rect 571794 73294 572414 93058
rect 571794 73058 571826 73294
rect 572062 73058 572146 73294
rect 572382 73058 572414 73294
rect 571794 53294 572414 73058
rect 571794 53058 571826 53294
rect 572062 53058 572146 53294
rect 572382 53058 572414 53294
rect 571794 33294 572414 53058
rect 571794 33058 571826 33294
rect 572062 33058 572146 33294
rect 572382 33058 572414 33294
rect 571794 13294 572414 33058
rect 571794 13058 571826 13294
rect 572062 13058 572146 13294
rect 572382 13058 572414 13294
rect 571794 -1306 572414 13058
rect 571794 -1542 571826 -1306
rect 572062 -1542 572146 -1306
rect 572382 -1542 572414 -1306
rect 571794 -1626 572414 -1542
rect 571794 -1862 571826 -1626
rect 572062 -1862 572146 -1626
rect 572382 -1862 572414 -1626
rect 571794 -1894 572414 -1862
rect 572954 694274 573574 710042
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 579234 709638 579854 709670
rect 579234 709402 579266 709638
rect 579502 709402 579586 709638
rect 579822 709402 579854 709638
rect 579234 709318 579854 709402
rect 579234 709082 579266 709318
rect 579502 709082 579586 709318
rect 579822 709082 579854 709318
rect 572954 694038 572986 694274
rect 573222 694038 573306 694274
rect 573542 694038 573574 694274
rect 572954 674274 573574 694038
rect 572954 674038 572986 674274
rect 573222 674038 573306 674274
rect 573542 674038 573574 674274
rect 572954 654274 573574 674038
rect 572954 654038 572986 654274
rect 573222 654038 573306 654274
rect 573542 654038 573574 654274
rect 572954 634274 573574 654038
rect 572954 634038 572986 634274
rect 573222 634038 573306 634274
rect 573542 634038 573574 634274
rect 572954 614274 573574 634038
rect 572954 614038 572986 614274
rect 573222 614038 573306 614274
rect 573542 614038 573574 614274
rect 572954 594274 573574 614038
rect 572954 594038 572986 594274
rect 573222 594038 573306 594274
rect 573542 594038 573574 594274
rect 572954 574274 573574 594038
rect 572954 574038 572986 574274
rect 573222 574038 573306 574274
rect 573542 574038 573574 574274
rect 572954 554274 573574 574038
rect 572954 554038 572986 554274
rect 573222 554038 573306 554274
rect 573542 554038 573574 554274
rect 572954 534274 573574 554038
rect 572954 534038 572986 534274
rect 573222 534038 573306 534274
rect 573542 534038 573574 534274
rect 572954 514274 573574 534038
rect 572954 514038 572986 514274
rect 573222 514038 573306 514274
rect 573542 514038 573574 514274
rect 572954 494274 573574 514038
rect 572954 494038 572986 494274
rect 573222 494038 573306 494274
rect 573542 494038 573574 494274
rect 572954 474274 573574 494038
rect 572954 474038 572986 474274
rect 573222 474038 573306 474274
rect 573542 474038 573574 474274
rect 572954 454274 573574 474038
rect 572954 454038 572986 454274
rect 573222 454038 573306 454274
rect 573542 454038 573574 454274
rect 572954 434274 573574 454038
rect 572954 434038 572986 434274
rect 573222 434038 573306 434274
rect 573542 434038 573574 434274
rect 572954 414274 573574 434038
rect 572954 414038 572986 414274
rect 573222 414038 573306 414274
rect 573542 414038 573574 414274
rect 572954 394274 573574 414038
rect 572954 394038 572986 394274
rect 573222 394038 573306 394274
rect 573542 394038 573574 394274
rect 572954 374274 573574 394038
rect 572954 374038 572986 374274
rect 573222 374038 573306 374274
rect 573542 374038 573574 374274
rect 572954 354274 573574 374038
rect 572954 354038 572986 354274
rect 573222 354038 573306 354274
rect 573542 354038 573574 354274
rect 572954 334274 573574 354038
rect 572954 334038 572986 334274
rect 573222 334038 573306 334274
rect 573542 334038 573574 334274
rect 572954 314274 573574 334038
rect 572954 314038 572986 314274
rect 573222 314038 573306 314274
rect 573542 314038 573574 314274
rect 572954 294274 573574 314038
rect 572954 294038 572986 294274
rect 573222 294038 573306 294274
rect 573542 294038 573574 294274
rect 572954 274274 573574 294038
rect 572954 274038 572986 274274
rect 573222 274038 573306 274274
rect 573542 274038 573574 274274
rect 572954 254274 573574 274038
rect 572954 254038 572986 254274
rect 573222 254038 573306 254274
rect 573542 254038 573574 254274
rect 572954 234274 573574 254038
rect 572954 234038 572986 234274
rect 573222 234038 573306 234274
rect 573542 234038 573574 234274
rect 572954 214274 573574 234038
rect 572954 214038 572986 214274
rect 573222 214038 573306 214274
rect 573542 214038 573574 214274
rect 572954 194274 573574 214038
rect 572954 194038 572986 194274
rect 573222 194038 573306 194274
rect 573542 194038 573574 194274
rect 572954 174274 573574 194038
rect 572954 174038 572986 174274
rect 573222 174038 573306 174274
rect 573542 174038 573574 174274
rect 572954 154274 573574 174038
rect 572954 154038 572986 154274
rect 573222 154038 573306 154274
rect 573542 154038 573574 154274
rect 572954 134274 573574 154038
rect 572954 134038 572986 134274
rect 573222 134038 573306 134274
rect 573542 134038 573574 134274
rect 572954 114274 573574 134038
rect 572954 114038 572986 114274
rect 573222 114038 573306 114274
rect 573542 114038 573574 114274
rect 572954 94274 573574 114038
rect 572954 94038 572986 94274
rect 573222 94038 573306 94274
rect 573542 94038 573574 94274
rect 572954 74274 573574 94038
rect 572954 74038 572986 74274
rect 573222 74038 573306 74274
rect 573542 74038 573574 74274
rect 572954 54274 573574 74038
rect 572954 54038 572986 54274
rect 573222 54038 573306 54274
rect 573542 54038 573574 54274
rect 572954 34274 573574 54038
rect 572954 34038 572986 34274
rect 573222 34038 573306 34274
rect 573542 34038 573574 34274
rect 572954 14274 573574 34038
rect 572954 14038 572986 14274
rect 573222 14038 573306 14274
rect 573542 14038 573574 14274
rect 569234 -4422 569266 -4186
rect 569502 -4422 569586 -4186
rect 569822 -4422 569854 -4186
rect 569234 -4506 569854 -4422
rect 569234 -4742 569266 -4506
rect 569502 -4742 569586 -4506
rect 569822 -4742 569854 -4506
rect 569234 -5734 569854 -4742
rect 562954 -7302 562986 -7066
rect 563222 -7302 563306 -7066
rect 563542 -7302 563574 -7066
rect 562954 -7386 563574 -7302
rect 562954 -7622 562986 -7386
rect 563222 -7622 563306 -7386
rect 563542 -7622 563574 -7386
rect 562954 -7654 563574 -7622
rect 572954 -6106 573574 14038
rect 575514 707718 576134 707750
rect 575514 707482 575546 707718
rect 575782 707482 575866 707718
rect 576102 707482 576134 707718
rect 575514 707398 576134 707482
rect 575514 707162 575546 707398
rect 575782 707162 575866 707398
rect 576102 707162 576134 707398
rect 575514 696954 576134 707162
rect 575514 696718 575546 696954
rect 575782 696718 575866 696954
rect 576102 696718 576134 696954
rect 575514 676954 576134 696718
rect 575514 676718 575546 676954
rect 575782 676718 575866 676954
rect 576102 676718 576134 676954
rect 575514 656954 576134 676718
rect 575514 656718 575546 656954
rect 575782 656718 575866 656954
rect 576102 656718 576134 656954
rect 575514 636954 576134 656718
rect 575514 636718 575546 636954
rect 575782 636718 575866 636954
rect 576102 636718 576134 636954
rect 575514 616954 576134 636718
rect 575514 616718 575546 616954
rect 575782 616718 575866 616954
rect 576102 616718 576134 616954
rect 575514 596954 576134 616718
rect 575514 596718 575546 596954
rect 575782 596718 575866 596954
rect 576102 596718 576134 596954
rect 575514 576954 576134 596718
rect 575514 576718 575546 576954
rect 575782 576718 575866 576954
rect 576102 576718 576134 576954
rect 575514 556954 576134 576718
rect 575514 556718 575546 556954
rect 575782 556718 575866 556954
rect 576102 556718 576134 556954
rect 575514 536954 576134 556718
rect 575514 536718 575546 536954
rect 575782 536718 575866 536954
rect 576102 536718 576134 536954
rect 575514 516954 576134 536718
rect 575514 516718 575546 516954
rect 575782 516718 575866 516954
rect 576102 516718 576134 516954
rect 575514 496954 576134 516718
rect 575514 496718 575546 496954
rect 575782 496718 575866 496954
rect 576102 496718 576134 496954
rect 575514 476954 576134 496718
rect 575514 476718 575546 476954
rect 575782 476718 575866 476954
rect 576102 476718 576134 476954
rect 575514 456954 576134 476718
rect 575514 456718 575546 456954
rect 575782 456718 575866 456954
rect 576102 456718 576134 456954
rect 575514 436954 576134 456718
rect 575514 436718 575546 436954
rect 575782 436718 575866 436954
rect 576102 436718 576134 436954
rect 575514 416954 576134 436718
rect 575514 416718 575546 416954
rect 575782 416718 575866 416954
rect 576102 416718 576134 416954
rect 575514 396954 576134 416718
rect 575514 396718 575546 396954
rect 575782 396718 575866 396954
rect 576102 396718 576134 396954
rect 575514 376954 576134 396718
rect 575514 376718 575546 376954
rect 575782 376718 575866 376954
rect 576102 376718 576134 376954
rect 575514 356954 576134 376718
rect 575514 356718 575546 356954
rect 575782 356718 575866 356954
rect 576102 356718 576134 356954
rect 575514 336954 576134 356718
rect 575514 336718 575546 336954
rect 575782 336718 575866 336954
rect 576102 336718 576134 336954
rect 575514 316954 576134 336718
rect 575514 316718 575546 316954
rect 575782 316718 575866 316954
rect 576102 316718 576134 316954
rect 575514 296954 576134 316718
rect 575514 296718 575546 296954
rect 575782 296718 575866 296954
rect 576102 296718 576134 296954
rect 575514 276954 576134 296718
rect 575514 276718 575546 276954
rect 575782 276718 575866 276954
rect 576102 276718 576134 276954
rect 575514 256954 576134 276718
rect 575514 256718 575546 256954
rect 575782 256718 575866 256954
rect 576102 256718 576134 256954
rect 575514 236954 576134 256718
rect 575514 236718 575546 236954
rect 575782 236718 575866 236954
rect 576102 236718 576134 236954
rect 575514 216954 576134 236718
rect 575514 216718 575546 216954
rect 575782 216718 575866 216954
rect 576102 216718 576134 216954
rect 575514 196954 576134 216718
rect 575514 196718 575546 196954
rect 575782 196718 575866 196954
rect 576102 196718 576134 196954
rect 575514 176954 576134 196718
rect 575514 176718 575546 176954
rect 575782 176718 575866 176954
rect 576102 176718 576134 176954
rect 575514 156954 576134 176718
rect 575514 156718 575546 156954
rect 575782 156718 575866 156954
rect 576102 156718 576134 156954
rect 575514 136954 576134 156718
rect 575514 136718 575546 136954
rect 575782 136718 575866 136954
rect 576102 136718 576134 136954
rect 575514 116954 576134 136718
rect 575514 116718 575546 116954
rect 575782 116718 575866 116954
rect 576102 116718 576134 116954
rect 575514 96954 576134 116718
rect 575514 96718 575546 96954
rect 575782 96718 575866 96954
rect 576102 96718 576134 96954
rect 575514 76954 576134 96718
rect 575514 76718 575546 76954
rect 575782 76718 575866 76954
rect 576102 76718 576134 76954
rect 575514 56954 576134 76718
rect 575514 56718 575546 56954
rect 575782 56718 575866 56954
rect 576102 56718 576134 56954
rect 575514 36954 576134 56718
rect 575514 36718 575546 36954
rect 575782 36718 575866 36954
rect 576102 36718 576134 36954
rect 575514 16954 576134 36718
rect 575514 16718 575546 16954
rect 575782 16718 575866 16954
rect 576102 16718 576134 16954
rect 575514 -3226 576134 16718
rect 575514 -3462 575546 -3226
rect 575782 -3462 575866 -3226
rect 576102 -3462 576134 -3226
rect 575514 -3546 576134 -3462
rect 575514 -3782 575546 -3546
rect 575782 -3782 575866 -3546
rect 576102 -3782 576134 -3546
rect 575514 -3814 576134 -3782
rect 579234 700614 579854 709082
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 579234 700378 579266 700614
rect 579502 700378 579586 700614
rect 579822 700378 579854 700614
rect 579234 680614 579854 700378
rect 579234 680378 579266 680614
rect 579502 680378 579586 680614
rect 579822 680378 579854 680614
rect 579234 660614 579854 680378
rect 579234 660378 579266 660614
rect 579502 660378 579586 660614
rect 579822 660378 579854 660614
rect 579234 640614 579854 660378
rect 579234 640378 579266 640614
rect 579502 640378 579586 640614
rect 579822 640378 579854 640614
rect 579234 620614 579854 640378
rect 579234 620378 579266 620614
rect 579502 620378 579586 620614
rect 579822 620378 579854 620614
rect 579234 600614 579854 620378
rect 579234 600378 579266 600614
rect 579502 600378 579586 600614
rect 579822 600378 579854 600614
rect 579234 580614 579854 600378
rect 579234 580378 579266 580614
rect 579502 580378 579586 580614
rect 579822 580378 579854 580614
rect 579234 560614 579854 580378
rect 579234 560378 579266 560614
rect 579502 560378 579586 560614
rect 579822 560378 579854 560614
rect 579234 540614 579854 560378
rect 579234 540378 579266 540614
rect 579502 540378 579586 540614
rect 579822 540378 579854 540614
rect 579234 520614 579854 540378
rect 579234 520378 579266 520614
rect 579502 520378 579586 520614
rect 579822 520378 579854 520614
rect 579234 500614 579854 520378
rect 579234 500378 579266 500614
rect 579502 500378 579586 500614
rect 579822 500378 579854 500614
rect 579234 480614 579854 500378
rect 579234 480378 579266 480614
rect 579502 480378 579586 480614
rect 579822 480378 579854 480614
rect 579234 460614 579854 480378
rect 579234 460378 579266 460614
rect 579502 460378 579586 460614
rect 579822 460378 579854 460614
rect 579234 440614 579854 460378
rect 579234 440378 579266 440614
rect 579502 440378 579586 440614
rect 579822 440378 579854 440614
rect 579234 420614 579854 440378
rect 579234 420378 579266 420614
rect 579502 420378 579586 420614
rect 579822 420378 579854 420614
rect 579234 400614 579854 420378
rect 579234 400378 579266 400614
rect 579502 400378 579586 400614
rect 579822 400378 579854 400614
rect 579234 380614 579854 400378
rect 579234 380378 579266 380614
rect 579502 380378 579586 380614
rect 579822 380378 579854 380614
rect 579234 360614 579854 380378
rect 579234 360378 579266 360614
rect 579502 360378 579586 360614
rect 579822 360378 579854 360614
rect 579234 340614 579854 360378
rect 579234 340378 579266 340614
rect 579502 340378 579586 340614
rect 579822 340378 579854 340614
rect 579234 320614 579854 340378
rect 579234 320378 579266 320614
rect 579502 320378 579586 320614
rect 579822 320378 579854 320614
rect 579234 300614 579854 320378
rect 579234 300378 579266 300614
rect 579502 300378 579586 300614
rect 579822 300378 579854 300614
rect 579234 280614 579854 300378
rect 579234 280378 579266 280614
rect 579502 280378 579586 280614
rect 579822 280378 579854 280614
rect 579234 260614 579854 280378
rect 579234 260378 579266 260614
rect 579502 260378 579586 260614
rect 579822 260378 579854 260614
rect 579234 240614 579854 260378
rect 579234 240378 579266 240614
rect 579502 240378 579586 240614
rect 579822 240378 579854 240614
rect 579234 220614 579854 240378
rect 579234 220378 579266 220614
rect 579502 220378 579586 220614
rect 579822 220378 579854 220614
rect 579234 200614 579854 220378
rect 579234 200378 579266 200614
rect 579502 200378 579586 200614
rect 579822 200378 579854 200614
rect 579234 180614 579854 200378
rect 579234 180378 579266 180614
rect 579502 180378 579586 180614
rect 579822 180378 579854 180614
rect 579234 160614 579854 180378
rect 579234 160378 579266 160614
rect 579502 160378 579586 160614
rect 579822 160378 579854 160614
rect 579234 140614 579854 160378
rect 579234 140378 579266 140614
rect 579502 140378 579586 140614
rect 579822 140378 579854 140614
rect 579234 120614 579854 140378
rect 579234 120378 579266 120614
rect 579502 120378 579586 120614
rect 579822 120378 579854 120614
rect 579234 100614 579854 120378
rect 579234 100378 579266 100614
rect 579502 100378 579586 100614
rect 579822 100378 579854 100614
rect 579234 80614 579854 100378
rect 579234 80378 579266 80614
rect 579502 80378 579586 80614
rect 579822 80378 579854 80614
rect 579234 60614 579854 80378
rect 579234 60378 579266 60614
rect 579502 60378 579586 60614
rect 579822 60378 579854 60614
rect 579234 40614 579854 60378
rect 579234 40378 579266 40614
rect 579502 40378 579586 40614
rect 579822 40378 579854 40614
rect 579234 20614 579854 40378
rect 579234 20378 579266 20614
rect 579502 20378 579586 20614
rect 579822 20378 579854 20614
rect 579234 -5146 579854 20378
rect 581794 704838 582414 705830
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581794 704602 581826 704838
rect 582062 704602 582146 704838
rect 582382 704602 582414 704838
rect 581794 704518 582414 704602
rect 581794 704282 581826 704518
rect 582062 704282 582146 704518
rect 582382 704282 582414 704518
rect 581794 683294 582414 704282
rect 581794 683058 581826 683294
rect 582062 683058 582146 683294
rect 582382 683058 582414 683294
rect 581794 663294 582414 683058
rect 581794 663058 581826 663294
rect 582062 663058 582146 663294
rect 582382 663058 582414 663294
rect 581794 643294 582414 663058
rect 581794 643058 581826 643294
rect 582062 643058 582146 643294
rect 582382 643058 582414 643294
rect 581794 623294 582414 643058
rect 581794 623058 581826 623294
rect 582062 623058 582146 623294
rect 582382 623058 582414 623294
rect 581794 603294 582414 623058
rect 581794 603058 581826 603294
rect 582062 603058 582146 603294
rect 582382 603058 582414 603294
rect 581794 583294 582414 603058
rect 581794 583058 581826 583294
rect 582062 583058 582146 583294
rect 582382 583058 582414 583294
rect 581794 563294 582414 583058
rect 581794 563058 581826 563294
rect 582062 563058 582146 563294
rect 582382 563058 582414 563294
rect 581794 543294 582414 563058
rect 581794 543058 581826 543294
rect 582062 543058 582146 543294
rect 582382 543058 582414 543294
rect 581794 523294 582414 543058
rect 581794 523058 581826 523294
rect 582062 523058 582146 523294
rect 582382 523058 582414 523294
rect 581794 503294 582414 523058
rect 581794 503058 581826 503294
rect 582062 503058 582146 503294
rect 582382 503058 582414 503294
rect 581794 483294 582414 503058
rect 581794 483058 581826 483294
rect 582062 483058 582146 483294
rect 582382 483058 582414 483294
rect 581794 463294 582414 483058
rect 581794 463058 581826 463294
rect 582062 463058 582146 463294
rect 582382 463058 582414 463294
rect 581794 443294 582414 463058
rect 581794 443058 581826 443294
rect 582062 443058 582146 443294
rect 582382 443058 582414 443294
rect 581794 423294 582414 443058
rect 581794 423058 581826 423294
rect 582062 423058 582146 423294
rect 582382 423058 582414 423294
rect 581794 403294 582414 423058
rect 581794 403058 581826 403294
rect 582062 403058 582146 403294
rect 582382 403058 582414 403294
rect 581794 383294 582414 403058
rect 581794 383058 581826 383294
rect 582062 383058 582146 383294
rect 582382 383058 582414 383294
rect 581794 363294 582414 383058
rect 581794 363058 581826 363294
rect 582062 363058 582146 363294
rect 582382 363058 582414 363294
rect 581794 343294 582414 363058
rect 581794 343058 581826 343294
rect 582062 343058 582146 343294
rect 582382 343058 582414 343294
rect 581794 323294 582414 343058
rect 581794 323058 581826 323294
rect 582062 323058 582146 323294
rect 582382 323058 582414 323294
rect 581794 303294 582414 323058
rect 581794 303058 581826 303294
rect 582062 303058 582146 303294
rect 582382 303058 582414 303294
rect 581794 283294 582414 303058
rect 581794 283058 581826 283294
rect 582062 283058 582146 283294
rect 582382 283058 582414 283294
rect 581794 263294 582414 283058
rect 581794 263058 581826 263294
rect 582062 263058 582146 263294
rect 582382 263058 582414 263294
rect 581794 243294 582414 263058
rect 581794 243058 581826 243294
rect 582062 243058 582146 243294
rect 582382 243058 582414 243294
rect 581794 223294 582414 243058
rect 581794 223058 581826 223294
rect 582062 223058 582146 223294
rect 582382 223058 582414 223294
rect 581794 203294 582414 223058
rect 581794 203058 581826 203294
rect 582062 203058 582146 203294
rect 582382 203058 582414 203294
rect 581794 183294 582414 203058
rect 581794 183058 581826 183294
rect 582062 183058 582146 183294
rect 582382 183058 582414 183294
rect 581794 163294 582414 183058
rect 581794 163058 581826 163294
rect 582062 163058 582146 163294
rect 582382 163058 582414 163294
rect 581794 143294 582414 163058
rect 581794 143058 581826 143294
rect 582062 143058 582146 143294
rect 582382 143058 582414 143294
rect 581794 123294 582414 143058
rect 581794 123058 581826 123294
rect 582062 123058 582146 123294
rect 582382 123058 582414 123294
rect 581794 103294 582414 123058
rect 581794 103058 581826 103294
rect 582062 103058 582146 103294
rect 582382 103058 582414 103294
rect 581794 83294 582414 103058
rect 581794 83058 581826 83294
rect 582062 83058 582146 83294
rect 582382 83058 582414 83294
rect 581794 63294 582414 83058
rect 581794 63058 581826 63294
rect 582062 63058 582146 63294
rect 582382 63058 582414 63294
rect 581794 43294 582414 63058
rect 581794 43058 581826 43294
rect 582062 43058 582146 43294
rect 582382 43058 582414 43294
rect 581794 23294 582414 43058
rect 581794 23058 581826 23294
rect 582062 23058 582146 23294
rect 582382 23058 582414 23294
rect 581794 3294 582414 23058
rect 581794 3058 581826 3294
rect 582062 3058 582146 3294
rect 582382 3058 582414 3294
rect 581794 -346 582414 3058
rect 581794 -582 581826 -346
rect 582062 -582 582146 -346
rect 582382 -582 582414 -346
rect 581794 -666 582414 -582
rect 581794 -902 581826 -666
rect 582062 -902 582146 -666
rect 582382 -902 582414 -666
rect 581794 -1894 582414 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 683294 585930 704282
rect 585310 683058 585342 683294
rect 585578 683058 585662 683294
rect 585898 683058 585930 683294
rect 585310 663294 585930 683058
rect 585310 663058 585342 663294
rect 585578 663058 585662 663294
rect 585898 663058 585930 663294
rect 585310 643294 585930 663058
rect 585310 643058 585342 643294
rect 585578 643058 585662 643294
rect 585898 643058 585930 643294
rect 585310 623294 585930 643058
rect 585310 623058 585342 623294
rect 585578 623058 585662 623294
rect 585898 623058 585930 623294
rect 585310 603294 585930 623058
rect 585310 603058 585342 603294
rect 585578 603058 585662 603294
rect 585898 603058 585930 603294
rect 585310 583294 585930 603058
rect 585310 583058 585342 583294
rect 585578 583058 585662 583294
rect 585898 583058 585930 583294
rect 585310 563294 585930 583058
rect 585310 563058 585342 563294
rect 585578 563058 585662 563294
rect 585898 563058 585930 563294
rect 585310 543294 585930 563058
rect 585310 543058 585342 543294
rect 585578 543058 585662 543294
rect 585898 543058 585930 543294
rect 585310 523294 585930 543058
rect 585310 523058 585342 523294
rect 585578 523058 585662 523294
rect 585898 523058 585930 523294
rect 585310 503294 585930 523058
rect 585310 503058 585342 503294
rect 585578 503058 585662 503294
rect 585898 503058 585930 503294
rect 585310 483294 585930 503058
rect 585310 483058 585342 483294
rect 585578 483058 585662 483294
rect 585898 483058 585930 483294
rect 585310 463294 585930 483058
rect 585310 463058 585342 463294
rect 585578 463058 585662 463294
rect 585898 463058 585930 463294
rect 585310 443294 585930 463058
rect 585310 443058 585342 443294
rect 585578 443058 585662 443294
rect 585898 443058 585930 443294
rect 585310 423294 585930 443058
rect 585310 423058 585342 423294
rect 585578 423058 585662 423294
rect 585898 423058 585930 423294
rect 585310 403294 585930 423058
rect 585310 403058 585342 403294
rect 585578 403058 585662 403294
rect 585898 403058 585930 403294
rect 585310 383294 585930 403058
rect 585310 383058 585342 383294
rect 585578 383058 585662 383294
rect 585898 383058 585930 383294
rect 585310 363294 585930 383058
rect 585310 363058 585342 363294
rect 585578 363058 585662 363294
rect 585898 363058 585930 363294
rect 585310 343294 585930 363058
rect 585310 343058 585342 343294
rect 585578 343058 585662 343294
rect 585898 343058 585930 343294
rect 585310 323294 585930 343058
rect 585310 323058 585342 323294
rect 585578 323058 585662 323294
rect 585898 323058 585930 323294
rect 585310 303294 585930 323058
rect 585310 303058 585342 303294
rect 585578 303058 585662 303294
rect 585898 303058 585930 303294
rect 585310 283294 585930 303058
rect 585310 283058 585342 283294
rect 585578 283058 585662 283294
rect 585898 283058 585930 283294
rect 585310 263294 585930 283058
rect 585310 263058 585342 263294
rect 585578 263058 585662 263294
rect 585898 263058 585930 263294
rect 585310 243294 585930 263058
rect 585310 243058 585342 243294
rect 585578 243058 585662 243294
rect 585898 243058 585930 243294
rect 585310 223294 585930 243058
rect 585310 223058 585342 223294
rect 585578 223058 585662 223294
rect 585898 223058 585930 223294
rect 585310 203294 585930 223058
rect 585310 203058 585342 203294
rect 585578 203058 585662 203294
rect 585898 203058 585930 203294
rect 585310 183294 585930 203058
rect 585310 183058 585342 183294
rect 585578 183058 585662 183294
rect 585898 183058 585930 183294
rect 585310 163294 585930 183058
rect 585310 163058 585342 163294
rect 585578 163058 585662 163294
rect 585898 163058 585930 163294
rect 585310 143294 585930 163058
rect 585310 143058 585342 143294
rect 585578 143058 585662 143294
rect 585898 143058 585930 143294
rect 585310 123294 585930 143058
rect 585310 123058 585342 123294
rect 585578 123058 585662 123294
rect 585898 123058 585930 123294
rect 585310 103294 585930 123058
rect 585310 103058 585342 103294
rect 585578 103058 585662 103294
rect 585898 103058 585930 103294
rect 585310 83294 585930 103058
rect 585310 83058 585342 83294
rect 585578 83058 585662 83294
rect 585898 83058 585930 83294
rect 585310 63294 585930 83058
rect 585310 63058 585342 63294
rect 585578 63058 585662 63294
rect 585898 63058 585930 63294
rect 585310 43294 585930 63058
rect 585310 43058 585342 43294
rect 585578 43058 585662 43294
rect 585898 43058 585930 43294
rect 585310 23294 585930 43058
rect 585310 23058 585342 23294
rect 585578 23058 585662 23294
rect 585898 23058 585930 23294
rect 585310 3294 585930 23058
rect 585310 3058 585342 3294
rect 585578 3058 585662 3294
rect 585898 3058 585930 3294
rect 585310 -346 585930 3058
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 693294 586890 705242
rect 586270 693058 586302 693294
rect 586538 693058 586622 693294
rect 586858 693058 586890 693294
rect 586270 673294 586890 693058
rect 586270 673058 586302 673294
rect 586538 673058 586622 673294
rect 586858 673058 586890 673294
rect 586270 653294 586890 673058
rect 586270 653058 586302 653294
rect 586538 653058 586622 653294
rect 586858 653058 586890 653294
rect 586270 633294 586890 653058
rect 586270 633058 586302 633294
rect 586538 633058 586622 633294
rect 586858 633058 586890 633294
rect 586270 613294 586890 633058
rect 586270 613058 586302 613294
rect 586538 613058 586622 613294
rect 586858 613058 586890 613294
rect 586270 593294 586890 613058
rect 586270 593058 586302 593294
rect 586538 593058 586622 593294
rect 586858 593058 586890 593294
rect 586270 573294 586890 593058
rect 586270 573058 586302 573294
rect 586538 573058 586622 573294
rect 586858 573058 586890 573294
rect 586270 553294 586890 573058
rect 586270 553058 586302 553294
rect 586538 553058 586622 553294
rect 586858 553058 586890 553294
rect 586270 533294 586890 553058
rect 586270 533058 586302 533294
rect 586538 533058 586622 533294
rect 586858 533058 586890 533294
rect 586270 513294 586890 533058
rect 586270 513058 586302 513294
rect 586538 513058 586622 513294
rect 586858 513058 586890 513294
rect 586270 493294 586890 513058
rect 586270 493058 586302 493294
rect 586538 493058 586622 493294
rect 586858 493058 586890 493294
rect 586270 473294 586890 493058
rect 586270 473058 586302 473294
rect 586538 473058 586622 473294
rect 586858 473058 586890 473294
rect 586270 453294 586890 473058
rect 586270 453058 586302 453294
rect 586538 453058 586622 453294
rect 586858 453058 586890 453294
rect 586270 433294 586890 453058
rect 586270 433058 586302 433294
rect 586538 433058 586622 433294
rect 586858 433058 586890 433294
rect 586270 413294 586890 433058
rect 586270 413058 586302 413294
rect 586538 413058 586622 413294
rect 586858 413058 586890 413294
rect 586270 393294 586890 413058
rect 586270 393058 586302 393294
rect 586538 393058 586622 393294
rect 586858 393058 586890 393294
rect 586270 373294 586890 393058
rect 586270 373058 586302 373294
rect 586538 373058 586622 373294
rect 586858 373058 586890 373294
rect 586270 353294 586890 373058
rect 586270 353058 586302 353294
rect 586538 353058 586622 353294
rect 586858 353058 586890 353294
rect 586270 333294 586890 353058
rect 586270 333058 586302 333294
rect 586538 333058 586622 333294
rect 586858 333058 586890 333294
rect 586270 313294 586890 333058
rect 586270 313058 586302 313294
rect 586538 313058 586622 313294
rect 586858 313058 586890 313294
rect 586270 293294 586890 313058
rect 586270 293058 586302 293294
rect 586538 293058 586622 293294
rect 586858 293058 586890 293294
rect 586270 273294 586890 293058
rect 586270 273058 586302 273294
rect 586538 273058 586622 273294
rect 586858 273058 586890 273294
rect 586270 253294 586890 273058
rect 586270 253058 586302 253294
rect 586538 253058 586622 253294
rect 586858 253058 586890 253294
rect 586270 233294 586890 253058
rect 586270 233058 586302 233294
rect 586538 233058 586622 233294
rect 586858 233058 586890 233294
rect 586270 213294 586890 233058
rect 586270 213058 586302 213294
rect 586538 213058 586622 213294
rect 586858 213058 586890 213294
rect 586270 193294 586890 213058
rect 586270 193058 586302 193294
rect 586538 193058 586622 193294
rect 586858 193058 586890 193294
rect 586270 173294 586890 193058
rect 586270 173058 586302 173294
rect 586538 173058 586622 173294
rect 586858 173058 586890 173294
rect 586270 153294 586890 173058
rect 586270 153058 586302 153294
rect 586538 153058 586622 153294
rect 586858 153058 586890 153294
rect 586270 133294 586890 153058
rect 586270 133058 586302 133294
rect 586538 133058 586622 133294
rect 586858 133058 586890 133294
rect 586270 113294 586890 133058
rect 586270 113058 586302 113294
rect 586538 113058 586622 113294
rect 586858 113058 586890 113294
rect 586270 93294 586890 113058
rect 586270 93058 586302 93294
rect 586538 93058 586622 93294
rect 586858 93058 586890 93294
rect 586270 73294 586890 93058
rect 586270 73058 586302 73294
rect 586538 73058 586622 73294
rect 586858 73058 586890 73294
rect 586270 53294 586890 73058
rect 586270 53058 586302 53294
rect 586538 53058 586622 53294
rect 586858 53058 586890 53294
rect 586270 33294 586890 53058
rect 586270 33058 586302 33294
rect 586538 33058 586622 33294
rect 586858 33058 586890 33294
rect 586270 13294 586890 33058
rect 586270 13058 586302 13294
rect 586538 13058 586622 13294
rect 586858 13058 586890 13294
rect 586270 -1306 586890 13058
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 686954 587850 706202
rect 587230 686718 587262 686954
rect 587498 686718 587582 686954
rect 587818 686718 587850 686954
rect 587230 666954 587850 686718
rect 587230 666718 587262 666954
rect 587498 666718 587582 666954
rect 587818 666718 587850 666954
rect 587230 646954 587850 666718
rect 587230 646718 587262 646954
rect 587498 646718 587582 646954
rect 587818 646718 587850 646954
rect 587230 626954 587850 646718
rect 587230 626718 587262 626954
rect 587498 626718 587582 626954
rect 587818 626718 587850 626954
rect 587230 606954 587850 626718
rect 587230 606718 587262 606954
rect 587498 606718 587582 606954
rect 587818 606718 587850 606954
rect 587230 586954 587850 606718
rect 587230 586718 587262 586954
rect 587498 586718 587582 586954
rect 587818 586718 587850 586954
rect 587230 566954 587850 586718
rect 587230 566718 587262 566954
rect 587498 566718 587582 566954
rect 587818 566718 587850 566954
rect 587230 546954 587850 566718
rect 587230 546718 587262 546954
rect 587498 546718 587582 546954
rect 587818 546718 587850 546954
rect 587230 526954 587850 546718
rect 587230 526718 587262 526954
rect 587498 526718 587582 526954
rect 587818 526718 587850 526954
rect 587230 506954 587850 526718
rect 587230 506718 587262 506954
rect 587498 506718 587582 506954
rect 587818 506718 587850 506954
rect 587230 486954 587850 506718
rect 587230 486718 587262 486954
rect 587498 486718 587582 486954
rect 587818 486718 587850 486954
rect 587230 466954 587850 486718
rect 587230 466718 587262 466954
rect 587498 466718 587582 466954
rect 587818 466718 587850 466954
rect 587230 446954 587850 466718
rect 587230 446718 587262 446954
rect 587498 446718 587582 446954
rect 587818 446718 587850 446954
rect 587230 426954 587850 446718
rect 587230 426718 587262 426954
rect 587498 426718 587582 426954
rect 587818 426718 587850 426954
rect 587230 406954 587850 426718
rect 587230 406718 587262 406954
rect 587498 406718 587582 406954
rect 587818 406718 587850 406954
rect 587230 386954 587850 406718
rect 587230 386718 587262 386954
rect 587498 386718 587582 386954
rect 587818 386718 587850 386954
rect 587230 366954 587850 386718
rect 587230 366718 587262 366954
rect 587498 366718 587582 366954
rect 587818 366718 587850 366954
rect 587230 346954 587850 366718
rect 587230 346718 587262 346954
rect 587498 346718 587582 346954
rect 587818 346718 587850 346954
rect 587230 326954 587850 346718
rect 587230 326718 587262 326954
rect 587498 326718 587582 326954
rect 587818 326718 587850 326954
rect 587230 306954 587850 326718
rect 587230 306718 587262 306954
rect 587498 306718 587582 306954
rect 587818 306718 587850 306954
rect 587230 286954 587850 306718
rect 587230 286718 587262 286954
rect 587498 286718 587582 286954
rect 587818 286718 587850 286954
rect 587230 266954 587850 286718
rect 587230 266718 587262 266954
rect 587498 266718 587582 266954
rect 587818 266718 587850 266954
rect 587230 246954 587850 266718
rect 587230 246718 587262 246954
rect 587498 246718 587582 246954
rect 587818 246718 587850 246954
rect 587230 226954 587850 246718
rect 587230 226718 587262 226954
rect 587498 226718 587582 226954
rect 587818 226718 587850 226954
rect 587230 206954 587850 226718
rect 587230 206718 587262 206954
rect 587498 206718 587582 206954
rect 587818 206718 587850 206954
rect 587230 186954 587850 206718
rect 587230 186718 587262 186954
rect 587498 186718 587582 186954
rect 587818 186718 587850 186954
rect 587230 166954 587850 186718
rect 587230 166718 587262 166954
rect 587498 166718 587582 166954
rect 587818 166718 587850 166954
rect 587230 146954 587850 166718
rect 587230 146718 587262 146954
rect 587498 146718 587582 146954
rect 587818 146718 587850 146954
rect 587230 126954 587850 146718
rect 587230 126718 587262 126954
rect 587498 126718 587582 126954
rect 587818 126718 587850 126954
rect 587230 106954 587850 126718
rect 587230 106718 587262 106954
rect 587498 106718 587582 106954
rect 587818 106718 587850 106954
rect 587230 86954 587850 106718
rect 587230 86718 587262 86954
rect 587498 86718 587582 86954
rect 587818 86718 587850 86954
rect 587230 66954 587850 86718
rect 587230 66718 587262 66954
rect 587498 66718 587582 66954
rect 587818 66718 587850 66954
rect 587230 46954 587850 66718
rect 587230 46718 587262 46954
rect 587498 46718 587582 46954
rect 587818 46718 587850 46954
rect 587230 26954 587850 46718
rect 587230 26718 587262 26954
rect 587498 26718 587582 26954
rect 587818 26718 587850 26954
rect 587230 6954 587850 26718
rect 587230 6718 587262 6954
rect 587498 6718 587582 6954
rect 587818 6718 587850 6954
rect 587230 -2266 587850 6718
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 696954 588810 707162
rect 588190 696718 588222 696954
rect 588458 696718 588542 696954
rect 588778 696718 588810 696954
rect 588190 676954 588810 696718
rect 588190 676718 588222 676954
rect 588458 676718 588542 676954
rect 588778 676718 588810 676954
rect 588190 656954 588810 676718
rect 588190 656718 588222 656954
rect 588458 656718 588542 656954
rect 588778 656718 588810 656954
rect 588190 636954 588810 656718
rect 588190 636718 588222 636954
rect 588458 636718 588542 636954
rect 588778 636718 588810 636954
rect 588190 616954 588810 636718
rect 588190 616718 588222 616954
rect 588458 616718 588542 616954
rect 588778 616718 588810 616954
rect 588190 596954 588810 616718
rect 588190 596718 588222 596954
rect 588458 596718 588542 596954
rect 588778 596718 588810 596954
rect 588190 576954 588810 596718
rect 588190 576718 588222 576954
rect 588458 576718 588542 576954
rect 588778 576718 588810 576954
rect 588190 556954 588810 576718
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 536954 588810 556718
rect 588190 536718 588222 536954
rect 588458 536718 588542 536954
rect 588778 536718 588810 536954
rect 588190 516954 588810 536718
rect 588190 516718 588222 516954
rect 588458 516718 588542 516954
rect 588778 516718 588810 516954
rect 588190 496954 588810 516718
rect 588190 496718 588222 496954
rect 588458 496718 588542 496954
rect 588778 496718 588810 496954
rect 588190 476954 588810 496718
rect 588190 476718 588222 476954
rect 588458 476718 588542 476954
rect 588778 476718 588810 476954
rect 588190 456954 588810 476718
rect 588190 456718 588222 456954
rect 588458 456718 588542 456954
rect 588778 456718 588810 456954
rect 588190 436954 588810 456718
rect 588190 436718 588222 436954
rect 588458 436718 588542 436954
rect 588778 436718 588810 436954
rect 588190 416954 588810 436718
rect 588190 416718 588222 416954
rect 588458 416718 588542 416954
rect 588778 416718 588810 416954
rect 588190 396954 588810 416718
rect 588190 396718 588222 396954
rect 588458 396718 588542 396954
rect 588778 396718 588810 396954
rect 588190 376954 588810 396718
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 356954 588810 376718
rect 588190 356718 588222 356954
rect 588458 356718 588542 356954
rect 588778 356718 588810 356954
rect 588190 336954 588810 356718
rect 588190 336718 588222 336954
rect 588458 336718 588542 336954
rect 588778 336718 588810 336954
rect 588190 316954 588810 336718
rect 588190 316718 588222 316954
rect 588458 316718 588542 316954
rect 588778 316718 588810 316954
rect 588190 296954 588810 316718
rect 588190 296718 588222 296954
rect 588458 296718 588542 296954
rect 588778 296718 588810 296954
rect 588190 276954 588810 296718
rect 588190 276718 588222 276954
rect 588458 276718 588542 276954
rect 588778 276718 588810 276954
rect 588190 256954 588810 276718
rect 588190 256718 588222 256954
rect 588458 256718 588542 256954
rect 588778 256718 588810 256954
rect 588190 236954 588810 256718
rect 588190 236718 588222 236954
rect 588458 236718 588542 236954
rect 588778 236718 588810 236954
rect 588190 216954 588810 236718
rect 588190 216718 588222 216954
rect 588458 216718 588542 216954
rect 588778 216718 588810 216954
rect 588190 196954 588810 216718
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 176954 588810 196718
rect 588190 176718 588222 176954
rect 588458 176718 588542 176954
rect 588778 176718 588810 176954
rect 588190 156954 588810 176718
rect 588190 156718 588222 156954
rect 588458 156718 588542 156954
rect 588778 156718 588810 156954
rect 588190 136954 588810 156718
rect 588190 136718 588222 136954
rect 588458 136718 588542 136954
rect 588778 136718 588810 136954
rect 588190 116954 588810 136718
rect 588190 116718 588222 116954
rect 588458 116718 588542 116954
rect 588778 116718 588810 116954
rect 588190 96954 588810 116718
rect 588190 96718 588222 96954
rect 588458 96718 588542 96954
rect 588778 96718 588810 96954
rect 588190 76954 588810 96718
rect 588190 76718 588222 76954
rect 588458 76718 588542 76954
rect 588778 76718 588810 76954
rect 588190 56954 588810 76718
rect 588190 56718 588222 56954
rect 588458 56718 588542 56954
rect 588778 56718 588810 56954
rect 588190 36954 588810 56718
rect 588190 36718 588222 36954
rect 588458 36718 588542 36954
rect 588778 36718 588810 36954
rect 588190 16954 588810 36718
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 -3226 588810 16718
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 690614 589770 708122
rect 589150 690378 589182 690614
rect 589418 690378 589502 690614
rect 589738 690378 589770 690614
rect 589150 670614 589770 690378
rect 589150 670378 589182 670614
rect 589418 670378 589502 670614
rect 589738 670378 589770 670614
rect 589150 650614 589770 670378
rect 589150 650378 589182 650614
rect 589418 650378 589502 650614
rect 589738 650378 589770 650614
rect 589150 630614 589770 650378
rect 589150 630378 589182 630614
rect 589418 630378 589502 630614
rect 589738 630378 589770 630614
rect 589150 610614 589770 630378
rect 589150 610378 589182 610614
rect 589418 610378 589502 610614
rect 589738 610378 589770 610614
rect 589150 590614 589770 610378
rect 589150 590378 589182 590614
rect 589418 590378 589502 590614
rect 589738 590378 589770 590614
rect 589150 570614 589770 590378
rect 589150 570378 589182 570614
rect 589418 570378 589502 570614
rect 589738 570378 589770 570614
rect 589150 550614 589770 570378
rect 589150 550378 589182 550614
rect 589418 550378 589502 550614
rect 589738 550378 589770 550614
rect 589150 530614 589770 550378
rect 589150 530378 589182 530614
rect 589418 530378 589502 530614
rect 589738 530378 589770 530614
rect 589150 510614 589770 530378
rect 589150 510378 589182 510614
rect 589418 510378 589502 510614
rect 589738 510378 589770 510614
rect 589150 490614 589770 510378
rect 589150 490378 589182 490614
rect 589418 490378 589502 490614
rect 589738 490378 589770 490614
rect 589150 470614 589770 490378
rect 589150 470378 589182 470614
rect 589418 470378 589502 470614
rect 589738 470378 589770 470614
rect 589150 450614 589770 470378
rect 589150 450378 589182 450614
rect 589418 450378 589502 450614
rect 589738 450378 589770 450614
rect 589150 430614 589770 450378
rect 589150 430378 589182 430614
rect 589418 430378 589502 430614
rect 589738 430378 589770 430614
rect 589150 410614 589770 430378
rect 589150 410378 589182 410614
rect 589418 410378 589502 410614
rect 589738 410378 589770 410614
rect 589150 390614 589770 410378
rect 589150 390378 589182 390614
rect 589418 390378 589502 390614
rect 589738 390378 589770 390614
rect 589150 370614 589770 390378
rect 589150 370378 589182 370614
rect 589418 370378 589502 370614
rect 589738 370378 589770 370614
rect 589150 350614 589770 370378
rect 589150 350378 589182 350614
rect 589418 350378 589502 350614
rect 589738 350378 589770 350614
rect 589150 330614 589770 350378
rect 589150 330378 589182 330614
rect 589418 330378 589502 330614
rect 589738 330378 589770 330614
rect 589150 310614 589770 330378
rect 589150 310378 589182 310614
rect 589418 310378 589502 310614
rect 589738 310378 589770 310614
rect 589150 290614 589770 310378
rect 589150 290378 589182 290614
rect 589418 290378 589502 290614
rect 589738 290378 589770 290614
rect 589150 270614 589770 290378
rect 589150 270378 589182 270614
rect 589418 270378 589502 270614
rect 589738 270378 589770 270614
rect 589150 250614 589770 270378
rect 589150 250378 589182 250614
rect 589418 250378 589502 250614
rect 589738 250378 589770 250614
rect 589150 230614 589770 250378
rect 589150 230378 589182 230614
rect 589418 230378 589502 230614
rect 589738 230378 589770 230614
rect 589150 210614 589770 230378
rect 589150 210378 589182 210614
rect 589418 210378 589502 210614
rect 589738 210378 589770 210614
rect 589150 190614 589770 210378
rect 589150 190378 589182 190614
rect 589418 190378 589502 190614
rect 589738 190378 589770 190614
rect 589150 170614 589770 190378
rect 589150 170378 589182 170614
rect 589418 170378 589502 170614
rect 589738 170378 589770 170614
rect 589150 150614 589770 170378
rect 589150 150378 589182 150614
rect 589418 150378 589502 150614
rect 589738 150378 589770 150614
rect 589150 130614 589770 150378
rect 589150 130378 589182 130614
rect 589418 130378 589502 130614
rect 589738 130378 589770 130614
rect 589150 110614 589770 130378
rect 589150 110378 589182 110614
rect 589418 110378 589502 110614
rect 589738 110378 589770 110614
rect 589150 90614 589770 110378
rect 589150 90378 589182 90614
rect 589418 90378 589502 90614
rect 589738 90378 589770 90614
rect 589150 70614 589770 90378
rect 589150 70378 589182 70614
rect 589418 70378 589502 70614
rect 589738 70378 589770 70614
rect 589150 50614 589770 70378
rect 589150 50378 589182 50614
rect 589418 50378 589502 50614
rect 589738 50378 589770 50614
rect 589150 30614 589770 50378
rect 589150 30378 589182 30614
rect 589418 30378 589502 30614
rect 589738 30378 589770 30614
rect 589150 10614 589770 30378
rect 589150 10378 589182 10614
rect 589418 10378 589502 10614
rect 589738 10378 589770 10614
rect 589150 -4186 589770 10378
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 700614 590730 709082
rect 590110 700378 590142 700614
rect 590378 700378 590462 700614
rect 590698 700378 590730 700614
rect 590110 680614 590730 700378
rect 590110 680378 590142 680614
rect 590378 680378 590462 680614
rect 590698 680378 590730 680614
rect 590110 660614 590730 680378
rect 590110 660378 590142 660614
rect 590378 660378 590462 660614
rect 590698 660378 590730 660614
rect 590110 640614 590730 660378
rect 590110 640378 590142 640614
rect 590378 640378 590462 640614
rect 590698 640378 590730 640614
rect 590110 620614 590730 640378
rect 590110 620378 590142 620614
rect 590378 620378 590462 620614
rect 590698 620378 590730 620614
rect 590110 600614 590730 620378
rect 590110 600378 590142 600614
rect 590378 600378 590462 600614
rect 590698 600378 590730 600614
rect 590110 580614 590730 600378
rect 590110 580378 590142 580614
rect 590378 580378 590462 580614
rect 590698 580378 590730 580614
rect 590110 560614 590730 580378
rect 590110 560378 590142 560614
rect 590378 560378 590462 560614
rect 590698 560378 590730 560614
rect 590110 540614 590730 560378
rect 590110 540378 590142 540614
rect 590378 540378 590462 540614
rect 590698 540378 590730 540614
rect 590110 520614 590730 540378
rect 590110 520378 590142 520614
rect 590378 520378 590462 520614
rect 590698 520378 590730 520614
rect 590110 500614 590730 520378
rect 590110 500378 590142 500614
rect 590378 500378 590462 500614
rect 590698 500378 590730 500614
rect 590110 480614 590730 500378
rect 590110 480378 590142 480614
rect 590378 480378 590462 480614
rect 590698 480378 590730 480614
rect 590110 460614 590730 480378
rect 590110 460378 590142 460614
rect 590378 460378 590462 460614
rect 590698 460378 590730 460614
rect 590110 440614 590730 460378
rect 590110 440378 590142 440614
rect 590378 440378 590462 440614
rect 590698 440378 590730 440614
rect 590110 420614 590730 440378
rect 590110 420378 590142 420614
rect 590378 420378 590462 420614
rect 590698 420378 590730 420614
rect 590110 400614 590730 420378
rect 590110 400378 590142 400614
rect 590378 400378 590462 400614
rect 590698 400378 590730 400614
rect 590110 380614 590730 400378
rect 590110 380378 590142 380614
rect 590378 380378 590462 380614
rect 590698 380378 590730 380614
rect 590110 360614 590730 380378
rect 590110 360378 590142 360614
rect 590378 360378 590462 360614
rect 590698 360378 590730 360614
rect 590110 340614 590730 360378
rect 590110 340378 590142 340614
rect 590378 340378 590462 340614
rect 590698 340378 590730 340614
rect 590110 320614 590730 340378
rect 590110 320378 590142 320614
rect 590378 320378 590462 320614
rect 590698 320378 590730 320614
rect 590110 300614 590730 320378
rect 590110 300378 590142 300614
rect 590378 300378 590462 300614
rect 590698 300378 590730 300614
rect 590110 280614 590730 300378
rect 590110 280378 590142 280614
rect 590378 280378 590462 280614
rect 590698 280378 590730 280614
rect 590110 260614 590730 280378
rect 590110 260378 590142 260614
rect 590378 260378 590462 260614
rect 590698 260378 590730 260614
rect 590110 240614 590730 260378
rect 590110 240378 590142 240614
rect 590378 240378 590462 240614
rect 590698 240378 590730 240614
rect 590110 220614 590730 240378
rect 590110 220378 590142 220614
rect 590378 220378 590462 220614
rect 590698 220378 590730 220614
rect 590110 200614 590730 220378
rect 590110 200378 590142 200614
rect 590378 200378 590462 200614
rect 590698 200378 590730 200614
rect 590110 180614 590730 200378
rect 590110 180378 590142 180614
rect 590378 180378 590462 180614
rect 590698 180378 590730 180614
rect 590110 160614 590730 180378
rect 590110 160378 590142 160614
rect 590378 160378 590462 160614
rect 590698 160378 590730 160614
rect 590110 140614 590730 160378
rect 590110 140378 590142 140614
rect 590378 140378 590462 140614
rect 590698 140378 590730 140614
rect 590110 120614 590730 140378
rect 590110 120378 590142 120614
rect 590378 120378 590462 120614
rect 590698 120378 590730 120614
rect 590110 100614 590730 120378
rect 590110 100378 590142 100614
rect 590378 100378 590462 100614
rect 590698 100378 590730 100614
rect 590110 80614 590730 100378
rect 590110 80378 590142 80614
rect 590378 80378 590462 80614
rect 590698 80378 590730 80614
rect 590110 60614 590730 80378
rect 590110 60378 590142 60614
rect 590378 60378 590462 60614
rect 590698 60378 590730 60614
rect 590110 40614 590730 60378
rect 590110 40378 590142 40614
rect 590378 40378 590462 40614
rect 590698 40378 590730 40614
rect 590110 20614 590730 40378
rect 590110 20378 590142 20614
rect 590378 20378 590462 20614
rect 590698 20378 590730 20614
rect 579234 -5382 579266 -5146
rect 579502 -5382 579586 -5146
rect 579822 -5382 579854 -5146
rect 579234 -5466 579854 -5382
rect 579234 -5702 579266 -5466
rect 579502 -5702 579586 -5466
rect 579822 -5702 579854 -5466
rect 579234 -5734 579854 -5702
rect 590110 -5146 590730 20378
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 694274 591690 710042
rect 591070 694038 591102 694274
rect 591338 694038 591422 694274
rect 591658 694038 591690 694274
rect 591070 674274 591690 694038
rect 591070 674038 591102 674274
rect 591338 674038 591422 674274
rect 591658 674038 591690 674274
rect 591070 654274 591690 674038
rect 591070 654038 591102 654274
rect 591338 654038 591422 654274
rect 591658 654038 591690 654274
rect 591070 634274 591690 654038
rect 591070 634038 591102 634274
rect 591338 634038 591422 634274
rect 591658 634038 591690 634274
rect 591070 614274 591690 634038
rect 591070 614038 591102 614274
rect 591338 614038 591422 614274
rect 591658 614038 591690 614274
rect 591070 594274 591690 614038
rect 591070 594038 591102 594274
rect 591338 594038 591422 594274
rect 591658 594038 591690 594274
rect 591070 574274 591690 594038
rect 591070 574038 591102 574274
rect 591338 574038 591422 574274
rect 591658 574038 591690 574274
rect 591070 554274 591690 574038
rect 591070 554038 591102 554274
rect 591338 554038 591422 554274
rect 591658 554038 591690 554274
rect 591070 534274 591690 554038
rect 591070 534038 591102 534274
rect 591338 534038 591422 534274
rect 591658 534038 591690 534274
rect 591070 514274 591690 534038
rect 591070 514038 591102 514274
rect 591338 514038 591422 514274
rect 591658 514038 591690 514274
rect 591070 494274 591690 514038
rect 591070 494038 591102 494274
rect 591338 494038 591422 494274
rect 591658 494038 591690 494274
rect 591070 474274 591690 494038
rect 591070 474038 591102 474274
rect 591338 474038 591422 474274
rect 591658 474038 591690 474274
rect 591070 454274 591690 474038
rect 591070 454038 591102 454274
rect 591338 454038 591422 454274
rect 591658 454038 591690 454274
rect 591070 434274 591690 454038
rect 591070 434038 591102 434274
rect 591338 434038 591422 434274
rect 591658 434038 591690 434274
rect 591070 414274 591690 434038
rect 591070 414038 591102 414274
rect 591338 414038 591422 414274
rect 591658 414038 591690 414274
rect 591070 394274 591690 414038
rect 591070 394038 591102 394274
rect 591338 394038 591422 394274
rect 591658 394038 591690 394274
rect 591070 374274 591690 394038
rect 591070 374038 591102 374274
rect 591338 374038 591422 374274
rect 591658 374038 591690 374274
rect 591070 354274 591690 374038
rect 591070 354038 591102 354274
rect 591338 354038 591422 354274
rect 591658 354038 591690 354274
rect 591070 334274 591690 354038
rect 591070 334038 591102 334274
rect 591338 334038 591422 334274
rect 591658 334038 591690 334274
rect 591070 314274 591690 334038
rect 591070 314038 591102 314274
rect 591338 314038 591422 314274
rect 591658 314038 591690 314274
rect 591070 294274 591690 314038
rect 591070 294038 591102 294274
rect 591338 294038 591422 294274
rect 591658 294038 591690 294274
rect 591070 274274 591690 294038
rect 591070 274038 591102 274274
rect 591338 274038 591422 274274
rect 591658 274038 591690 274274
rect 591070 254274 591690 274038
rect 591070 254038 591102 254274
rect 591338 254038 591422 254274
rect 591658 254038 591690 254274
rect 591070 234274 591690 254038
rect 591070 234038 591102 234274
rect 591338 234038 591422 234274
rect 591658 234038 591690 234274
rect 591070 214274 591690 234038
rect 591070 214038 591102 214274
rect 591338 214038 591422 214274
rect 591658 214038 591690 214274
rect 591070 194274 591690 214038
rect 591070 194038 591102 194274
rect 591338 194038 591422 194274
rect 591658 194038 591690 194274
rect 591070 174274 591690 194038
rect 591070 174038 591102 174274
rect 591338 174038 591422 174274
rect 591658 174038 591690 174274
rect 591070 154274 591690 174038
rect 591070 154038 591102 154274
rect 591338 154038 591422 154274
rect 591658 154038 591690 154274
rect 591070 134274 591690 154038
rect 591070 134038 591102 134274
rect 591338 134038 591422 134274
rect 591658 134038 591690 134274
rect 591070 114274 591690 134038
rect 591070 114038 591102 114274
rect 591338 114038 591422 114274
rect 591658 114038 591690 114274
rect 591070 94274 591690 114038
rect 591070 94038 591102 94274
rect 591338 94038 591422 94274
rect 591658 94038 591690 94274
rect 591070 74274 591690 94038
rect 591070 74038 591102 74274
rect 591338 74038 591422 74274
rect 591658 74038 591690 74274
rect 591070 54274 591690 74038
rect 591070 54038 591102 54274
rect 591338 54038 591422 54274
rect 591658 54038 591690 54274
rect 591070 34274 591690 54038
rect 591070 34038 591102 34274
rect 591338 34038 591422 34274
rect 591658 34038 591690 34274
rect 591070 14274 591690 34038
rect 591070 14038 591102 14274
rect 591338 14038 591422 14274
rect 591658 14038 591690 14274
rect 572954 -6342 572986 -6106
rect 573222 -6342 573306 -6106
rect 573542 -6342 573574 -6106
rect 572954 -6426 573574 -6342
rect 572954 -6662 572986 -6426
rect 573222 -6662 573306 -6426
rect 573542 -6662 573574 -6426
rect 572954 -7654 573574 -6662
rect 591070 -6106 591690 14038
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 684274 592650 711002
rect 592030 684038 592062 684274
rect 592298 684038 592382 684274
rect 592618 684038 592650 684274
rect 592030 664274 592650 684038
rect 592030 664038 592062 664274
rect 592298 664038 592382 664274
rect 592618 664038 592650 664274
rect 592030 644274 592650 664038
rect 592030 644038 592062 644274
rect 592298 644038 592382 644274
rect 592618 644038 592650 644274
rect 592030 624274 592650 644038
rect 592030 624038 592062 624274
rect 592298 624038 592382 624274
rect 592618 624038 592650 624274
rect 592030 604274 592650 624038
rect 592030 604038 592062 604274
rect 592298 604038 592382 604274
rect 592618 604038 592650 604274
rect 592030 584274 592650 604038
rect 592030 584038 592062 584274
rect 592298 584038 592382 584274
rect 592618 584038 592650 584274
rect 592030 564274 592650 584038
rect 592030 564038 592062 564274
rect 592298 564038 592382 564274
rect 592618 564038 592650 564274
rect 592030 544274 592650 564038
rect 592030 544038 592062 544274
rect 592298 544038 592382 544274
rect 592618 544038 592650 544274
rect 592030 524274 592650 544038
rect 592030 524038 592062 524274
rect 592298 524038 592382 524274
rect 592618 524038 592650 524274
rect 592030 504274 592650 524038
rect 592030 504038 592062 504274
rect 592298 504038 592382 504274
rect 592618 504038 592650 504274
rect 592030 484274 592650 504038
rect 592030 484038 592062 484274
rect 592298 484038 592382 484274
rect 592618 484038 592650 484274
rect 592030 464274 592650 484038
rect 592030 464038 592062 464274
rect 592298 464038 592382 464274
rect 592618 464038 592650 464274
rect 592030 444274 592650 464038
rect 592030 444038 592062 444274
rect 592298 444038 592382 444274
rect 592618 444038 592650 444274
rect 592030 424274 592650 444038
rect 592030 424038 592062 424274
rect 592298 424038 592382 424274
rect 592618 424038 592650 424274
rect 592030 404274 592650 424038
rect 592030 404038 592062 404274
rect 592298 404038 592382 404274
rect 592618 404038 592650 404274
rect 592030 384274 592650 404038
rect 592030 384038 592062 384274
rect 592298 384038 592382 384274
rect 592618 384038 592650 384274
rect 592030 364274 592650 384038
rect 592030 364038 592062 364274
rect 592298 364038 592382 364274
rect 592618 364038 592650 364274
rect 592030 344274 592650 364038
rect 592030 344038 592062 344274
rect 592298 344038 592382 344274
rect 592618 344038 592650 344274
rect 592030 324274 592650 344038
rect 592030 324038 592062 324274
rect 592298 324038 592382 324274
rect 592618 324038 592650 324274
rect 592030 304274 592650 324038
rect 592030 304038 592062 304274
rect 592298 304038 592382 304274
rect 592618 304038 592650 304274
rect 592030 284274 592650 304038
rect 592030 284038 592062 284274
rect 592298 284038 592382 284274
rect 592618 284038 592650 284274
rect 592030 264274 592650 284038
rect 592030 264038 592062 264274
rect 592298 264038 592382 264274
rect 592618 264038 592650 264274
rect 592030 244274 592650 264038
rect 592030 244038 592062 244274
rect 592298 244038 592382 244274
rect 592618 244038 592650 244274
rect 592030 224274 592650 244038
rect 592030 224038 592062 224274
rect 592298 224038 592382 224274
rect 592618 224038 592650 224274
rect 592030 204274 592650 224038
rect 592030 204038 592062 204274
rect 592298 204038 592382 204274
rect 592618 204038 592650 204274
rect 592030 184274 592650 204038
rect 592030 184038 592062 184274
rect 592298 184038 592382 184274
rect 592618 184038 592650 184274
rect 592030 164274 592650 184038
rect 592030 164038 592062 164274
rect 592298 164038 592382 164274
rect 592618 164038 592650 164274
rect 592030 144274 592650 164038
rect 592030 144038 592062 144274
rect 592298 144038 592382 144274
rect 592618 144038 592650 144274
rect 592030 124274 592650 144038
rect 592030 124038 592062 124274
rect 592298 124038 592382 124274
rect 592618 124038 592650 124274
rect 592030 104274 592650 124038
rect 592030 104038 592062 104274
rect 592298 104038 592382 104274
rect 592618 104038 592650 104274
rect 592030 84274 592650 104038
rect 592030 84038 592062 84274
rect 592298 84038 592382 84274
rect 592618 84038 592650 84274
rect 592030 64274 592650 84038
rect 592030 64038 592062 64274
rect 592298 64038 592382 64274
rect 592618 64038 592650 64274
rect 592030 44274 592650 64038
rect 592030 44038 592062 44274
rect 592298 44038 592382 44274
rect 592618 44038 592650 44274
rect 592030 24274 592650 44038
rect 592030 24038 592062 24274
rect 592298 24038 592382 24274
rect 592618 24038 592650 24274
rect 592030 -7066 592650 24038
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 684038 -8458 684274
rect -8374 684038 -8138 684274
rect -8694 664038 -8458 664274
rect -8374 664038 -8138 664274
rect -8694 644038 -8458 644274
rect -8374 644038 -8138 644274
rect -8694 624038 -8458 624274
rect -8374 624038 -8138 624274
rect -8694 604038 -8458 604274
rect -8374 604038 -8138 604274
rect -8694 584038 -8458 584274
rect -8374 584038 -8138 584274
rect -8694 564038 -8458 564274
rect -8374 564038 -8138 564274
rect -8694 544038 -8458 544274
rect -8374 544038 -8138 544274
rect -8694 524038 -8458 524274
rect -8374 524038 -8138 524274
rect -8694 504038 -8458 504274
rect -8374 504038 -8138 504274
rect -8694 484038 -8458 484274
rect -8374 484038 -8138 484274
rect -8694 464038 -8458 464274
rect -8374 464038 -8138 464274
rect -8694 444038 -8458 444274
rect -8374 444038 -8138 444274
rect -8694 424038 -8458 424274
rect -8374 424038 -8138 424274
rect -8694 404038 -8458 404274
rect -8374 404038 -8138 404274
rect -8694 384038 -8458 384274
rect -8374 384038 -8138 384274
rect -8694 364038 -8458 364274
rect -8374 364038 -8138 364274
rect -8694 344038 -8458 344274
rect -8374 344038 -8138 344274
rect -8694 324038 -8458 324274
rect -8374 324038 -8138 324274
rect -8694 304038 -8458 304274
rect -8374 304038 -8138 304274
rect -8694 284038 -8458 284274
rect -8374 284038 -8138 284274
rect -8694 264038 -8458 264274
rect -8374 264038 -8138 264274
rect -8694 244038 -8458 244274
rect -8374 244038 -8138 244274
rect -8694 224038 -8458 224274
rect -8374 224038 -8138 224274
rect -8694 204038 -8458 204274
rect -8374 204038 -8138 204274
rect -8694 184038 -8458 184274
rect -8374 184038 -8138 184274
rect -8694 164038 -8458 164274
rect -8374 164038 -8138 164274
rect -8694 144038 -8458 144274
rect -8374 144038 -8138 144274
rect -8694 124038 -8458 124274
rect -8374 124038 -8138 124274
rect -8694 104038 -8458 104274
rect -8374 104038 -8138 104274
rect -8694 84038 -8458 84274
rect -8374 84038 -8138 84274
rect -8694 64038 -8458 64274
rect -8374 64038 -8138 64274
rect -8694 44038 -8458 44274
rect -8374 44038 -8138 44274
rect -8694 24038 -8458 24274
rect -8374 24038 -8138 24274
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 694038 -7498 694274
rect -7414 694038 -7178 694274
rect -7734 674038 -7498 674274
rect -7414 674038 -7178 674274
rect -7734 654038 -7498 654274
rect -7414 654038 -7178 654274
rect -7734 634038 -7498 634274
rect -7414 634038 -7178 634274
rect -7734 614038 -7498 614274
rect -7414 614038 -7178 614274
rect -7734 594038 -7498 594274
rect -7414 594038 -7178 594274
rect -7734 574038 -7498 574274
rect -7414 574038 -7178 574274
rect -7734 554038 -7498 554274
rect -7414 554038 -7178 554274
rect -7734 534038 -7498 534274
rect -7414 534038 -7178 534274
rect -7734 514038 -7498 514274
rect -7414 514038 -7178 514274
rect -7734 494038 -7498 494274
rect -7414 494038 -7178 494274
rect -7734 474038 -7498 474274
rect -7414 474038 -7178 474274
rect -7734 454038 -7498 454274
rect -7414 454038 -7178 454274
rect -7734 434038 -7498 434274
rect -7414 434038 -7178 434274
rect -7734 414038 -7498 414274
rect -7414 414038 -7178 414274
rect -7734 394038 -7498 394274
rect -7414 394038 -7178 394274
rect -7734 374038 -7498 374274
rect -7414 374038 -7178 374274
rect -7734 354038 -7498 354274
rect -7414 354038 -7178 354274
rect -7734 334038 -7498 334274
rect -7414 334038 -7178 334274
rect -7734 314038 -7498 314274
rect -7414 314038 -7178 314274
rect -7734 294038 -7498 294274
rect -7414 294038 -7178 294274
rect -7734 274038 -7498 274274
rect -7414 274038 -7178 274274
rect -7734 254038 -7498 254274
rect -7414 254038 -7178 254274
rect -7734 234038 -7498 234274
rect -7414 234038 -7178 234274
rect -7734 214038 -7498 214274
rect -7414 214038 -7178 214274
rect -7734 194038 -7498 194274
rect -7414 194038 -7178 194274
rect -7734 174038 -7498 174274
rect -7414 174038 -7178 174274
rect -7734 154038 -7498 154274
rect -7414 154038 -7178 154274
rect -7734 134038 -7498 134274
rect -7414 134038 -7178 134274
rect -7734 114038 -7498 114274
rect -7414 114038 -7178 114274
rect -7734 94038 -7498 94274
rect -7414 94038 -7178 94274
rect -7734 74038 -7498 74274
rect -7414 74038 -7178 74274
rect -7734 54038 -7498 54274
rect -7414 54038 -7178 54274
rect -7734 34038 -7498 34274
rect -7414 34038 -7178 34274
rect -7734 14038 -7498 14274
rect -7414 14038 -7178 14274
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 700378 -6538 700614
rect -6454 700378 -6218 700614
rect -6774 680378 -6538 680614
rect -6454 680378 -6218 680614
rect -6774 660378 -6538 660614
rect -6454 660378 -6218 660614
rect -6774 640378 -6538 640614
rect -6454 640378 -6218 640614
rect -6774 620378 -6538 620614
rect -6454 620378 -6218 620614
rect -6774 600378 -6538 600614
rect -6454 600378 -6218 600614
rect -6774 580378 -6538 580614
rect -6454 580378 -6218 580614
rect -6774 560378 -6538 560614
rect -6454 560378 -6218 560614
rect -6774 540378 -6538 540614
rect -6454 540378 -6218 540614
rect -6774 520378 -6538 520614
rect -6454 520378 -6218 520614
rect -6774 500378 -6538 500614
rect -6454 500378 -6218 500614
rect -6774 480378 -6538 480614
rect -6454 480378 -6218 480614
rect -6774 460378 -6538 460614
rect -6454 460378 -6218 460614
rect -6774 440378 -6538 440614
rect -6454 440378 -6218 440614
rect -6774 420378 -6538 420614
rect -6454 420378 -6218 420614
rect -6774 400378 -6538 400614
rect -6454 400378 -6218 400614
rect -6774 380378 -6538 380614
rect -6454 380378 -6218 380614
rect -6774 360378 -6538 360614
rect -6454 360378 -6218 360614
rect -6774 340378 -6538 340614
rect -6454 340378 -6218 340614
rect -6774 320378 -6538 320614
rect -6454 320378 -6218 320614
rect -6774 300378 -6538 300614
rect -6454 300378 -6218 300614
rect -6774 280378 -6538 280614
rect -6454 280378 -6218 280614
rect -6774 260378 -6538 260614
rect -6454 260378 -6218 260614
rect -6774 240378 -6538 240614
rect -6454 240378 -6218 240614
rect -6774 220378 -6538 220614
rect -6454 220378 -6218 220614
rect -6774 200378 -6538 200614
rect -6454 200378 -6218 200614
rect -6774 180378 -6538 180614
rect -6454 180378 -6218 180614
rect -6774 160378 -6538 160614
rect -6454 160378 -6218 160614
rect -6774 140378 -6538 140614
rect -6454 140378 -6218 140614
rect -6774 120378 -6538 120614
rect -6454 120378 -6218 120614
rect -6774 100378 -6538 100614
rect -6454 100378 -6218 100614
rect -6774 80378 -6538 80614
rect -6454 80378 -6218 80614
rect -6774 60378 -6538 60614
rect -6454 60378 -6218 60614
rect -6774 40378 -6538 40614
rect -6454 40378 -6218 40614
rect -6774 20378 -6538 20614
rect -6454 20378 -6218 20614
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 690378 -5578 690614
rect -5494 690378 -5258 690614
rect -5814 670378 -5578 670614
rect -5494 670378 -5258 670614
rect -5814 650378 -5578 650614
rect -5494 650378 -5258 650614
rect -5814 630378 -5578 630614
rect -5494 630378 -5258 630614
rect -5814 610378 -5578 610614
rect -5494 610378 -5258 610614
rect -5814 590378 -5578 590614
rect -5494 590378 -5258 590614
rect -5814 570378 -5578 570614
rect -5494 570378 -5258 570614
rect -5814 550378 -5578 550614
rect -5494 550378 -5258 550614
rect -5814 530378 -5578 530614
rect -5494 530378 -5258 530614
rect -5814 510378 -5578 510614
rect -5494 510378 -5258 510614
rect -5814 490378 -5578 490614
rect -5494 490378 -5258 490614
rect -5814 470378 -5578 470614
rect -5494 470378 -5258 470614
rect -5814 450378 -5578 450614
rect -5494 450378 -5258 450614
rect -5814 430378 -5578 430614
rect -5494 430378 -5258 430614
rect -5814 410378 -5578 410614
rect -5494 410378 -5258 410614
rect -5814 390378 -5578 390614
rect -5494 390378 -5258 390614
rect -5814 370378 -5578 370614
rect -5494 370378 -5258 370614
rect -5814 350378 -5578 350614
rect -5494 350378 -5258 350614
rect -5814 330378 -5578 330614
rect -5494 330378 -5258 330614
rect -5814 310378 -5578 310614
rect -5494 310378 -5258 310614
rect -5814 290378 -5578 290614
rect -5494 290378 -5258 290614
rect -5814 270378 -5578 270614
rect -5494 270378 -5258 270614
rect -5814 250378 -5578 250614
rect -5494 250378 -5258 250614
rect -5814 230378 -5578 230614
rect -5494 230378 -5258 230614
rect -5814 210378 -5578 210614
rect -5494 210378 -5258 210614
rect -5814 190378 -5578 190614
rect -5494 190378 -5258 190614
rect -5814 170378 -5578 170614
rect -5494 170378 -5258 170614
rect -5814 150378 -5578 150614
rect -5494 150378 -5258 150614
rect -5814 130378 -5578 130614
rect -5494 130378 -5258 130614
rect -5814 110378 -5578 110614
rect -5494 110378 -5258 110614
rect -5814 90378 -5578 90614
rect -5494 90378 -5258 90614
rect -5814 70378 -5578 70614
rect -5494 70378 -5258 70614
rect -5814 50378 -5578 50614
rect -5494 50378 -5258 50614
rect -5814 30378 -5578 30614
rect -5494 30378 -5258 30614
rect -5814 10378 -5578 10614
rect -5494 10378 -5258 10614
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 696718 -4618 696954
rect -4534 696718 -4298 696954
rect -4854 676718 -4618 676954
rect -4534 676718 -4298 676954
rect -4854 656718 -4618 656954
rect -4534 656718 -4298 656954
rect -4854 636718 -4618 636954
rect -4534 636718 -4298 636954
rect -4854 616718 -4618 616954
rect -4534 616718 -4298 616954
rect -4854 596718 -4618 596954
rect -4534 596718 -4298 596954
rect -4854 576718 -4618 576954
rect -4534 576718 -4298 576954
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 536718 -4618 536954
rect -4534 536718 -4298 536954
rect -4854 516718 -4618 516954
rect -4534 516718 -4298 516954
rect -4854 496718 -4618 496954
rect -4534 496718 -4298 496954
rect -4854 476718 -4618 476954
rect -4534 476718 -4298 476954
rect -4854 456718 -4618 456954
rect -4534 456718 -4298 456954
rect -4854 436718 -4618 436954
rect -4534 436718 -4298 436954
rect -4854 416718 -4618 416954
rect -4534 416718 -4298 416954
rect -4854 396718 -4618 396954
rect -4534 396718 -4298 396954
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 356718 -4618 356954
rect -4534 356718 -4298 356954
rect -4854 336718 -4618 336954
rect -4534 336718 -4298 336954
rect -4854 316718 -4618 316954
rect -4534 316718 -4298 316954
rect -4854 296718 -4618 296954
rect -4534 296718 -4298 296954
rect -4854 276718 -4618 276954
rect -4534 276718 -4298 276954
rect -4854 256718 -4618 256954
rect -4534 256718 -4298 256954
rect -4854 236718 -4618 236954
rect -4534 236718 -4298 236954
rect -4854 216718 -4618 216954
rect -4534 216718 -4298 216954
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 176718 -4618 176954
rect -4534 176718 -4298 176954
rect -4854 156718 -4618 156954
rect -4534 156718 -4298 156954
rect -4854 136718 -4618 136954
rect -4534 136718 -4298 136954
rect -4854 116718 -4618 116954
rect -4534 116718 -4298 116954
rect -4854 96718 -4618 96954
rect -4534 96718 -4298 96954
rect -4854 76718 -4618 76954
rect -4534 76718 -4298 76954
rect -4854 56718 -4618 56954
rect -4534 56718 -4298 56954
rect -4854 36718 -4618 36954
rect -4534 36718 -4298 36954
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 686718 -3658 686954
rect -3574 686718 -3338 686954
rect -3894 666718 -3658 666954
rect -3574 666718 -3338 666954
rect -3894 646718 -3658 646954
rect -3574 646718 -3338 646954
rect -3894 626718 -3658 626954
rect -3574 626718 -3338 626954
rect -3894 606718 -3658 606954
rect -3574 606718 -3338 606954
rect -3894 586718 -3658 586954
rect -3574 586718 -3338 586954
rect -3894 566718 -3658 566954
rect -3574 566718 -3338 566954
rect -3894 546718 -3658 546954
rect -3574 546718 -3338 546954
rect -3894 526718 -3658 526954
rect -3574 526718 -3338 526954
rect -3894 506718 -3658 506954
rect -3574 506718 -3338 506954
rect -3894 486718 -3658 486954
rect -3574 486718 -3338 486954
rect -3894 466718 -3658 466954
rect -3574 466718 -3338 466954
rect -3894 446718 -3658 446954
rect -3574 446718 -3338 446954
rect -3894 426718 -3658 426954
rect -3574 426718 -3338 426954
rect -3894 406718 -3658 406954
rect -3574 406718 -3338 406954
rect -3894 386718 -3658 386954
rect -3574 386718 -3338 386954
rect -3894 366718 -3658 366954
rect -3574 366718 -3338 366954
rect -3894 346718 -3658 346954
rect -3574 346718 -3338 346954
rect -3894 326718 -3658 326954
rect -3574 326718 -3338 326954
rect -3894 306718 -3658 306954
rect -3574 306718 -3338 306954
rect -3894 286718 -3658 286954
rect -3574 286718 -3338 286954
rect -3894 266718 -3658 266954
rect -3574 266718 -3338 266954
rect -3894 246718 -3658 246954
rect -3574 246718 -3338 246954
rect -3894 226718 -3658 226954
rect -3574 226718 -3338 226954
rect -3894 206718 -3658 206954
rect -3574 206718 -3338 206954
rect -3894 186718 -3658 186954
rect -3574 186718 -3338 186954
rect -3894 166718 -3658 166954
rect -3574 166718 -3338 166954
rect -3894 146718 -3658 146954
rect -3574 146718 -3338 146954
rect -3894 126718 -3658 126954
rect -3574 126718 -3338 126954
rect -3894 106718 -3658 106954
rect -3574 106718 -3338 106954
rect -3894 86718 -3658 86954
rect -3574 86718 -3338 86954
rect -3894 66718 -3658 66954
rect -3574 66718 -3338 66954
rect -3894 46718 -3658 46954
rect -3574 46718 -3338 46954
rect -3894 26718 -3658 26954
rect -3574 26718 -3338 26954
rect -3894 6718 -3658 6954
rect -3574 6718 -3338 6954
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 693058 -2698 693294
rect -2614 693058 -2378 693294
rect -2934 673058 -2698 673294
rect -2614 673058 -2378 673294
rect -2934 653058 -2698 653294
rect -2614 653058 -2378 653294
rect -2934 633058 -2698 633294
rect -2614 633058 -2378 633294
rect -2934 613058 -2698 613294
rect -2614 613058 -2378 613294
rect -2934 593058 -2698 593294
rect -2614 593058 -2378 593294
rect -2934 573058 -2698 573294
rect -2614 573058 -2378 573294
rect -2934 553058 -2698 553294
rect -2614 553058 -2378 553294
rect -2934 533058 -2698 533294
rect -2614 533058 -2378 533294
rect -2934 513058 -2698 513294
rect -2614 513058 -2378 513294
rect -2934 493058 -2698 493294
rect -2614 493058 -2378 493294
rect -2934 473058 -2698 473294
rect -2614 473058 -2378 473294
rect -2934 453058 -2698 453294
rect -2614 453058 -2378 453294
rect -2934 433058 -2698 433294
rect -2614 433058 -2378 433294
rect -2934 413058 -2698 413294
rect -2614 413058 -2378 413294
rect -2934 393058 -2698 393294
rect -2614 393058 -2378 393294
rect -2934 373058 -2698 373294
rect -2614 373058 -2378 373294
rect -2934 353058 -2698 353294
rect -2614 353058 -2378 353294
rect -2934 333058 -2698 333294
rect -2614 333058 -2378 333294
rect -2934 313058 -2698 313294
rect -2614 313058 -2378 313294
rect -2934 293058 -2698 293294
rect -2614 293058 -2378 293294
rect -2934 273058 -2698 273294
rect -2614 273058 -2378 273294
rect -2934 253058 -2698 253294
rect -2614 253058 -2378 253294
rect -2934 233058 -2698 233294
rect -2614 233058 -2378 233294
rect -2934 213058 -2698 213294
rect -2614 213058 -2378 213294
rect -2934 193058 -2698 193294
rect -2614 193058 -2378 193294
rect -2934 173058 -2698 173294
rect -2614 173058 -2378 173294
rect -2934 153058 -2698 153294
rect -2614 153058 -2378 153294
rect -2934 133058 -2698 133294
rect -2614 133058 -2378 133294
rect -2934 113058 -2698 113294
rect -2614 113058 -2378 113294
rect -2934 93058 -2698 93294
rect -2614 93058 -2378 93294
rect -2934 73058 -2698 73294
rect -2614 73058 -2378 73294
rect -2934 53058 -2698 53294
rect -2614 53058 -2378 53294
rect -2934 33058 -2698 33294
rect -2614 33058 -2378 33294
rect -2934 13058 -2698 13294
rect -2614 13058 -2378 13294
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 683058 -1738 683294
rect -1654 683058 -1418 683294
rect -1974 663058 -1738 663294
rect -1654 663058 -1418 663294
rect -1974 643058 -1738 643294
rect -1654 643058 -1418 643294
rect -1974 623058 -1738 623294
rect -1654 623058 -1418 623294
rect -1974 603058 -1738 603294
rect -1654 603058 -1418 603294
rect -1974 583058 -1738 583294
rect -1654 583058 -1418 583294
rect -1974 563058 -1738 563294
rect -1654 563058 -1418 563294
rect -1974 543058 -1738 543294
rect -1654 543058 -1418 543294
rect -1974 523058 -1738 523294
rect -1654 523058 -1418 523294
rect -1974 503058 -1738 503294
rect -1654 503058 -1418 503294
rect -1974 483058 -1738 483294
rect -1654 483058 -1418 483294
rect -1974 463058 -1738 463294
rect -1654 463058 -1418 463294
rect -1974 443058 -1738 443294
rect -1654 443058 -1418 443294
rect -1974 423058 -1738 423294
rect -1654 423058 -1418 423294
rect -1974 403058 -1738 403294
rect -1654 403058 -1418 403294
rect -1974 383058 -1738 383294
rect -1654 383058 -1418 383294
rect -1974 363058 -1738 363294
rect -1654 363058 -1418 363294
rect -1974 343058 -1738 343294
rect -1654 343058 -1418 343294
rect -1974 323058 -1738 323294
rect -1654 323058 -1418 323294
rect -1974 303058 -1738 303294
rect -1654 303058 -1418 303294
rect -1974 283058 -1738 283294
rect -1654 283058 -1418 283294
rect -1974 263058 -1738 263294
rect -1654 263058 -1418 263294
rect -1974 243058 -1738 243294
rect -1654 243058 -1418 243294
rect -1974 223058 -1738 223294
rect -1654 223058 -1418 223294
rect -1974 203058 -1738 203294
rect -1654 203058 -1418 203294
rect -1974 183058 -1738 183294
rect -1654 183058 -1418 183294
rect -1974 163058 -1738 163294
rect -1654 163058 -1418 163294
rect -1974 143058 -1738 143294
rect -1654 143058 -1418 143294
rect -1974 123058 -1738 123294
rect -1654 123058 -1418 123294
rect -1974 103058 -1738 103294
rect -1654 103058 -1418 103294
rect -1974 83058 -1738 83294
rect -1654 83058 -1418 83294
rect -1974 63058 -1738 63294
rect -1654 63058 -1418 63294
rect -1974 43058 -1738 43294
rect -1654 43058 -1418 43294
rect -1974 23058 -1738 23294
rect -1654 23058 -1418 23294
rect -1974 3058 -1738 3294
rect -1654 3058 -1418 3294
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 683058 2062 683294
rect 2146 683058 2382 683294
rect 1826 663058 2062 663294
rect 2146 663058 2382 663294
rect 1826 643058 2062 643294
rect 2146 643058 2382 643294
rect 1826 623058 2062 623294
rect 2146 623058 2382 623294
rect 1826 603058 2062 603294
rect 2146 603058 2382 603294
rect 1826 583058 2062 583294
rect 2146 583058 2382 583294
rect 1826 563058 2062 563294
rect 2146 563058 2382 563294
rect 1826 543058 2062 543294
rect 2146 543058 2382 543294
rect 1826 523058 2062 523294
rect 2146 523058 2382 523294
rect 1826 503058 2062 503294
rect 2146 503058 2382 503294
rect 1826 483058 2062 483294
rect 2146 483058 2382 483294
rect 1826 463058 2062 463294
rect 2146 463058 2382 463294
rect 1826 443058 2062 443294
rect 2146 443058 2382 443294
rect 1826 423058 2062 423294
rect 2146 423058 2382 423294
rect 1826 403058 2062 403294
rect 2146 403058 2382 403294
rect 1826 383058 2062 383294
rect 2146 383058 2382 383294
rect 1826 363058 2062 363294
rect 2146 363058 2382 363294
rect 1826 343058 2062 343294
rect 2146 343058 2382 343294
rect 1826 323058 2062 323294
rect 2146 323058 2382 323294
rect 1826 303058 2062 303294
rect 2146 303058 2382 303294
rect 1826 283058 2062 283294
rect 2146 283058 2382 283294
rect 1826 263058 2062 263294
rect 2146 263058 2382 263294
rect 1826 243058 2062 243294
rect 2146 243058 2382 243294
rect 1826 223058 2062 223294
rect 2146 223058 2382 223294
rect 1826 203058 2062 203294
rect 2146 203058 2382 203294
rect 1826 183058 2062 183294
rect 2146 183058 2382 183294
rect 1826 163058 2062 163294
rect 2146 163058 2382 163294
rect 1826 143058 2062 143294
rect 2146 143058 2382 143294
rect 1826 123058 2062 123294
rect 2146 123058 2382 123294
rect 1826 103058 2062 103294
rect 2146 103058 2382 103294
rect 1826 83058 2062 83294
rect 2146 83058 2382 83294
rect 1826 63058 2062 63294
rect 2146 63058 2382 63294
rect 1826 43058 2062 43294
rect 2146 43058 2382 43294
rect 1826 23058 2062 23294
rect 2146 23058 2382 23294
rect 1826 3058 2062 3294
rect 2146 3058 2382 3294
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 686718 5782 686954
rect 5866 686718 6102 686954
rect 5546 666718 5782 666954
rect 5866 666718 6102 666954
rect 5546 646718 5782 646954
rect 5866 646718 6102 646954
rect 5546 626718 5782 626954
rect 5866 626718 6102 626954
rect 5546 606718 5782 606954
rect 5866 606718 6102 606954
rect 5546 586718 5782 586954
rect 5866 586718 6102 586954
rect 5546 566718 5782 566954
rect 5866 566718 6102 566954
rect 5546 546718 5782 546954
rect 5866 546718 6102 546954
rect 5546 526718 5782 526954
rect 5866 526718 6102 526954
rect 5546 506718 5782 506954
rect 5866 506718 6102 506954
rect 5546 486718 5782 486954
rect 5866 486718 6102 486954
rect 5546 466718 5782 466954
rect 5866 466718 6102 466954
rect 5546 446718 5782 446954
rect 5866 446718 6102 446954
rect 5546 426718 5782 426954
rect 5866 426718 6102 426954
rect 5546 406718 5782 406954
rect 5866 406718 6102 406954
rect 5546 386718 5782 386954
rect 5866 386718 6102 386954
rect 5546 366718 5782 366954
rect 5866 366718 6102 366954
rect 5546 346718 5782 346954
rect 5866 346718 6102 346954
rect 5546 326718 5782 326954
rect 5866 326718 6102 326954
rect 5546 306718 5782 306954
rect 5866 306718 6102 306954
rect 5546 286718 5782 286954
rect 5866 286718 6102 286954
rect 5546 266718 5782 266954
rect 5866 266718 6102 266954
rect 5546 246718 5782 246954
rect 5866 246718 6102 246954
rect 5546 226718 5782 226954
rect 5866 226718 6102 226954
rect 5546 206718 5782 206954
rect 5866 206718 6102 206954
rect 5546 186718 5782 186954
rect 5866 186718 6102 186954
rect 5546 166718 5782 166954
rect 5866 166718 6102 166954
rect 5546 146718 5782 146954
rect 5866 146718 6102 146954
rect 5546 126718 5782 126954
rect 5866 126718 6102 126954
rect 5546 106718 5782 106954
rect 5866 106718 6102 106954
rect 5546 86718 5782 86954
rect 5866 86718 6102 86954
rect 5546 66718 5782 66954
rect 5866 66718 6102 66954
rect 5546 46718 5782 46954
rect 5866 46718 6102 46954
rect 5546 26718 5782 26954
rect 5866 26718 6102 26954
rect 5546 6718 5782 6954
rect 5866 6718 6102 6954
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 690378 9502 690614
rect 9586 690378 9822 690614
rect 9266 670378 9502 670614
rect 9586 670378 9822 670614
rect 9266 650378 9502 650614
rect 9586 650378 9822 650614
rect 9266 630378 9502 630614
rect 9586 630378 9822 630614
rect 9266 610378 9502 610614
rect 9586 610378 9822 610614
rect 9266 590378 9502 590614
rect 9586 590378 9822 590614
rect 9266 570378 9502 570614
rect 9586 570378 9822 570614
rect 9266 550378 9502 550614
rect 9586 550378 9822 550614
rect 9266 530378 9502 530614
rect 9586 530378 9822 530614
rect 9266 510378 9502 510614
rect 9586 510378 9822 510614
rect 9266 490378 9502 490614
rect 9586 490378 9822 490614
rect 9266 470378 9502 470614
rect 9586 470378 9822 470614
rect 9266 450378 9502 450614
rect 9586 450378 9822 450614
rect 9266 430378 9502 430614
rect 9586 430378 9822 430614
rect 9266 410378 9502 410614
rect 9586 410378 9822 410614
rect 9266 390378 9502 390614
rect 9586 390378 9822 390614
rect 9266 370378 9502 370614
rect 9586 370378 9822 370614
rect 9266 350378 9502 350614
rect 9586 350378 9822 350614
rect 9266 330378 9502 330614
rect 9586 330378 9822 330614
rect 9266 310378 9502 310614
rect 9586 310378 9822 310614
rect 9266 290378 9502 290614
rect 9586 290378 9822 290614
rect 9266 270378 9502 270614
rect 9586 270378 9822 270614
rect 9266 250378 9502 250614
rect 9586 250378 9822 250614
rect 9266 230378 9502 230614
rect 9586 230378 9822 230614
rect 9266 210378 9502 210614
rect 9586 210378 9822 210614
rect 9266 190378 9502 190614
rect 9586 190378 9822 190614
rect 9266 170378 9502 170614
rect 9586 170378 9822 170614
rect 9266 150378 9502 150614
rect 9586 150378 9822 150614
rect 9266 130378 9502 130614
rect 9586 130378 9822 130614
rect 9266 110378 9502 110614
rect 9586 110378 9822 110614
rect 9266 90378 9502 90614
rect 9586 90378 9822 90614
rect 9266 70378 9502 70614
rect 9586 70378 9822 70614
rect 9266 50378 9502 50614
rect 9586 50378 9822 50614
rect 9266 30378 9502 30614
rect 9586 30378 9822 30614
rect 9266 10378 9502 10614
rect 9586 10378 9822 10614
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 11826 705562 12062 705798
rect 12146 705562 12382 705798
rect 11826 705242 12062 705478
rect 12146 705242 12382 705478
rect 11826 693058 12062 693294
rect 12146 693058 12382 693294
rect 11826 673058 12062 673294
rect 12146 673058 12382 673294
rect 11826 653058 12062 653294
rect 12146 653058 12382 653294
rect 11826 633058 12062 633294
rect 12146 633058 12382 633294
rect 11826 613058 12062 613294
rect 12146 613058 12382 613294
rect 11826 593058 12062 593294
rect 12146 593058 12382 593294
rect 11826 573058 12062 573294
rect 12146 573058 12382 573294
rect 11826 553058 12062 553294
rect 12146 553058 12382 553294
rect 11826 533058 12062 533294
rect 12146 533058 12382 533294
rect 11826 513058 12062 513294
rect 12146 513058 12382 513294
rect 11826 493058 12062 493294
rect 12146 493058 12382 493294
rect 11826 473058 12062 473294
rect 12146 473058 12382 473294
rect 11826 453058 12062 453294
rect 12146 453058 12382 453294
rect 11826 433058 12062 433294
rect 12146 433058 12382 433294
rect 11826 413058 12062 413294
rect 12146 413058 12382 413294
rect 11826 393058 12062 393294
rect 12146 393058 12382 393294
rect 11826 373058 12062 373294
rect 12146 373058 12382 373294
rect 11826 353058 12062 353294
rect 12146 353058 12382 353294
rect 11826 333058 12062 333294
rect 12146 333058 12382 333294
rect 11826 313058 12062 313294
rect 12146 313058 12382 313294
rect 11826 293058 12062 293294
rect 12146 293058 12382 293294
rect 11826 273058 12062 273294
rect 12146 273058 12382 273294
rect 11826 253058 12062 253294
rect 12146 253058 12382 253294
rect 11826 233058 12062 233294
rect 12146 233058 12382 233294
rect 11826 213058 12062 213294
rect 12146 213058 12382 213294
rect 11826 193058 12062 193294
rect 12146 193058 12382 193294
rect 11826 173058 12062 173294
rect 12146 173058 12382 173294
rect 11826 153058 12062 153294
rect 12146 153058 12382 153294
rect 11826 133058 12062 133294
rect 12146 133058 12382 133294
rect 11826 113058 12062 113294
rect 12146 113058 12382 113294
rect 11826 93058 12062 93294
rect 12146 93058 12382 93294
rect 11826 73058 12062 73294
rect 12146 73058 12382 73294
rect 11826 53058 12062 53294
rect 12146 53058 12382 53294
rect 11826 33058 12062 33294
rect 12146 33058 12382 33294
rect 11826 13058 12062 13294
rect 12146 13058 12382 13294
rect 11826 -1542 12062 -1306
rect 12146 -1542 12382 -1306
rect 11826 -1862 12062 -1626
rect 12146 -1862 12382 -1626
rect 22986 711322 23222 711558
rect 23306 711322 23542 711558
rect 22986 711002 23222 711238
rect 23306 711002 23542 711238
rect 19266 709402 19502 709638
rect 19586 709402 19822 709638
rect 19266 709082 19502 709318
rect 19586 709082 19822 709318
rect 12986 694038 13222 694274
rect 13306 694038 13542 694274
rect 12986 674038 13222 674274
rect 13306 674038 13542 674274
rect 12986 654038 13222 654274
rect 13306 654038 13542 654274
rect 12986 634038 13222 634274
rect 13306 634038 13542 634274
rect 12986 614038 13222 614274
rect 13306 614038 13542 614274
rect 12986 594038 13222 594274
rect 13306 594038 13542 594274
rect 12986 574038 13222 574274
rect 13306 574038 13542 574274
rect 12986 554038 13222 554274
rect 13306 554038 13542 554274
rect 12986 534038 13222 534274
rect 13306 534038 13542 534274
rect 12986 514038 13222 514274
rect 13306 514038 13542 514274
rect 12986 494038 13222 494274
rect 13306 494038 13542 494274
rect 12986 474038 13222 474274
rect 13306 474038 13542 474274
rect 12986 454038 13222 454274
rect 13306 454038 13542 454274
rect 12986 434038 13222 434274
rect 13306 434038 13542 434274
rect 12986 414038 13222 414274
rect 13306 414038 13542 414274
rect 12986 394038 13222 394274
rect 13306 394038 13542 394274
rect 12986 374038 13222 374274
rect 13306 374038 13542 374274
rect 12986 354038 13222 354274
rect 13306 354038 13542 354274
rect 12986 334038 13222 334274
rect 13306 334038 13542 334274
rect 12986 314038 13222 314274
rect 13306 314038 13542 314274
rect 12986 294038 13222 294274
rect 13306 294038 13542 294274
rect 12986 274038 13222 274274
rect 13306 274038 13542 274274
rect 12986 254038 13222 254274
rect 13306 254038 13542 254274
rect 12986 234038 13222 234274
rect 13306 234038 13542 234274
rect 12986 214038 13222 214274
rect 13306 214038 13542 214274
rect 12986 194038 13222 194274
rect 13306 194038 13542 194274
rect 12986 174038 13222 174274
rect 13306 174038 13542 174274
rect 12986 154038 13222 154274
rect 13306 154038 13542 154274
rect 12986 134038 13222 134274
rect 13306 134038 13542 134274
rect 12986 114038 13222 114274
rect 13306 114038 13542 114274
rect 12986 94038 13222 94274
rect 13306 94038 13542 94274
rect 12986 74038 13222 74274
rect 13306 74038 13542 74274
rect 12986 54038 13222 54274
rect 13306 54038 13542 54274
rect 12986 34038 13222 34274
rect 13306 34038 13542 34274
rect 12986 14038 13222 14274
rect 13306 14038 13542 14274
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 15546 707482 15782 707718
rect 15866 707482 16102 707718
rect 15546 707162 15782 707398
rect 15866 707162 16102 707398
rect 15546 696718 15782 696954
rect 15866 696718 16102 696954
rect 15546 676718 15782 676954
rect 15866 676718 16102 676954
rect 15546 656718 15782 656954
rect 15866 656718 16102 656954
rect 15546 636718 15782 636954
rect 15866 636718 16102 636954
rect 15546 616718 15782 616954
rect 15866 616718 16102 616954
rect 15546 596718 15782 596954
rect 15866 596718 16102 596954
rect 15546 576718 15782 576954
rect 15866 576718 16102 576954
rect 15546 556718 15782 556954
rect 15866 556718 16102 556954
rect 15546 536718 15782 536954
rect 15866 536718 16102 536954
rect 15546 516718 15782 516954
rect 15866 516718 16102 516954
rect 15546 496718 15782 496954
rect 15866 496718 16102 496954
rect 15546 476718 15782 476954
rect 15866 476718 16102 476954
rect 15546 456718 15782 456954
rect 15866 456718 16102 456954
rect 15546 436718 15782 436954
rect 15866 436718 16102 436954
rect 15546 416718 15782 416954
rect 15866 416718 16102 416954
rect 15546 396718 15782 396954
rect 15866 396718 16102 396954
rect 15546 376718 15782 376954
rect 15866 376718 16102 376954
rect 15546 356718 15782 356954
rect 15866 356718 16102 356954
rect 15546 336718 15782 336954
rect 15866 336718 16102 336954
rect 15546 316718 15782 316954
rect 15866 316718 16102 316954
rect 15546 296718 15782 296954
rect 15866 296718 16102 296954
rect 15546 276718 15782 276954
rect 15866 276718 16102 276954
rect 15546 256718 15782 256954
rect 15866 256718 16102 256954
rect 15546 236718 15782 236954
rect 15866 236718 16102 236954
rect 15546 216718 15782 216954
rect 15866 216718 16102 216954
rect 15546 196718 15782 196954
rect 15866 196718 16102 196954
rect 15546 176718 15782 176954
rect 15866 176718 16102 176954
rect 15546 156718 15782 156954
rect 15866 156718 16102 156954
rect 15546 136718 15782 136954
rect 15866 136718 16102 136954
rect 15546 116718 15782 116954
rect 15866 116718 16102 116954
rect 15546 96718 15782 96954
rect 15866 96718 16102 96954
rect 15546 76718 15782 76954
rect 15866 76718 16102 76954
rect 15546 56718 15782 56954
rect 15866 56718 16102 56954
rect 15546 36718 15782 36954
rect 15866 36718 16102 36954
rect 15546 16718 15782 16954
rect 15866 16718 16102 16954
rect 15546 -3462 15782 -3226
rect 15866 -3462 16102 -3226
rect 15546 -3782 15782 -3546
rect 15866 -3782 16102 -3546
rect 19266 700378 19502 700614
rect 19586 700378 19822 700614
rect 19266 680378 19502 680614
rect 19586 680378 19822 680614
rect 19266 660378 19502 660614
rect 19586 660378 19822 660614
rect 19266 640378 19502 640614
rect 19586 640378 19822 640614
rect 19266 620378 19502 620614
rect 19586 620378 19822 620614
rect 19266 600378 19502 600614
rect 19586 600378 19822 600614
rect 19266 580378 19502 580614
rect 19586 580378 19822 580614
rect 19266 560378 19502 560614
rect 19586 560378 19822 560614
rect 19266 540378 19502 540614
rect 19586 540378 19822 540614
rect 19266 520378 19502 520614
rect 19586 520378 19822 520614
rect 19266 500378 19502 500614
rect 19586 500378 19822 500614
rect 19266 480378 19502 480614
rect 19586 480378 19822 480614
rect 19266 460378 19502 460614
rect 19586 460378 19822 460614
rect 19266 440378 19502 440614
rect 19586 440378 19822 440614
rect 19266 420378 19502 420614
rect 19586 420378 19822 420614
rect 19266 400378 19502 400614
rect 19586 400378 19822 400614
rect 19266 380378 19502 380614
rect 19586 380378 19822 380614
rect 19266 360378 19502 360614
rect 19586 360378 19822 360614
rect 19266 340378 19502 340614
rect 19586 340378 19822 340614
rect 19266 320378 19502 320614
rect 19586 320378 19822 320614
rect 19266 300378 19502 300614
rect 19586 300378 19822 300614
rect 19266 280378 19502 280614
rect 19586 280378 19822 280614
rect 19266 260378 19502 260614
rect 19586 260378 19822 260614
rect 19266 240378 19502 240614
rect 19586 240378 19822 240614
rect 19266 220378 19502 220614
rect 19586 220378 19822 220614
rect 19266 200378 19502 200614
rect 19586 200378 19822 200614
rect 19266 180378 19502 180614
rect 19586 180378 19822 180614
rect 19266 160378 19502 160614
rect 19586 160378 19822 160614
rect 19266 140378 19502 140614
rect 19586 140378 19822 140614
rect 19266 120378 19502 120614
rect 19586 120378 19822 120614
rect 19266 100378 19502 100614
rect 19586 100378 19822 100614
rect 19266 80378 19502 80614
rect 19586 80378 19822 80614
rect 19266 60378 19502 60614
rect 19586 60378 19822 60614
rect 19266 40378 19502 40614
rect 19586 40378 19822 40614
rect 19266 20378 19502 20614
rect 19586 20378 19822 20614
rect 21826 704602 22062 704838
rect 22146 704602 22382 704838
rect 21826 704282 22062 704518
rect 22146 704282 22382 704518
rect 21826 683058 22062 683294
rect 22146 683058 22382 683294
rect 21826 663058 22062 663294
rect 22146 663058 22382 663294
rect 21826 643058 22062 643294
rect 22146 643058 22382 643294
rect 21826 623058 22062 623294
rect 22146 623058 22382 623294
rect 21826 603058 22062 603294
rect 22146 603058 22382 603294
rect 21826 583058 22062 583294
rect 22146 583058 22382 583294
rect 21826 563058 22062 563294
rect 22146 563058 22382 563294
rect 21826 543058 22062 543294
rect 22146 543058 22382 543294
rect 21826 523058 22062 523294
rect 22146 523058 22382 523294
rect 21826 503058 22062 503294
rect 22146 503058 22382 503294
rect 21826 483058 22062 483294
rect 22146 483058 22382 483294
rect 21826 463058 22062 463294
rect 22146 463058 22382 463294
rect 21826 443058 22062 443294
rect 22146 443058 22382 443294
rect 21826 423058 22062 423294
rect 22146 423058 22382 423294
rect 21826 403058 22062 403294
rect 22146 403058 22382 403294
rect 21826 383058 22062 383294
rect 22146 383058 22382 383294
rect 21826 363058 22062 363294
rect 22146 363058 22382 363294
rect 21826 343058 22062 343294
rect 22146 343058 22382 343294
rect 21826 323058 22062 323294
rect 22146 323058 22382 323294
rect 21826 303058 22062 303294
rect 22146 303058 22382 303294
rect 21826 283058 22062 283294
rect 22146 283058 22382 283294
rect 21826 263058 22062 263294
rect 22146 263058 22382 263294
rect 21826 243058 22062 243294
rect 22146 243058 22382 243294
rect 21826 223058 22062 223294
rect 22146 223058 22382 223294
rect 21826 203058 22062 203294
rect 22146 203058 22382 203294
rect 21826 183058 22062 183294
rect 22146 183058 22382 183294
rect 21826 163058 22062 163294
rect 22146 163058 22382 163294
rect 21826 143058 22062 143294
rect 22146 143058 22382 143294
rect 21826 123058 22062 123294
rect 22146 123058 22382 123294
rect 21826 103058 22062 103294
rect 22146 103058 22382 103294
rect 21826 83058 22062 83294
rect 22146 83058 22382 83294
rect 21826 63058 22062 63294
rect 22146 63058 22382 63294
rect 21826 43058 22062 43294
rect 22146 43058 22382 43294
rect 21826 23058 22062 23294
rect 22146 23058 22382 23294
rect 21826 3058 22062 3294
rect 22146 3058 22382 3294
rect 21826 -582 22062 -346
rect 22146 -582 22382 -346
rect 21826 -902 22062 -666
rect 22146 -902 22382 -666
rect 32986 710362 33222 710598
rect 33306 710362 33542 710598
rect 32986 710042 33222 710278
rect 33306 710042 33542 710278
rect 29266 708442 29502 708678
rect 29586 708442 29822 708678
rect 29266 708122 29502 708358
rect 29586 708122 29822 708358
rect 22986 684038 23222 684274
rect 23306 684038 23542 684274
rect 22986 664038 23222 664274
rect 23306 664038 23542 664274
rect 22986 644038 23222 644274
rect 23306 644038 23542 644274
rect 22986 624038 23222 624274
rect 23306 624038 23542 624274
rect 22986 604038 23222 604274
rect 23306 604038 23542 604274
rect 22986 584038 23222 584274
rect 23306 584038 23542 584274
rect 22986 564038 23222 564274
rect 23306 564038 23542 564274
rect 22986 544038 23222 544274
rect 23306 544038 23542 544274
rect 22986 524038 23222 524274
rect 23306 524038 23542 524274
rect 22986 504038 23222 504274
rect 23306 504038 23542 504274
rect 22986 484038 23222 484274
rect 23306 484038 23542 484274
rect 22986 464038 23222 464274
rect 23306 464038 23542 464274
rect 22986 444038 23222 444274
rect 23306 444038 23542 444274
rect 22986 424038 23222 424274
rect 23306 424038 23542 424274
rect 22986 404038 23222 404274
rect 23306 404038 23542 404274
rect 22986 384038 23222 384274
rect 23306 384038 23542 384274
rect 22986 364038 23222 364274
rect 23306 364038 23542 364274
rect 22986 344038 23222 344274
rect 23306 344038 23542 344274
rect 22986 324038 23222 324274
rect 23306 324038 23542 324274
rect 22986 304038 23222 304274
rect 23306 304038 23542 304274
rect 22986 284038 23222 284274
rect 23306 284038 23542 284274
rect 22986 264038 23222 264274
rect 23306 264038 23542 264274
rect 22986 244038 23222 244274
rect 23306 244038 23542 244274
rect 22986 224038 23222 224274
rect 23306 224038 23542 224274
rect 22986 204038 23222 204274
rect 23306 204038 23542 204274
rect 22986 184038 23222 184274
rect 23306 184038 23542 184274
rect 22986 164038 23222 164274
rect 23306 164038 23542 164274
rect 22986 144038 23222 144274
rect 23306 144038 23542 144274
rect 22986 124038 23222 124274
rect 23306 124038 23542 124274
rect 22986 104038 23222 104274
rect 23306 104038 23542 104274
rect 22986 84038 23222 84274
rect 23306 84038 23542 84274
rect 22986 64038 23222 64274
rect 23306 64038 23542 64274
rect 22986 44038 23222 44274
rect 23306 44038 23542 44274
rect 22986 24038 23222 24274
rect 23306 24038 23542 24274
rect 19266 -5382 19502 -5146
rect 19586 -5382 19822 -5146
rect 19266 -5702 19502 -5466
rect 19586 -5702 19822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 25546 706522 25782 706758
rect 25866 706522 26102 706758
rect 25546 706202 25782 706438
rect 25866 706202 26102 706438
rect 25546 686718 25782 686954
rect 25866 686718 26102 686954
rect 29266 690378 29502 690614
rect 29586 690378 29822 690614
rect 31826 705562 32062 705798
rect 32146 705562 32382 705798
rect 31826 705242 32062 705478
rect 32146 705242 32382 705478
rect 31826 693058 32062 693294
rect 32146 693058 32382 693294
rect 42986 711322 43222 711558
rect 43306 711322 43542 711558
rect 42986 711002 43222 711238
rect 43306 711002 43542 711238
rect 39266 709402 39502 709638
rect 39586 709402 39822 709638
rect 39266 709082 39502 709318
rect 39586 709082 39822 709318
rect 32986 694038 33222 694274
rect 33306 694038 33542 694274
rect 35546 707482 35782 707718
rect 35866 707482 36102 707718
rect 35546 707162 35782 707398
rect 35866 707162 36102 707398
rect 35546 696718 35782 696954
rect 35866 696718 36102 696954
rect 35546 676718 35782 676954
rect 35866 676718 36102 676954
rect 39266 700378 39502 700614
rect 39586 700378 39822 700614
rect 39266 680378 39502 680614
rect 39586 680378 39822 680614
rect 41826 704602 42062 704838
rect 42146 704602 42382 704838
rect 41826 704282 42062 704518
rect 42146 704282 42382 704518
rect 41826 683058 42062 683294
rect 42146 683058 42382 683294
rect 52986 710362 53222 710598
rect 53306 710362 53542 710598
rect 52986 710042 53222 710278
rect 53306 710042 53542 710278
rect 49266 708442 49502 708678
rect 49586 708442 49822 708678
rect 49266 708122 49502 708358
rect 49586 708122 49822 708358
rect 42986 684038 43222 684274
rect 43306 684038 43542 684274
rect 45546 706522 45782 706758
rect 45866 706522 46102 706758
rect 45546 706202 45782 706438
rect 45866 706202 46102 706438
rect 45546 686718 45782 686954
rect 45866 686718 46102 686954
rect 49266 690378 49502 690614
rect 49586 690378 49822 690614
rect 51826 705562 52062 705798
rect 52146 705562 52382 705798
rect 51826 705242 52062 705478
rect 52146 705242 52382 705478
rect 51826 693058 52062 693294
rect 52146 693058 52382 693294
rect 62986 711322 63222 711558
rect 63306 711322 63542 711558
rect 62986 711002 63222 711238
rect 63306 711002 63542 711238
rect 59266 709402 59502 709638
rect 59586 709402 59822 709638
rect 59266 709082 59502 709318
rect 59586 709082 59822 709318
rect 52986 694038 53222 694274
rect 53306 694038 53542 694274
rect 55546 707482 55782 707718
rect 55866 707482 56102 707718
rect 55546 707162 55782 707398
rect 55866 707162 56102 707398
rect 55546 696718 55782 696954
rect 55866 696718 56102 696954
rect 55546 676718 55782 676954
rect 55866 676718 56102 676954
rect 59266 700378 59502 700614
rect 59586 700378 59822 700614
rect 59266 680378 59502 680614
rect 59586 680378 59822 680614
rect 61826 704602 62062 704838
rect 62146 704602 62382 704838
rect 61826 704282 62062 704518
rect 62146 704282 62382 704518
rect 61826 683058 62062 683294
rect 62146 683058 62382 683294
rect 72986 710362 73222 710598
rect 73306 710362 73542 710598
rect 72986 710042 73222 710278
rect 73306 710042 73542 710278
rect 69266 708442 69502 708678
rect 69586 708442 69822 708678
rect 69266 708122 69502 708358
rect 69586 708122 69822 708358
rect 62986 684038 63222 684274
rect 63306 684038 63542 684274
rect 65546 706522 65782 706758
rect 65866 706522 66102 706758
rect 65546 706202 65782 706438
rect 65866 706202 66102 706438
rect 65546 686718 65782 686954
rect 65866 686718 66102 686954
rect 69266 690378 69502 690614
rect 69586 690378 69822 690614
rect 71826 705562 72062 705798
rect 72146 705562 72382 705798
rect 71826 705242 72062 705478
rect 72146 705242 72382 705478
rect 71826 693058 72062 693294
rect 72146 693058 72382 693294
rect 82986 711322 83222 711558
rect 83306 711322 83542 711558
rect 82986 711002 83222 711238
rect 83306 711002 83542 711238
rect 79266 709402 79502 709638
rect 79586 709402 79822 709638
rect 79266 709082 79502 709318
rect 79586 709082 79822 709318
rect 72986 694038 73222 694274
rect 73306 694038 73542 694274
rect 75546 707482 75782 707718
rect 75866 707482 76102 707718
rect 75546 707162 75782 707398
rect 75866 707162 76102 707398
rect 75546 696718 75782 696954
rect 75866 696718 76102 696954
rect 75546 676718 75782 676954
rect 75866 676718 76102 676954
rect 79266 700378 79502 700614
rect 79586 700378 79822 700614
rect 79266 680378 79502 680614
rect 79586 680378 79822 680614
rect 81826 704602 82062 704838
rect 82146 704602 82382 704838
rect 81826 704282 82062 704518
rect 82146 704282 82382 704518
rect 81826 683058 82062 683294
rect 82146 683058 82382 683294
rect 92986 710362 93222 710598
rect 93306 710362 93542 710598
rect 92986 710042 93222 710278
rect 93306 710042 93542 710278
rect 89266 708442 89502 708678
rect 89586 708442 89822 708678
rect 89266 708122 89502 708358
rect 89586 708122 89822 708358
rect 82986 684038 83222 684274
rect 83306 684038 83542 684274
rect 85546 706522 85782 706758
rect 85866 706522 86102 706758
rect 85546 706202 85782 706438
rect 85866 706202 86102 706438
rect 85546 686718 85782 686954
rect 85866 686718 86102 686954
rect 89266 690378 89502 690614
rect 89586 690378 89822 690614
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 693058 92062 693294
rect 92146 693058 92382 693294
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 92986 694038 93222 694274
rect 93306 694038 93542 694274
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 95546 696718 95782 696954
rect 95866 696718 96102 696954
rect 95546 676718 95782 676954
rect 95866 676718 96102 676954
rect 99266 700378 99502 700614
rect 99586 700378 99822 700614
rect 99266 680378 99502 680614
rect 99586 680378 99822 680614
rect 101826 704602 102062 704838
rect 102146 704602 102382 704838
rect 101826 704282 102062 704518
rect 102146 704282 102382 704518
rect 101826 683058 102062 683294
rect 102146 683058 102382 683294
rect 112986 710362 113222 710598
rect 113306 710362 113542 710598
rect 112986 710042 113222 710278
rect 113306 710042 113542 710278
rect 109266 708442 109502 708678
rect 109586 708442 109822 708678
rect 109266 708122 109502 708358
rect 109586 708122 109822 708358
rect 102986 684038 103222 684274
rect 103306 684038 103542 684274
rect 105546 706522 105782 706758
rect 105866 706522 106102 706758
rect 105546 706202 105782 706438
rect 105866 706202 106102 706438
rect 105546 686718 105782 686954
rect 105866 686718 106102 686954
rect 109266 690378 109502 690614
rect 109586 690378 109822 690614
rect 111826 705562 112062 705798
rect 112146 705562 112382 705798
rect 111826 705242 112062 705478
rect 112146 705242 112382 705478
rect 111826 693058 112062 693294
rect 112146 693058 112382 693294
rect 122986 711322 123222 711558
rect 123306 711322 123542 711558
rect 122986 711002 123222 711238
rect 123306 711002 123542 711238
rect 119266 709402 119502 709638
rect 119586 709402 119822 709638
rect 119266 709082 119502 709318
rect 119586 709082 119822 709318
rect 112986 694038 113222 694274
rect 113306 694038 113542 694274
rect 115546 707482 115782 707718
rect 115866 707482 116102 707718
rect 115546 707162 115782 707398
rect 115866 707162 116102 707398
rect 115546 696718 115782 696954
rect 115866 696718 116102 696954
rect 115546 676718 115782 676954
rect 115866 676718 116102 676954
rect 119266 700378 119502 700614
rect 119586 700378 119822 700614
rect 119266 680378 119502 680614
rect 119586 680378 119822 680614
rect 121826 704602 122062 704838
rect 122146 704602 122382 704838
rect 121826 704282 122062 704518
rect 122146 704282 122382 704518
rect 121826 683058 122062 683294
rect 122146 683058 122382 683294
rect 132986 710362 133222 710598
rect 133306 710362 133542 710598
rect 132986 710042 133222 710278
rect 133306 710042 133542 710278
rect 129266 708442 129502 708678
rect 129586 708442 129822 708678
rect 129266 708122 129502 708358
rect 129586 708122 129822 708358
rect 122986 684038 123222 684274
rect 123306 684038 123542 684274
rect 125546 706522 125782 706758
rect 125866 706522 126102 706758
rect 125546 706202 125782 706438
rect 125866 706202 126102 706438
rect 125546 686718 125782 686954
rect 125866 686718 126102 686954
rect 129266 690378 129502 690614
rect 129586 690378 129822 690614
rect 131826 705562 132062 705798
rect 132146 705562 132382 705798
rect 131826 705242 132062 705478
rect 132146 705242 132382 705478
rect 131826 693058 132062 693294
rect 132146 693058 132382 693294
rect 142986 711322 143222 711558
rect 143306 711322 143542 711558
rect 142986 711002 143222 711238
rect 143306 711002 143542 711238
rect 139266 709402 139502 709638
rect 139586 709402 139822 709638
rect 139266 709082 139502 709318
rect 139586 709082 139822 709318
rect 132986 694038 133222 694274
rect 133306 694038 133542 694274
rect 135546 707482 135782 707718
rect 135866 707482 136102 707718
rect 135546 707162 135782 707398
rect 135866 707162 136102 707398
rect 135546 696718 135782 696954
rect 135866 696718 136102 696954
rect 135546 676718 135782 676954
rect 135866 676718 136102 676954
rect 139266 700378 139502 700614
rect 139586 700378 139822 700614
rect 139266 680378 139502 680614
rect 139586 680378 139822 680614
rect 141826 704602 142062 704838
rect 142146 704602 142382 704838
rect 141826 704282 142062 704518
rect 142146 704282 142382 704518
rect 141826 683058 142062 683294
rect 142146 683058 142382 683294
rect 152986 710362 153222 710598
rect 153306 710362 153542 710598
rect 152986 710042 153222 710278
rect 153306 710042 153542 710278
rect 149266 708442 149502 708678
rect 149586 708442 149822 708678
rect 149266 708122 149502 708358
rect 149586 708122 149822 708358
rect 142986 684038 143222 684274
rect 143306 684038 143542 684274
rect 145546 706522 145782 706758
rect 145866 706522 146102 706758
rect 145546 706202 145782 706438
rect 145866 706202 146102 706438
rect 145546 686718 145782 686954
rect 145866 686718 146102 686954
rect 149266 690378 149502 690614
rect 149586 690378 149822 690614
rect 151826 705562 152062 705798
rect 152146 705562 152382 705798
rect 151826 705242 152062 705478
rect 152146 705242 152382 705478
rect 151826 693058 152062 693294
rect 152146 693058 152382 693294
rect 162986 711322 163222 711558
rect 163306 711322 163542 711558
rect 162986 711002 163222 711238
rect 163306 711002 163542 711238
rect 159266 709402 159502 709638
rect 159586 709402 159822 709638
rect 159266 709082 159502 709318
rect 159586 709082 159822 709318
rect 152986 694038 153222 694274
rect 153306 694038 153542 694274
rect 155546 707482 155782 707718
rect 155866 707482 156102 707718
rect 155546 707162 155782 707398
rect 155866 707162 156102 707398
rect 155546 696718 155782 696954
rect 155866 696718 156102 696954
rect 155546 676718 155782 676954
rect 155866 676718 156102 676954
rect 159266 700378 159502 700614
rect 159586 700378 159822 700614
rect 159266 680378 159502 680614
rect 159586 680378 159822 680614
rect 161826 704602 162062 704838
rect 162146 704602 162382 704838
rect 161826 704282 162062 704518
rect 162146 704282 162382 704518
rect 161826 683058 162062 683294
rect 162146 683058 162382 683294
rect 172986 710362 173222 710598
rect 173306 710362 173542 710598
rect 172986 710042 173222 710278
rect 173306 710042 173542 710278
rect 169266 708442 169502 708678
rect 169586 708442 169822 708678
rect 169266 708122 169502 708358
rect 169586 708122 169822 708358
rect 162986 684038 163222 684274
rect 163306 684038 163542 684274
rect 165546 706522 165782 706758
rect 165866 706522 166102 706758
rect 165546 706202 165782 706438
rect 165866 706202 166102 706438
rect 165546 686718 165782 686954
rect 165866 686718 166102 686954
rect 169266 690378 169502 690614
rect 169586 690378 169822 690614
rect 25546 666718 25782 666954
rect 25866 666718 26102 666954
rect 169266 670378 169502 670614
rect 169586 670378 169822 670614
rect 31008 663058 31244 663294
rect 165376 663058 165612 663294
rect 30328 653058 30564 653294
rect 166056 653058 166292 653294
rect 25546 646718 25782 646954
rect 25866 646718 26102 646954
rect 169266 650378 169502 650614
rect 169586 650378 169822 650614
rect 31008 643058 31244 643294
rect 165376 643058 165612 643294
rect 30328 633058 30564 633294
rect 166056 633058 166292 633294
rect 25546 626718 25782 626954
rect 25866 626718 26102 626954
rect 169266 630378 169502 630614
rect 169586 630378 169822 630614
rect 31008 623058 31244 623294
rect 165376 623058 165612 623294
rect 30328 613058 30564 613294
rect 166056 613058 166292 613294
rect 25546 606718 25782 606954
rect 25866 606718 26102 606954
rect 169266 610378 169502 610614
rect 169586 610378 169822 610614
rect 31008 603058 31244 603294
rect 165376 603058 165612 603294
rect 30328 593058 30564 593294
rect 166056 593058 166292 593294
rect 169266 590378 169502 590614
rect 169586 590378 169822 590614
rect 25546 586718 25782 586954
rect 25866 586718 26102 586954
rect 25546 566718 25782 566954
rect 25866 566718 26102 566954
rect 29266 570378 29502 570614
rect 29586 570378 29822 570614
rect 31826 573058 32062 573294
rect 32146 573058 32382 573294
rect 32986 574038 33222 574274
rect 33306 574038 33542 574274
rect 35546 576718 35782 576954
rect 35866 576718 36102 576954
rect 39266 580378 39502 580614
rect 39586 580378 39822 580614
rect 41826 583058 42062 583294
rect 42146 583058 42382 583294
rect 42986 584038 43222 584274
rect 43306 584038 43542 584274
rect 42986 564038 43222 564274
rect 43306 564038 43542 564274
rect 45546 586718 45782 586954
rect 45866 586718 46102 586954
rect 45546 566718 45782 566954
rect 45866 566718 46102 566954
rect 49266 570378 49502 570614
rect 49586 570378 49822 570614
rect 51826 573058 52062 573294
rect 52146 573058 52382 573294
rect 52986 574038 53222 574274
rect 53306 574038 53542 574274
rect 55546 576718 55782 576954
rect 55866 576718 56102 576954
rect 59266 580378 59502 580614
rect 59586 580378 59822 580614
rect 61826 583058 62062 583294
rect 62146 583058 62382 583294
rect 65546 586718 65782 586954
rect 65866 586718 66102 586954
rect 62986 584038 63222 584274
rect 63306 584038 63542 584274
rect 62986 564038 63222 564274
rect 63306 564038 63542 564274
rect 65546 566718 65782 566954
rect 65866 566718 66102 566954
rect 69266 570378 69502 570614
rect 69586 570378 69822 570614
rect 71826 573058 72062 573294
rect 72146 573058 72382 573294
rect 72986 574038 73222 574274
rect 73306 574038 73542 574274
rect 75546 576718 75782 576954
rect 75866 576718 76102 576954
rect 79266 580378 79502 580614
rect 79586 580378 79822 580614
rect 81826 583058 82062 583294
rect 82146 583058 82382 583294
rect 82986 584038 83222 584274
rect 83306 584038 83542 584274
rect 82986 564038 83222 564274
rect 83306 564038 83542 564274
rect 85546 586718 85782 586954
rect 85866 586718 86102 586954
rect 85546 566718 85782 566954
rect 85866 566718 86102 566954
rect 89266 570378 89502 570614
rect 89586 570378 89822 570614
rect 91826 573058 92062 573294
rect 92146 573058 92382 573294
rect 92986 574038 93222 574274
rect 93306 574038 93542 574274
rect 95546 576718 95782 576954
rect 95866 576718 96102 576954
rect 99266 580378 99502 580614
rect 99586 580378 99822 580614
rect 101826 583058 102062 583294
rect 102146 583058 102382 583294
rect 102986 584038 103222 584274
rect 103306 584038 103542 584274
rect 102986 564038 103222 564274
rect 103306 564038 103542 564274
rect 105546 586718 105782 586954
rect 105866 586718 106102 586954
rect 105546 566718 105782 566954
rect 105866 566718 106102 566954
rect 109266 570378 109502 570614
rect 109586 570378 109822 570614
rect 111826 573058 112062 573294
rect 112146 573058 112382 573294
rect 112986 574038 113222 574274
rect 113306 574038 113542 574274
rect 115546 576718 115782 576954
rect 115866 576718 116102 576954
rect 119266 580378 119502 580614
rect 119586 580378 119822 580614
rect 121826 583058 122062 583294
rect 122146 583058 122382 583294
rect 125546 586718 125782 586954
rect 125866 586718 126102 586954
rect 122986 584038 123222 584274
rect 123306 584038 123542 584274
rect 122986 564038 123222 564274
rect 123306 564038 123542 564274
rect 125546 566718 125782 566954
rect 125866 566718 126102 566954
rect 129266 570378 129502 570614
rect 129586 570378 129822 570614
rect 131826 573058 132062 573294
rect 132146 573058 132382 573294
rect 132986 574038 133222 574274
rect 133306 574038 133542 574274
rect 135546 576718 135782 576954
rect 135866 576718 136102 576954
rect 139266 580378 139502 580614
rect 139586 580378 139822 580614
rect 141826 583058 142062 583294
rect 142146 583058 142382 583294
rect 142986 584038 143222 584274
rect 143306 584038 143542 584274
rect 142986 564038 143222 564274
rect 143306 564038 143542 564274
rect 145546 586718 145782 586954
rect 145866 586718 146102 586954
rect 145546 566718 145782 566954
rect 145866 566718 146102 566954
rect 149266 570378 149502 570614
rect 149586 570378 149822 570614
rect 151826 573058 152062 573294
rect 152146 573058 152382 573294
rect 152986 574038 153222 574274
rect 153306 574038 153542 574274
rect 155546 576718 155782 576954
rect 155866 576718 156102 576954
rect 159266 580378 159502 580614
rect 159586 580378 159822 580614
rect 161826 583058 162062 583294
rect 162146 583058 162382 583294
rect 162986 584038 163222 584274
rect 163306 584038 163542 584274
rect 162986 564038 163222 564274
rect 163306 564038 163542 564274
rect 165546 586718 165782 586954
rect 165866 586718 166102 586954
rect 165546 566718 165782 566954
rect 165866 566718 166102 566954
rect 30328 553058 30564 553294
rect 166056 553058 166292 553294
rect 25546 546718 25782 546954
rect 25866 546718 26102 546954
rect 31008 543058 31244 543294
rect 165376 543058 165612 543294
rect 30328 533058 30564 533294
rect 166056 533058 166292 533294
rect 25546 526718 25782 526954
rect 25866 526718 26102 526954
rect 31008 523058 31244 523294
rect 165376 523058 165612 523294
rect 30328 513058 30564 513294
rect 166056 513058 166292 513294
rect 25546 506718 25782 506954
rect 25866 506718 26102 506954
rect 31008 503058 31244 503294
rect 165376 503058 165612 503294
rect 30328 493058 30564 493294
rect 166056 493058 166292 493294
rect 25546 486718 25782 486954
rect 25866 486718 26102 486954
rect 31008 483058 31244 483294
rect 165376 483058 165612 483294
rect 25546 466718 25782 466954
rect 25866 466718 26102 466954
rect 29266 470378 29502 470614
rect 29586 470378 29822 470614
rect 31826 473058 32062 473294
rect 32146 473058 32382 473294
rect 31826 453058 32062 453294
rect 32146 453058 32382 453294
rect 32986 474038 33222 474274
rect 33306 474038 33542 474274
rect 32986 454038 33222 454274
rect 33306 454038 33542 454274
rect 35546 456718 35782 456954
rect 35866 456718 36102 456954
rect 39266 460378 39502 460614
rect 39586 460378 39822 460614
rect 41826 463058 42062 463294
rect 42146 463058 42382 463294
rect 42986 464038 43222 464274
rect 43306 464038 43542 464274
rect 45546 466718 45782 466954
rect 45866 466718 46102 466954
rect 49266 470378 49502 470614
rect 49586 470378 49822 470614
rect 51826 473058 52062 473294
rect 52146 473058 52382 473294
rect 51826 453058 52062 453294
rect 52146 453058 52382 453294
rect 52986 474038 53222 474274
rect 53306 474038 53542 474274
rect 52986 454038 53222 454274
rect 53306 454038 53542 454274
rect 55546 456718 55782 456954
rect 55866 456718 56102 456954
rect 59266 460378 59502 460614
rect 59586 460378 59822 460614
rect 61826 463058 62062 463294
rect 62146 463058 62382 463294
rect 62986 464038 63222 464274
rect 63306 464038 63542 464274
rect 65546 466718 65782 466954
rect 65866 466718 66102 466954
rect 69266 470378 69502 470614
rect 69586 470378 69822 470614
rect 71826 473058 72062 473294
rect 72146 473058 72382 473294
rect 71826 453058 72062 453294
rect 72146 453058 72382 453294
rect 72986 474038 73222 474274
rect 73306 474038 73542 474274
rect 72986 454038 73222 454274
rect 73306 454038 73542 454274
rect 75546 456718 75782 456954
rect 75866 456718 76102 456954
rect 79266 460378 79502 460614
rect 79586 460378 79822 460614
rect 81826 463058 82062 463294
rect 82146 463058 82382 463294
rect 82986 464038 83222 464274
rect 83306 464038 83542 464274
rect 85546 466718 85782 466954
rect 85866 466718 86102 466954
rect 89266 470378 89502 470614
rect 89586 470378 89822 470614
rect 91826 473058 92062 473294
rect 92146 473058 92382 473294
rect 91826 453058 92062 453294
rect 92146 453058 92382 453294
rect 92986 474038 93222 474274
rect 93306 474038 93542 474274
rect 92986 454038 93222 454274
rect 93306 454038 93542 454274
rect 95546 456718 95782 456954
rect 95866 456718 96102 456954
rect 99266 460378 99502 460614
rect 99586 460378 99822 460614
rect 101826 463058 102062 463294
rect 102146 463058 102382 463294
rect 102986 464038 103222 464274
rect 103306 464038 103542 464274
rect 105546 466718 105782 466954
rect 105866 466718 106102 466954
rect 109266 470378 109502 470614
rect 109586 470378 109822 470614
rect 111826 473058 112062 473294
rect 112146 473058 112382 473294
rect 111826 453058 112062 453294
rect 112146 453058 112382 453294
rect 112986 474038 113222 474274
rect 113306 474038 113542 474274
rect 112986 454038 113222 454274
rect 113306 454038 113542 454274
rect 115546 456718 115782 456954
rect 115866 456718 116102 456954
rect 119266 460378 119502 460614
rect 119586 460378 119822 460614
rect 121826 463058 122062 463294
rect 122146 463058 122382 463294
rect 122986 464038 123222 464274
rect 123306 464038 123542 464274
rect 125546 466718 125782 466954
rect 125866 466718 126102 466954
rect 129266 470378 129502 470614
rect 129586 470378 129822 470614
rect 131826 473058 132062 473294
rect 132146 473058 132382 473294
rect 131826 453058 132062 453294
rect 132146 453058 132382 453294
rect 132986 474038 133222 474274
rect 133306 474038 133542 474274
rect 132986 454038 133222 454274
rect 133306 454038 133542 454274
rect 135546 456718 135782 456954
rect 135866 456718 136102 456954
rect 139266 460378 139502 460614
rect 139586 460378 139822 460614
rect 141826 463058 142062 463294
rect 142146 463058 142382 463294
rect 142986 464038 143222 464274
rect 143306 464038 143542 464274
rect 145546 466718 145782 466954
rect 145866 466718 146102 466954
rect 149266 470378 149502 470614
rect 149586 470378 149822 470614
rect 151826 473058 152062 473294
rect 152146 473058 152382 473294
rect 151826 453058 152062 453294
rect 152146 453058 152382 453294
rect 152986 474038 153222 474274
rect 153306 474038 153542 474274
rect 152986 454038 153222 454274
rect 153306 454038 153542 454274
rect 155546 456718 155782 456954
rect 155866 456718 156102 456954
rect 159266 460378 159502 460614
rect 159586 460378 159822 460614
rect 161826 463058 162062 463294
rect 162146 463058 162382 463294
rect 162986 464038 163222 464274
rect 163306 464038 163542 464274
rect 165546 466718 165782 466954
rect 165866 466718 166102 466954
rect 25546 446718 25782 446954
rect 25866 446718 26102 446954
rect 31008 443058 31244 443294
rect 165376 443058 165612 443294
rect 30328 433058 30564 433294
rect 166056 433058 166292 433294
rect 25546 426718 25782 426954
rect 25866 426718 26102 426954
rect 31008 423058 31244 423294
rect 165376 423058 165612 423294
rect 30328 413058 30564 413294
rect 166056 413058 166292 413294
rect 25546 406718 25782 406954
rect 25866 406718 26102 406954
rect 31008 403058 31244 403294
rect 165376 403058 165612 403294
rect 30328 393058 30564 393294
rect 166056 393058 166292 393294
rect 25546 386718 25782 386954
rect 25866 386718 26102 386954
rect 31008 383058 31244 383294
rect 165376 383058 165612 383294
rect 30328 373058 30564 373294
rect 166056 373058 166292 373294
rect 25546 366718 25782 366954
rect 25866 366718 26102 366954
rect 25546 346718 25782 346954
rect 25866 346718 26102 346954
rect 29266 350378 29502 350614
rect 29586 350378 29822 350614
rect 31826 353058 32062 353294
rect 32146 353058 32382 353294
rect 32986 354038 33222 354274
rect 33306 354038 33542 354274
rect 35546 356718 35782 356954
rect 35866 356718 36102 356954
rect 39266 360378 39502 360614
rect 39586 360378 39822 360614
rect 39266 340378 39502 340614
rect 39586 340378 39822 340614
rect 41826 363058 42062 363294
rect 42146 363058 42382 363294
rect 41826 343058 42062 343294
rect 42146 343058 42382 343294
rect 42986 344038 43222 344274
rect 43306 344038 43542 344274
rect 45546 346718 45782 346954
rect 45866 346718 46102 346954
rect 49266 350378 49502 350614
rect 49586 350378 49822 350614
rect 51826 353058 52062 353294
rect 52146 353058 52382 353294
rect 52986 354038 53222 354274
rect 53306 354038 53542 354274
rect 55546 356718 55782 356954
rect 55866 356718 56102 356954
rect 61826 363058 62062 363294
rect 62146 363058 62382 363294
rect 59266 360378 59502 360614
rect 59586 360378 59822 360614
rect 59266 340378 59502 340614
rect 59586 340378 59822 340614
rect 61826 343058 62062 343294
rect 62146 343058 62382 343294
rect 62986 344038 63222 344274
rect 63306 344038 63542 344274
rect 65546 346718 65782 346954
rect 65866 346718 66102 346954
rect 69266 350378 69502 350614
rect 69586 350378 69822 350614
rect 71826 353058 72062 353294
rect 72146 353058 72382 353294
rect 72986 354038 73222 354274
rect 73306 354038 73542 354274
rect 75546 356718 75782 356954
rect 75866 356718 76102 356954
rect 81826 363058 82062 363294
rect 82146 363058 82382 363294
rect 79266 360378 79502 360614
rect 79586 360378 79822 360614
rect 79266 340378 79502 340614
rect 79586 340378 79822 340614
rect 81826 343058 82062 343294
rect 82146 343058 82382 343294
rect 82986 344038 83222 344274
rect 83306 344038 83542 344274
rect 85546 346718 85782 346954
rect 85866 346718 86102 346954
rect 89266 350378 89502 350614
rect 89586 350378 89822 350614
rect 91826 353058 92062 353294
rect 92146 353058 92382 353294
rect 92986 354038 93222 354274
rect 93306 354038 93542 354274
rect 95546 356718 95782 356954
rect 95866 356718 96102 356954
rect 101826 363058 102062 363294
rect 102146 363058 102382 363294
rect 99266 360378 99502 360614
rect 99586 360378 99822 360614
rect 99266 340378 99502 340614
rect 99586 340378 99822 340614
rect 101826 343058 102062 343294
rect 102146 343058 102382 343294
rect 102986 344038 103222 344274
rect 103306 344038 103542 344274
rect 105546 346718 105782 346954
rect 105866 346718 106102 346954
rect 109266 350378 109502 350614
rect 109586 350378 109822 350614
rect 111826 353058 112062 353294
rect 112146 353058 112382 353294
rect 112986 354038 113222 354274
rect 113306 354038 113542 354274
rect 115546 356718 115782 356954
rect 115866 356718 116102 356954
rect 121826 363058 122062 363294
rect 122146 363058 122382 363294
rect 119266 360378 119502 360614
rect 119586 360378 119822 360614
rect 119266 340378 119502 340614
rect 119586 340378 119822 340614
rect 121826 343058 122062 343294
rect 122146 343058 122382 343294
rect 122986 344038 123222 344274
rect 123306 344038 123542 344274
rect 125546 346718 125782 346954
rect 125866 346718 126102 346954
rect 129266 350378 129502 350614
rect 129586 350378 129822 350614
rect 131826 353058 132062 353294
rect 132146 353058 132382 353294
rect 132986 354038 133222 354274
rect 133306 354038 133542 354274
rect 135546 356718 135782 356954
rect 135866 356718 136102 356954
rect 141826 363058 142062 363294
rect 142146 363058 142382 363294
rect 139266 360378 139502 360614
rect 139586 360378 139822 360614
rect 139266 340378 139502 340614
rect 139586 340378 139822 340614
rect 141826 343058 142062 343294
rect 142146 343058 142382 343294
rect 142986 344038 143222 344274
rect 143306 344038 143542 344274
rect 145546 346718 145782 346954
rect 145866 346718 146102 346954
rect 149266 350378 149502 350614
rect 149586 350378 149822 350614
rect 151826 353058 152062 353294
rect 152146 353058 152382 353294
rect 152986 354038 153222 354274
rect 153306 354038 153542 354274
rect 155546 356718 155782 356954
rect 155866 356718 156102 356954
rect 159266 360378 159502 360614
rect 159586 360378 159822 360614
rect 159266 340378 159502 340614
rect 159586 340378 159822 340614
rect 161826 363058 162062 363294
rect 162146 363058 162382 363294
rect 161826 343058 162062 343294
rect 162146 343058 162382 343294
rect 162986 344038 163222 344274
rect 163306 344038 163542 344274
rect 165546 346718 165782 346954
rect 165866 346718 166102 346954
rect 30328 333058 30564 333294
rect 166056 333058 166292 333294
rect 25546 326718 25782 326954
rect 25866 326718 26102 326954
rect 31008 323058 31244 323294
rect 165376 323058 165612 323294
rect 30328 313058 30564 313294
rect 166056 313058 166292 313294
rect 25546 306718 25782 306954
rect 25866 306718 26102 306954
rect 31008 303058 31244 303294
rect 165376 303058 165612 303294
rect 30328 293058 30564 293294
rect 166056 293058 166292 293294
rect 25546 286718 25782 286954
rect 25866 286718 26102 286954
rect 31008 283058 31244 283294
rect 165376 283058 165612 283294
rect 30328 273058 30564 273294
rect 166056 273058 166292 273294
rect 25546 266718 25782 266954
rect 25866 266718 26102 266954
rect 31008 263058 31244 263294
rect 165376 263058 165612 263294
rect 25546 246718 25782 246954
rect 25866 246718 26102 246954
rect 29266 250378 29502 250614
rect 29586 250378 29822 250614
rect 29266 230378 29502 230614
rect 29586 230378 29822 230614
rect 31826 233058 32062 233294
rect 32146 233058 32382 233294
rect 32986 234038 33222 234274
rect 33306 234038 33542 234274
rect 35546 236718 35782 236954
rect 35866 236718 36102 236954
rect 25546 226718 25782 226954
rect 25866 226718 26102 226954
rect 39266 240378 39502 240614
rect 39586 240378 39822 240614
rect 41826 243058 42062 243294
rect 42146 243058 42382 243294
rect 42986 244038 43222 244274
rect 43306 244038 43542 244274
rect 45546 246718 45782 246954
rect 45866 246718 46102 246954
rect 49266 250378 49502 250614
rect 49586 250378 49822 250614
rect 49266 230378 49502 230614
rect 49586 230378 49822 230614
rect 51826 233058 52062 233294
rect 52146 233058 52382 233294
rect 52986 234038 53222 234274
rect 53306 234038 53542 234274
rect 55546 236718 55782 236954
rect 55866 236718 56102 236954
rect 59266 240378 59502 240614
rect 59586 240378 59822 240614
rect 61826 243058 62062 243294
rect 62146 243058 62382 243294
rect 62986 244038 63222 244274
rect 63306 244038 63542 244274
rect 65546 246718 65782 246954
rect 65866 246718 66102 246954
rect 69266 250378 69502 250614
rect 69586 250378 69822 250614
rect 69266 230378 69502 230614
rect 69586 230378 69822 230614
rect 71826 233058 72062 233294
rect 72146 233058 72382 233294
rect 72986 234038 73222 234274
rect 73306 234038 73542 234274
rect 75546 236718 75782 236954
rect 75866 236718 76102 236954
rect 79266 240378 79502 240614
rect 79586 240378 79822 240614
rect 81826 243058 82062 243294
rect 82146 243058 82382 243294
rect 82986 244038 83222 244274
rect 83306 244038 83542 244274
rect 85546 246718 85782 246954
rect 85866 246718 86102 246954
rect 89266 250378 89502 250614
rect 89586 250378 89822 250614
rect 89266 230378 89502 230614
rect 89586 230378 89822 230614
rect 91826 233058 92062 233294
rect 92146 233058 92382 233294
rect 92986 234038 93222 234274
rect 93306 234038 93542 234274
rect 95546 236718 95782 236954
rect 95866 236718 96102 236954
rect 99266 240378 99502 240614
rect 99586 240378 99822 240614
rect 101826 243058 102062 243294
rect 102146 243058 102382 243294
rect 102986 244038 103222 244274
rect 103306 244038 103542 244274
rect 105546 246718 105782 246954
rect 105866 246718 106102 246954
rect 109266 250378 109502 250614
rect 109586 250378 109822 250614
rect 109266 230378 109502 230614
rect 109586 230378 109822 230614
rect 111826 233058 112062 233294
rect 112146 233058 112382 233294
rect 112986 234038 113222 234274
rect 113306 234038 113542 234274
rect 115546 236718 115782 236954
rect 115866 236718 116102 236954
rect 119266 240378 119502 240614
rect 119586 240378 119822 240614
rect 121826 243058 122062 243294
rect 122146 243058 122382 243294
rect 122986 244038 123222 244274
rect 123306 244038 123542 244274
rect 125546 246718 125782 246954
rect 125866 246718 126102 246954
rect 129266 250378 129502 250614
rect 129586 250378 129822 250614
rect 129266 230378 129502 230614
rect 129586 230378 129822 230614
rect 131826 233058 132062 233294
rect 132146 233058 132382 233294
rect 132986 234038 133222 234274
rect 133306 234038 133542 234274
rect 135546 236718 135782 236954
rect 135866 236718 136102 236954
rect 139266 240378 139502 240614
rect 139586 240378 139822 240614
rect 141826 243058 142062 243294
rect 142146 243058 142382 243294
rect 142986 244038 143222 244274
rect 143306 244038 143542 244274
rect 145546 246718 145782 246954
rect 145866 246718 146102 246954
rect 149266 250378 149502 250614
rect 149586 250378 149822 250614
rect 149266 230378 149502 230614
rect 149586 230378 149822 230614
rect 151826 233058 152062 233294
rect 152146 233058 152382 233294
rect 152986 234038 153222 234274
rect 153306 234038 153542 234274
rect 155546 236718 155782 236954
rect 155866 236718 156102 236954
rect 159266 240378 159502 240614
rect 159586 240378 159822 240614
rect 161826 243058 162062 243294
rect 162146 243058 162382 243294
rect 162986 244038 163222 244274
rect 163306 244038 163542 244274
rect 165546 246718 165782 246954
rect 165866 246718 166102 246954
rect 171826 705562 172062 705798
rect 172146 705562 172382 705798
rect 171826 705242 172062 705478
rect 172146 705242 172382 705478
rect 171826 693058 172062 693294
rect 172146 693058 172382 693294
rect 171826 673058 172062 673294
rect 172146 673058 172382 673294
rect 171826 653058 172062 653294
rect 172146 653058 172382 653294
rect 171826 633058 172062 633294
rect 172146 633058 172382 633294
rect 171826 613058 172062 613294
rect 172146 613058 172382 613294
rect 171826 593058 172062 593294
rect 172146 593058 172382 593294
rect 169266 570378 169502 570614
rect 169586 570378 169822 570614
rect 169266 550378 169502 550614
rect 169586 550378 169822 550614
rect 169266 530378 169502 530614
rect 169586 530378 169822 530614
rect 169266 510378 169502 510614
rect 169586 510378 169822 510614
rect 169266 490378 169502 490614
rect 169586 490378 169822 490614
rect 169266 470378 169502 470614
rect 169586 470378 169822 470614
rect 169266 450378 169502 450614
rect 169586 450378 169822 450614
rect 169266 430378 169502 430614
rect 169586 430378 169822 430614
rect 182986 711322 183222 711558
rect 183306 711322 183542 711558
rect 182986 711002 183222 711238
rect 183306 711002 183542 711238
rect 179266 709402 179502 709638
rect 179586 709402 179822 709638
rect 179266 709082 179502 709318
rect 179586 709082 179822 709318
rect 175546 707482 175782 707718
rect 175866 707482 176102 707718
rect 175546 707162 175782 707398
rect 175866 707162 176102 707398
rect 172986 694038 173222 694274
rect 173306 694038 173542 694274
rect 172986 674038 173222 674274
rect 173306 674038 173542 674274
rect 172986 654038 173222 654274
rect 173306 654038 173542 654274
rect 172986 634038 173222 634274
rect 173306 634038 173542 634274
rect 172986 614038 173222 614274
rect 173306 614038 173542 614274
rect 172986 594038 173222 594274
rect 173306 594038 173542 594274
rect 171826 573058 172062 573294
rect 172146 573058 172382 573294
rect 171826 553058 172062 553294
rect 172146 553058 172382 553294
rect 171826 533058 172062 533294
rect 172146 533058 172382 533294
rect 171826 513058 172062 513294
rect 172146 513058 172382 513294
rect 171826 493058 172062 493294
rect 172146 493058 172382 493294
rect 171826 473058 172062 473294
rect 172146 473058 172382 473294
rect 171826 453058 172062 453294
rect 172146 453058 172382 453294
rect 169266 410378 169502 410614
rect 169586 410378 169822 410614
rect 169266 390378 169502 390614
rect 169586 390378 169822 390614
rect 169266 370378 169502 370614
rect 169586 370378 169822 370614
rect 169266 350378 169502 350614
rect 169586 350378 169822 350614
rect 169266 330378 169502 330614
rect 169586 330378 169822 330614
rect 169266 310378 169502 310614
rect 169586 310378 169822 310614
rect 169266 290378 169502 290614
rect 169586 290378 169822 290614
rect 169266 270378 169502 270614
rect 169586 270378 169822 270614
rect 169266 250378 169502 250614
rect 169586 250378 169822 250614
rect 169266 230378 169502 230614
rect 169586 230378 169822 230614
rect 31008 223058 31244 223294
rect 165376 223058 165612 223294
rect 30328 213058 30564 213294
rect 166056 213058 166292 213294
rect 25546 206718 25782 206954
rect 25866 206718 26102 206954
rect 171826 433058 172062 433294
rect 172146 433058 172382 433294
rect 171826 413058 172062 413294
rect 172146 413058 172382 413294
rect 171826 393058 172062 393294
rect 172146 393058 172382 393294
rect 171826 373058 172062 373294
rect 172146 373058 172382 373294
rect 171826 353058 172062 353294
rect 172146 353058 172382 353294
rect 172986 574038 173222 574274
rect 173306 574038 173542 574274
rect 172986 554038 173222 554274
rect 173306 554038 173542 554274
rect 172986 534038 173222 534274
rect 173306 534038 173542 534274
rect 172986 514038 173222 514274
rect 173306 514038 173542 514274
rect 172986 494038 173222 494274
rect 173306 494038 173542 494274
rect 172986 474038 173222 474274
rect 173306 474038 173542 474274
rect 172986 454038 173222 454274
rect 173306 454038 173542 454274
rect 175546 696718 175782 696954
rect 175866 696718 176102 696954
rect 175546 676718 175782 676954
rect 175866 676718 176102 676954
rect 175546 656718 175782 656954
rect 175866 656718 176102 656954
rect 175546 636718 175782 636954
rect 175866 636718 176102 636954
rect 175546 616718 175782 616954
rect 175866 616718 176102 616954
rect 175546 596718 175782 596954
rect 175866 596718 176102 596954
rect 175546 576718 175782 576954
rect 175866 576718 176102 576954
rect 175546 556718 175782 556954
rect 175866 556718 176102 556954
rect 175546 536718 175782 536954
rect 175866 536718 176102 536954
rect 175546 516718 175782 516954
rect 175866 516718 176102 516954
rect 175546 496718 175782 496954
rect 175866 496718 176102 496954
rect 175546 476718 175782 476954
rect 175866 476718 176102 476954
rect 175546 456718 175782 456954
rect 175866 456718 176102 456954
rect 172986 434038 173222 434274
rect 173306 434038 173542 434274
rect 175546 436718 175782 436954
rect 175866 436718 176102 436954
rect 172986 414038 173222 414274
rect 173306 414038 173542 414274
rect 172986 394038 173222 394274
rect 173306 394038 173542 394274
rect 172986 374038 173222 374274
rect 173306 374038 173542 374274
rect 172986 354038 173222 354274
rect 173306 354038 173542 354274
rect 171826 333058 172062 333294
rect 172146 333058 172382 333294
rect 171826 313058 172062 313294
rect 172146 313058 172382 313294
rect 171826 293058 172062 293294
rect 172146 293058 172382 293294
rect 171826 273058 172062 273294
rect 172146 273058 172382 273294
rect 171826 253058 172062 253294
rect 172146 253058 172382 253294
rect 171826 233058 172062 233294
rect 172146 233058 172382 233294
rect 169266 210378 169502 210614
rect 169586 210378 169822 210614
rect 31008 203058 31244 203294
rect 165376 203058 165612 203294
rect 30328 193058 30564 193294
rect 166056 193058 166292 193294
rect 25546 186718 25782 186954
rect 25866 186718 26102 186954
rect 169266 190378 169502 190614
rect 169586 190378 169822 190614
rect 31008 183058 31244 183294
rect 165376 183058 165612 183294
rect 30328 173058 30564 173294
rect 166056 173058 166292 173294
rect 25546 166718 25782 166954
rect 25866 166718 26102 166954
rect 169266 170378 169502 170614
rect 169586 170378 169822 170614
rect 31008 163058 31244 163294
rect 165376 163058 165612 163294
rect 30328 153058 30564 153294
rect 166056 153058 166292 153294
rect 25546 146718 25782 146954
rect 25866 146718 26102 146954
rect 169266 150378 169502 150614
rect 169586 150378 169822 150614
rect 25546 126718 25782 126954
rect 25866 126718 26102 126954
rect 29266 130378 29502 130614
rect 29586 130378 29822 130614
rect 31826 133058 32062 133294
rect 32146 133058 32382 133294
rect 32986 134038 33222 134274
rect 33306 134038 33542 134274
rect 35546 136718 35782 136954
rect 35866 136718 36102 136954
rect 35546 116718 35782 116954
rect 35866 116718 36102 116954
rect 39266 120378 39502 120614
rect 39586 120378 39822 120614
rect 41826 123058 42062 123294
rect 42146 123058 42382 123294
rect 42986 124038 43222 124274
rect 43306 124038 43542 124274
rect 45546 126718 45782 126954
rect 45866 126718 46102 126954
rect 49266 130378 49502 130614
rect 49586 130378 49822 130614
rect 51826 133058 52062 133294
rect 52146 133058 52382 133294
rect 52986 134038 53222 134274
rect 53306 134038 53542 134274
rect 55546 136718 55782 136954
rect 55866 136718 56102 136954
rect 55546 116718 55782 116954
rect 55866 116718 56102 116954
rect 59266 120378 59502 120614
rect 59586 120378 59822 120614
rect 61826 123058 62062 123294
rect 62146 123058 62382 123294
rect 62986 124038 63222 124274
rect 63306 124038 63542 124274
rect 65546 126718 65782 126954
rect 65866 126718 66102 126954
rect 69266 130378 69502 130614
rect 69586 130378 69822 130614
rect 71826 133058 72062 133294
rect 72146 133058 72382 133294
rect 72986 134038 73222 134274
rect 73306 134038 73542 134274
rect 75546 136718 75782 136954
rect 75866 136718 76102 136954
rect 75546 116718 75782 116954
rect 75866 116718 76102 116954
rect 79266 120378 79502 120614
rect 79586 120378 79822 120614
rect 81826 123058 82062 123294
rect 82146 123058 82382 123294
rect 82986 124038 83222 124274
rect 83306 124038 83542 124274
rect 85546 126718 85782 126954
rect 85866 126718 86102 126954
rect 89266 130378 89502 130614
rect 89586 130378 89822 130614
rect 91826 133058 92062 133294
rect 92146 133058 92382 133294
rect 92986 134038 93222 134274
rect 93306 134038 93542 134274
rect 95546 136718 95782 136954
rect 95866 136718 96102 136954
rect 95546 116718 95782 116954
rect 95866 116718 96102 116954
rect 99266 120378 99502 120614
rect 99586 120378 99822 120614
rect 101826 123058 102062 123294
rect 102146 123058 102382 123294
rect 102986 124038 103222 124274
rect 103306 124038 103542 124274
rect 105546 126718 105782 126954
rect 105866 126718 106102 126954
rect 109266 130378 109502 130614
rect 109586 130378 109822 130614
rect 111826 133058 112062 133294
rect 112146 133058 112382 133294
rect 112986 134038 113222 134274
rect 113306 134038 113542 134274
rect 115546 136718 115782 136954
rect 115866 136718 116102 136954
rect 115546 116718 115782 116954
rect 115866 116718 116102 116954
rect 119266 120378 119502 120614
rect 119586 120378 119822 120614
rect 121826 123058 122062 123294
rect 122146 123058 122382 123294
rect 122986 124038 123222 124274
rect 123306 124038 123542 124274
rect 125546 126718 125782 126954
rect 125866 126718 126102 126954
rect 129266 130378 129502 130614
rect 129586 130378 129822 130614
rect 131826 133058 132062 133294
rect 132146 133058 132382 133294
rect 132986 134038 133222 134274
rect 133306 134038 133542 134274
rect 135546 136718 135782 136954
rect 135866 136718 136102 136954
rect 135546 116718 135782 116954
rect 135866 116718 136102 116954
rect 139266 120378 139502 120614
rect 139586 120378 139822 120614
rect 141826 123058 142062 123294
rect 142146 123058 142382 123294
rect 142986 124038 143222 124274
rect 143306 124038 143542 124274
rect 145546 126718 145782 126954
rect 145866 126718 146102 126954
rect 149266 130378 149502 130614
rect 149586 130378 149822 130614
rect 151826 133058 152062 133294
rect 152146 133058 152382 133294
rect 152986 134038 153222 134274
rect 153306 134038 153542 134274
rect 155546 136718 155782 136954
rect 155866 136718 156102 136954
rect 155546 116718 155782 116954
rect 155866 116718 156102 116954
rect 159266 120378 159502 120614
rect 159586 120378 159822 120614
rect 161826 123058 162062 123294
rect 162146 123058 162382 123294
rect 162986 124038 163222 124274
rect 163306 124038 163542 124274
rect 165546 126718 165782 126954
rect 165866 126718 166102 126954
rect 169266 130378 169502 130614
rect 169586 130378 169822 130614
rect 25546 106718 25782 106954
rect 25866 106718 26102 106954
rect 169266 110378 169502 110614
rect 169586 110378 169822 110614
rect 31008 103058 31244 103294
rect 165376 103058 165612 103294
rect 30328 93058 30564 93294
rect 166056 93058 166292 93294
rect 25546 86718 25782 86954
rect 25866 86718 26102 86954
rect 169266 90378 169502 90614
rect 169586 90378 169822 90614
rect 31008 83058 31244 83294
rect 165376 83058 165612 83294
rect 30328 73058 30564 73294
rect 166056 73058 166292 73294
rect 25546 66718 25782 66954
rect 25866 66718 26102 66954
rect 169266 70378 169502 70614
rect 169586 70378 169822 70614
rect 31008 63058 31244 63294
rect 165376 63058 165612 63294
rect 30328 53058 30564 53294
rect 166056 53058 166292 53294
rect 25546 46718 25782 46954
rect 25866 46718 26102 46954
rect 169266 50378 169502 50614
rect 169586 50378 169822 50614
rect 31008 43058 31244 43294
rect 165376 43058 165612 43294
rect 30328 33058 30564 33294
rect 166056 33058 166292 33294
rect 169266 30378 169502 30614
rect 169586 30378 169822 30614
rect 25546 26718 25782 26954
rect 25866 26718 26102 26954
rect 25546 6718 25782 6954
rect 25866 6718 26102 6954
rect 25546 -2502 25782 -2266
rect 25866 -2502 26102 -2266
rect 25546 -2822 25782 -2586
rect 25866 -2822 26102 -2586
rect 29266 10378 29502 10614
rect 29586 10378 29822 10614
rect 31826 13058 32062 13294
rect 32146 13058 32382 13294
rect 31826 -1542 32062 -1306
rect 32146 -1542 32382 -1306
rect 31826 -1862 32062 -1626
rect 32146 -1862 32382 -1626
rect 32986 14038 33222 14274
rect 33306 14038 33542 14274
rect 29266 -4422 29502 -4186
rect 29586 -4422 29822 -4186
rect 29266 -4742 29502 -4506
rect 29586 -4742 29822 -4506
rect 22986 -7302 23222 -7066
rect 23306 -7302 23542 -7066
rect 22986 -7622 23222 -7386
rect 23306 -7622 23542 -7386
rect 35546 16718 35782 16954
rect 35866 16718 36102 16954
rect 35546 -3462 35782 -3226
rect 35866 -3462 36102 -3226
rect 35546 -3782 35782 -3546
rect 35866 -3782 36102 -3546
rect 39266 20378 39502 20614
rect 39586 20378 39822 20614
rect 41826 23058 42062 23294
rect 42146 23058 42382 23294
rect 41826 3058 42062 3294
rect 42146 3058 42382 3294
rect 41826 -582 42062 -346
rect 42146 -582 42382 -346
rect 41826 -902 42062 -666
rect 42146 -902 42382 -666
rect 42986 24038 43222 24274
rect 43306 24038 43542 24274
rect 39266 -5382 39502 -5146
rect 39586 -5382 39822 -5146
rect 39266 -5702 39502 -5466
rect 39586 -5702 39822 -5466
rect 32986 -6342 33222 -6106
rect 33306 -6342 33542 -6106
rect 32986 -6662 33222 -6426
rect 33306 -6662 33542 -6426
rect 45546 26718 45782 26954
rect 45866 26718 46102 26954
rect 45546 6718 45782 6954
rect 45866 6718 46102 6954
rect 45546 -2502 45782 -2266
rect 45866 -2502 46102 -2266
rect 45546 -2822 45782 -2586
rect 45866 -2822 46102 -2586
rect 49266 10378 49502 10614
rect 49586 10378 49822 10614
rect 51826 13058 52062 13294
rect 52146 13058 52382 13294
rect 51826 -1542 52062 -1306
rect 52146 -1542 52382 -1306
rect 51826 -1862 52062 -1626
rect 52146 -1862 52382 -1626
rect 52986 14038 53222 14274
rect 53306 14038 53542 14274
rect 49266 -4422 49502 -4186
rect 49586 -4422 49822 -4186
rect 49266 -4742 49502 -4506
rect 49586 -4742 49822 -4506
rect 42986 -7302 43222 -7066
rect 43306 -7302 43542 -7066
rect 42986 -7622 43222 -7386
rect 43306 -7622 43542 -7386
rect 55546 16718 55782 16954
rect 55866 16718 56102 16954
rect 55546 -3462 55782 -3226
rect 55866 -3462 56102 -3226
rect 55546 -3782 55782 -3546
rect 55866 -3782 56102 -3546
rect 59266 20378 59502 20614
rect 59586 20378 59822 20614
rect 61826 23058 62062 23294
rect 62146 23058 62382 23294
rect 61826 3058 62062 3294
rect 62146 3058 62382 3294
rect 61826 -582 62062 -346
rect 62146 -582 62382 -346
rect 61826 -902 62062 -666
rect 62146 -902 62382 -666
rect 62986 24038 63222 24274
rect 63306 24038 63542 24274
rect 59266 -5382 59502 -5146
rect 59586 -5382 59822 -5146
rect 59266 -5702 59502 -5466
rect 59586 -5702 59822 -5466
rect 52986 -6342 53222 -6106
rect 53306 -6342 53542 -6106
rect 52986 -6662 53222 -6426
rect 53306 -6662 53542 -6426
rect 65546 26718 65782 26954
rect 65866 26718 66102 26954
rect 65546 6718 65782 6954
rect 65866 6718 66102 6954
rect 65546 -2502 65782 -2266
rect 65866 -2502 66102 -2266
rect 65546 -2822 65782 -2586
rect 65866 -2822 66102 -2586
rect 69266 10378 69502 10614
rect 69586 10378 69822 10614
rect 71826 13058 72062 13294
rect 72146 13058 72382 13294
rect 71826 -1542 72062 -1306
rect 72146 -1542 72382 -1306
rect 71826 -1862 72062 -1626
rect 72146 -1862 72382 -1626
rect 72986 14038 73222 14274
rect 73306 14038 73542 14274
rect 69266 -4422 69502 -4186
rect 69586 -4422 69822 -4186
rect 69266 -4742 69502 -4506
rect 69586 -4742 69822 -4506
rect 62986 -7302 63222 -7066
rect 63306 -7302 63542 -7066
rect 62986 -7622 63222 -7386
rect 63306 -7622 63542 -7386
rect 75546 16718 75782 16954
rect 75866 16718 76102 16954
rect 75546 -3462 75782 -3226
rect 75866 -3462 76102 -3226
rect 75546 -3782 75782 -3546
rect 75866 -3782 76102 -3546
rect 79266 20378 79502 20614
rect 79586 20378 79822 20614
rect 81826 23058 82062 23294
rect 82146 23058 82382 23294
rect 81826 3058 82062 3294
rect 82146 3058 82382 3294
rect 81826 -582 82062 -346
rect 82146 -582 82382 -346
rect 81826 -902 82062 -666
rect 82146 -902 82382 -666
rect 82986 24038 83222 24274
rect 83306 24038 83542 24274
rect 79266 -5382 79502 -5146
rect 79586 -5382 79822 -5146
rect 79266 -5702 79502 -5466
rect 79586 -5702 79822 -5466
rect 72986 -6342 73222 -6106
rect 73306 -6342 73542 -6106
rect 72986 -6662 73222 -6426
rect 73306 -6662 73542 -6426
rect 85546 26718 85782 26954
rect 85866 26718 86102 26954
rect 85546 6718 85782 6954
rect 85866 6718 86102 6954
rect 85546 -2502 85782 -2266
rect 85866 -2502 86102 -2266
rect 85546 -2822 85782 -2586
rect 85866 -2822 86102 -2586
rect 89266 10378 89502 10614
rect 89586 10378 89822 10614
rect 91826 13058 92062 13294
rect 92146 13058 92382 13294
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 92986 14038 93222 14274
rect 93306 14038 93542 14274
rect 89266 -4422 89502 -4186
rect 89586 -4422 89822 -4186
rect 89266 -4742 89502 -4506
rect 89586 -4742 89822 -4506
rect 82986 -7302 83222 -7066
rect 83306 -7302 83542 -7066
rect 82986 -7622 83222 -7386
rect 83306 -7622 83542 -7386
rect 95546 16718 95782 16954
rect 95866 16718 96102 16954
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 20378 99502 20614
rect 99586 20378 99822 20614
rect 101826 23058 102062 23294
rect 102146 23058 102382 23294
rect 101826 3058 102062 3294
rect 102146 3058 102382 3294
rect 101826 -582 102062 -346
rect 102146 -582 102382 -346
rect 101826 -902 102062 -666
rect 102146 -902 102382 -666
rect 102986 24038 103222 24274
rect 103306 24038 103542 24274
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 92986 -6342 93222 -6106
rect 93306 -6342 93542 -6106
rect 92986 -6662 93222 -6426
rect 93306 -6662 93542 -6426
rect 105546 26718 105782 26954
rect 105866 26718 106102 26954
rect 105546 6718 105782 6954
rect 105866 6718 106102 6954
rect 105546 -2502 105782 -2266
rect 105866 -2502 106102 -2266
rect 105546 -2822 105782 -2586
rect 105866 -2822 106102 -2586
rect 109266 10378 109502 10614
rect 109586 10378 109822 10614
rect 111826 13058 112062 13294
rect 112146 13058 112382 13294
rect 111826 -1542 112062 -1306
rect 112146 -1542 112382 -1306
rect 111826 -1862 112062 -1626
rect 112146 -1862 112382 -1626
rect 112986 14038 113222 14274
rect 113306 14038 113542 14274
rect 109266 -4422 109502 -4186
rect 109586 -4422 109822 -4186
rect 109266 -4742 109502 -4506
rect 109586 -4742 109822 -4506
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 115546 16718 115782 16954
rect 115866 16718 116102 16954
rect 115546 -3462 115782 -3226
rect 115866 -3462 116102 -3226
rect 115546 -3782 115782 -3546
rect 115866 -3782 116102 -3546
rect 119266 20378 119502 20614
rect 119586 20378 119822 20614
rect 121826 23058 122062 23294
rect 122146 23058 122382 23294
rect 121826 3058 122062 3294
rect 122146 3058 122382 3294
rect 121826 -582 122062 -346
rect 122146 -582 122382 -346
rect 121826 -902 122062 -666
rect 122146 -902 122382 -666
rect 122986 24038 123222 24274
rect 123306 24038 123542 24274
rect 119266 -5382 119502 -5146
rect 119586 -5382 119822 -5146
rect 119266 -5702 119502 -5466
rect 119586 -5702 119822 -5466
rect 112986 -6342 113222 -6106
rect 113306 -6342 113542 -6106
rect 112986 -6662 113222 -6426
rect 113306 -6662 113542 -6426
rect 125546 26718 125782 26954
rect 125866 26718 126102 26954
rect 125546 6718 125782 6954
rect 125866 6718 126102 6954
rect 125546 -2502 125782 -2266
rect 125866 -2502 126102 -2266
rect 125546 -2822 125782 -2586
rect 125866 -2822 126102 -2586
rect 129266 10378 129502 10614
rect 129586 10378 129822 10614
rect 131826 13058 132062 13294
rect 132146 13058 132382 13294
rect 131826 -1542 132062 -1306
rect 132146 -1542 132382 -1306
rect 131826 -1862 132062 -1626
rect 132146 -1862 132382 -1626
rect 132986 14038 133222 14274
rect 133306 14038 133542 14274
rect 129266 -4422 129502 -4186
rect 129586 -4422 129822 -4186
rect 129266 -4742 129502 -4506
rect 129586 -4742 129822 -4506
rect 122986 -7302 123222 -7066
rect 123306 -7302 123542 -7066
rect 122986 -7622 123222 -7386
rect 123306 -7622 123542 -7386
rect 135546 16718 135782 16954
rect 135866 16718 136102 16954
rect 135546 -3462 135782 -3226
rect 135866 -3462 136102 -3226
rect 135546 -3782 135782 -3546
rect 135866 -3782 136102 -3546
rect 139266 20378 139502 20614
rect 139586 20378 139822 20614
rect 141826 23058 142062 23294
rect 142146 23058 142382 23294
rect 141826 3058 142062 3294
rect 142146 3058 142382 3294
rect 141826 -582 142062 -346
rect 142146 -582 142382 -346
rect 141826 -902 142062 -666
rect 142146 -902 142382 -666
rect 142986 24038 143222 24274
rect 143306 24038 143542 24274
rect 139266 -5382 139502 -5146
rect 139586 -5382 139822 -5146
rect 139266 -5702 139502 -5466
rect 139586 -5702 139822 -5466
rect 132986 -6342 133222 -6106
rect 133306 -6342 133542 -6106
rect 132986 -6662 133222 -6426
rect 133306 -6662 133542 -6426
rect 145546 26718 145782 26954
rect 145866 26718 146102 26954
rect 145546 6718 145782 6954
rect 145866 6718 146102 6954
rect 145546 -2502 145782 -2266
rect 145866 -2502 146102 -2266
rect 145546 -2822 145782 -2586
rect 145866 -2822 146102 -2586
rect 149266 10378 149502 10614
rect 149586 10378 149822 10614
rect 151826 13058 152062 13294
rect 152146 13058 152382 13294
rect 151826 -1542 152062 -1306
rect 152146 -1542 152382 -1306
rect 151826 -1862 152062 -1626
rect 152146 -1862 152382 -1626
rect 152986 14038 153222 14274
rect 153306 14038 153542 14274
rect 149266 -4422 149502 -4186
rect 149586 -4422 149822 -4186
rect 149266 -4742 149502 -4506
rect 149586 -4742 149822 -4506
rect 142986 -7302 143222 -7066
rect 143306 -7302 143542 -7066
rect 142986 -7622 143222 -7386
rect 143306 -7622 143542 -7386
rect 155546 16718 155782 16954
rect 155866 16718 156102 16954
rect 155546 -3462 155782 -3226
rect 155866 -3462 156102 -3226
rect 155546 -3782 155782 -3546
rect 155866 -3782 156102 -3546
rect 159266 20378 159502 20614
rect 159586 20378 159822 20614
rect 161826 23058 162062 23294
rect 162146 23058 162382 23294
rect 161826 3058 162062 3294
rect 162146 3058 162382 3294
rect 161826 -582 162062 -346
rect 162146 -582 162382 -346
rect 161826 -902 162062 -666
rect 162146 -902 162382 -666
rect 162986 24038 163222 24274
rect 163306 24038 163542 24274
rect 159266 -5382 159502 -5146
rect 159586 -5382 159822 -5146
rect 159266 -5702 159502 -5466
rect 159586 -5702 159822 -5466
rect 152986 -6342 153222 -6106
rect 153306 -6342 153542 -6106
rect 152986 -6662 153222 -6426
rect 153306 -6662 153542 -6426
rect 165546 26718 165782 26954
rect 165866 26718 166102 26954
rect 165546 6718 165782 6954
rect 165866 6718 166102 6954
rect 165546 -2502 165782 -2266
rect 165866 -2502 166102 -2266
rect 165546 -2822 165782 -2586
rect 165866 -2822 166102 -2586
rect 169266 10378 169502 10614
rect 169586 10378 169822 10614
rect 171826 213058 172062 213294
rect 172146 213058 172382 213294
rect 171826 193058 172062 193294
rect 172146 193058 172382 193294
rect 171826 173058 172062 173294
rect 172146 173058 172382 173294
rect 171826 153058 172062 153294
rect 172146 153058 172382 153294
rect 171826 133058 172062 133294
rect 172146 133058 172382 133294
rect 171826 113058 172062 113294
rect 172146 113058 172382 113294
rect 171826 93058 172062 93294
rect 172146 93058 172382 93294
rect 171826 73058 172062 73294
rect 172146 73058 172382 73294
rect 171826 53058 172062 53294
rect 172146 53058 172382 53294
rect 171826 33058 172062 33294
rect 172146 33058 172382 33294
rect 171826 13058 172062 13294
rect 172146 13058 172382 13294
rect 171826 -1542 172062 -1306
rect 172146 -1542 172382 -1306
rect 171826 -1862 172062 -1626
rect 172146 -1862 172382 -1626
rect 172986 334038 173222 334274
rect 173306 334038 173542 334274
rect 172986 314038 173222 314274
rect 173306 314038 173542 314274
rect 172986 294038 173222 294274
rect 173306 294038 173542 294274
rect 172986 274038 173222 274274
rect 173306 274038 173542 274274
rect 172986 254038 173222 254274
rect 173306 254038 173542 254274
rect 172986 234038 173222 234274
rect 173306 234038 173542 234274
rect 172986 214038 173222 214274
rect 173306 214038 173542 214274
rect 172986 194038 173222 194274
rect 173306 194038 173542 194274
rect 172986 174038 173222 174274
rect 173306 174038 173542 174274
rect 172986 154038 173222 154274
rect 173306 154038 173542 154274
rect 172986 134038 173222 134274
rect 173306 134038 173542 134274
rect 172986 114038 173222 114274
rect 173306 114038 173542 114274
rect 172986 94038 173222 94274
rect 173306 94038 173542 94274
rect 172986 74038 173222 74274
rect 173306 74038 173542 74274
rect 172986 54038 173222 54274
rect 173306 54038 173542 54274
rect 172986 34038 173222 34274
rect 173306 34038 173542 34274
rect 172986 14038 173222 14274
rect 173306 14038 173542 14274
rect 169266 -4422 169502 -4186
rect 169586 -4422 169822 -4186
rect 169266 -4742 169502 -4506
rect 169586 -4742 169822 -4506
rect 162986 -7302 163222 -7066
rect 163306 -7302 163542 -7066
rect 162986 -7622 163222 -7386
rect 163306 -7622 163542 -7386
rect 175546 416718 175782 416954
rect 175866 416718 176102 416954
rect 175546 396718 175782 396954
rect 175866 396718 176102 396954
rect 175546 376718 175782 376954
rect 175866 376718 176102 376954
rect 175546 356718 175782 356954
rect 175866 356718 176102 356954
rect 175546 336718 175782 336954
rect 175866 336718 176102 336954
rect 175546 316718 175782 316954
rect 175866 316718 176102 316954
rect 175546 296718 175782 296954
rect 175866 296718 176102 296954
rect 175546 276718 175782 276954
rect 175866 276718 176102 276954
rect 175546 256718 175782 256954
rect 175866 256718 176102 256954
rect 175546 236718 175782 236954
rect 175866 236718 176102 236954
rect 175546 216718 175782 216954
rect 175866 216718 176102 216954
rect 175546 196718 175782 196954
rect 175866 196718 176102 196954
rect 175546 176718 175782 176954
rect 175866 176718 176102 176954
rect 175546 156718 175782 156954
rect 175866 156718 176102 156954
rect 175546 136718 175782 136954
rect 175866 136718 176102 136954
rect 175546 116718 175782 116954
rect 175866 116718 176102 116954
rect 175546 96718 175782 96954
rect 175866 96718 176102 96954
rect 175546 76718 175782 76954
rect 175866 76718 176102 76954
rect 175546 56718 175782 56954
rect 175866 56718 176102 56954
rect 175546 36718 175782 36954
rect 175866 36718 176102 36954
rect 175546 16718 175782 16954
rect 175866 16718 176102 16954
rect 175546 -3462 175782 -3226
rect 175866 -3462 176102 -3226
rect 175546 -3782 175782 -3546
rect 175866 -3782 176102 -3546
rect 179266 700378 179502 700614
rect 179586 700378 179822 700614
rect 179266 680378 179502 680614
rect 179586 680378 179822 680614
rect 179266 660378 179502 660614
rect 179586 660378 179822 660614
rect 179266 640378 179502 640614
rect 179586 640378 179822 640614
rect 179266 620378 179502 620614
rect 179586 620378 179822 620614
rect 179266 600378 179502 600614
rect 179586 600378 179822 600614
rect 179266 580378 179502 580614
rect 179586 580378 179822 580614
rect 179266 560378 179502 560614
rect 179586 560378 179822 560614
rect 179266 540378 179502 540614
rect 179586 540378 179822 540614
rect 179266 520378 179502 520614
rect 179586 520378 179822 520614
rect 179266 500378 179502 500614
rect 179586 500378 179822 500614
rect 179266 480378 179502 480614
rect 179586 480378 179822 480614
rect 179266 460378 179502 460614
rect 179586 460378 179822 460614
rect 179266 440378 179502 440614
rect 179586 440378 179822 440614
rect 179266 420378 179502 420614
rect 179586 420378 179822 420614
rect 179266 400378 179502 400614
rect 179586 400378 179822 400614
rect 179266 380378 179502 380614
rect 179586 380378 179822 380614
rect 179266 360378 179502 360614
rect 179586 360378 179822 360614
rect 179266 340378 179502 340614
rect 179586 340378 179822 340614
rect 179266 320378 179502 320614
rect 179586 320378 179822 320614
rect 179266 300378 179502 300614
rect 179586 300378 179822 300614
rect 179266 280378 179502 280614
rect 179586 280378 179822 280614
rect 179266 260378 179502 260614
rect 179586 260378 179822 260614
rect 179266 240378 179502 240614
rect 179586 240378 179822 240614
rect 179266 220378 179502 220614
rect 179586 220378 179822 220614
rect 179266 200378 179502 200614
rect 179586 200378 179822 200614
rect 179266 180378 179502 180614
rect 179586 180378 179822 180614
rect 179266 160378 179502 160614
rect 179586 160378 179822 160614
rect 179266 140378 179502 140614
rect 179586 140378 179822 140614
rect 179266 120378 179502 120614
rect 179586 120378 179822 120614
rect 179266 100378 179502 100614
rect 179586 100378 179822 100614
rect 179266 80378 179502 80614
rect 179586 80378 179822 80614
rect 179266 60378 179502 60614
rect 179586 60378 179822 60614
rect 179266 40378 179502 40614
rect 179586 40378 179822 40614
rect 179266 20378 179502 20614
rect 179586 20378 179822 20614
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 683058 182062 683294
rect 182146 683058 182382 683294
rect 181826 663058 182062 663294
rect 182146 663058 182382 663294
rect 181826 643058 182062 643294
rect 182146 643058 182382 643294
rect 181826 623058 182062 623294
rect 182146 623058 182382 623294
rect 181826 603058 182062 603294
rect 182146 603058 182382 603294
rect 181826 583058 182062 583294
rect 182146 583058 182382 583294
rect 181826 563058 182062 563294
rect 182146 563058 182382 563294
rect 181826 543058 182062 543294
rect 182146 543058 182382 543294
rect 181826 523058 182062 523294
rect 182146 523058 182382 523294
rect 181826 503058 182062 503294
rect 182146 503058 182382 503294
rect 181826 483058 182062 483294
rect 182146 483058 182382 483294
rect 181826 463058 182062 463294
rect 182146 463058 182382 463294
rect 181826 443058 182062 443294
rect 182146 443058 182382 443294
rect 181826 423058 182062 423294
rect 182146 423058 182382 423294
rect 181826 403058 182062 403294
rect 182146 403058 182382 403294
rect 181826 383058 182062 383294
rect 182146 383058 182382 383294
rect 181826 363058 182062 363294
rect 182146 363058 182382 363294
rect 181826 343058 182062 343294
rect 182146 343058 182382 343294
rect 181826 323058 182062 323294
rect 182146 323058 182382 323294
rect 181826 303058 182062 303294
rect 182146 303058 182382 303294
rect 181826 283058 182062 283294
rect 182146 283058 182382 283294
rect 181826 263058 182062 263294
rect 182146 263058 182382 263294
rect 181826 243058 182062 243294
rect 182146 243058 182382 243294
rect 181826 223058 182062 223294
rect 182146 223058 182382 223294
rect 181826 203058 182062 203294
rect 182146 203058 182382 203294
rect 181826 183058 182062 183294
rect 182146 183058 182382 183294
rect 181826 163058 182062 163294
rect 182146 163058 182382 163294
rect 181826 143058 182062 143294
rect 182146 143058 182382 143294
rect 181826 123058 182062 123294
rect 182146 123058 182382 123294
rect 181826 103058 182062 103294
rect 182146 103058 182382 103294
rect 181826 83058 182062 83294
rect 182146 83058 182382 83294
rect 181826 63058 182062 63294
rect 182146 63058 182382 63294
rect 181826 43058 182062 43294
rect 182146 43058 182382 43294
rect 181826 23058 182062 23294
rect 182146 23058 182382 23294
rect 181826 3058 182062 3294
rect 182146 3058 182382 3294
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 182986 684038 183222 684274
rect 183306 684038 183542 684274
rect 182986 664038 183222 664274
rect 183306 664038 183542 664274
rect 182986 644038 183222 644274
rect 183306 644038 183542 644274
rect 182986 624038 183222 624274
rect 183306 624038 183542 624274
rect 182986 604038 183222 604274
rect 183306 604038 183542 604274
rect 182986 584038 183222 584274
rect 183306 584038 183542 584274
rect 182986 564038 183222 564274
rect 183306 564038 183542 564274
rect 182986 544038 183222 544274
rect 183306 544038 183542 544274
rect 182986 524038 183222 524274
rect 183306 524038 183542 524274
rect 182986 504038 183222 504274
rect 183306 504038 183542 504274
rect 182986 484038 183222 484274
rect 183306 484038 183542 484274
rect 182986 464038 183222 464274
rect 183306 464038 183542 464274
rect 182986 444038 183222 444274
rect 183306 444038 183542 444274
rect 182986 424038 183222 424274
rect 183306 424038 183542 424274
rect 182986 404038 183222 404274
rect 183306 404038 183542 404274
rect 182986 384038 183222 384274
rect 183306 384038 183542 384274
rect 182986 364038 183222 364274
rect 183306 364038 183542 364274
rect 182986 344038 183222 344274
rect 183306 344038 183542 344274
rect 182986 324038 183222 324274
rect 183306 324038 183542 324274
rect 182986 304038 183222 304274
rect 183306 304038 183542 304274
rect 182986 284038 183222 284274
rect 183306 284038 183542 284274
rect 182986 264038 183222 264274
rect 183306 264038 183542 264274
rect 182986 244038 183222 244274
rect 183306 244038 183542 244274
rect 182986 224038 183222 224274
rect 183306 224038 183542 224274
rect 182986 204038 183222 204274
rect 183306 204038 183542 204274
rect 182986 184038 183222 184274
rect 183306 184038 183542 184274
rect 182986 164038 183222 164274
rect 183306 164038 183542 164274
rect 182986 144038 183222 144274
rect 183306 144038 183542 144274
rect 182986 124038 183222 124274
rect 183306 124038 183542 124274
rect 182986 104038 183222 104274
rect 183306 104038 183542 104274
rect 182986 84038 183222 84274
rect 183306 84038 183542 84274
rect 182986 64038 183222 64274
rect 183306 64038 183542 64274
rect 182986 44038 183222 44274
rect 183306 44038 183542 44274
rect 182986 24038 183222 24274
rect 183306 24038 183542 24274
rect 179266 -5382 179502 -5146
rect 179586 -5382 179822 -5146
rect 179266 -5702 179502 -5466
rect 179586 -5702 179822 -5466
rect 172986 -6342 173222 -6106
rect 173306 -6342 173542 -6106
rect 172986 -6662 173222 -6426
rect 173306 -6662 173542 -6426
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 185546 686718 185782 686954
rect 185866 686718 186102 686954
rect 185546 666718 185782 666954
rect 185866 666718 186102 666954
rect 185546 646718 185782 646954
rect 185866 646718 186102 646954
rect 185546 626718 185782 626954
rect 185866 626718 186102 626954
rect 185546 606718 185782 606954
rect 185866 606718 186102 606954
rect 185546 586718 185782 586954
rect 185866 586718 186102 586954
rect 185546 566718 185782 566954
rect 185866 566718 186102 566954
rect 185546 546718 185782 546954
rect 185866 546718 186102 546954
rect 185546 526718 185782 526954
rect 185866 526718 186102 526954
rect 185546 506718 185782 506954
rect 185866 506718 186102 506954
rect 185546 486718 185782 486954
rect 185866 486718 186102 486954
rect 185546 466718 185782 466954
rect 185866 466718 186102 466954
rect 185546 446718 185782 446954
rect 185866 446718 186102 446954
rect 185546 426718 185782 426954
rect 185866 426718 186102 426954
rect 185546 406718 185782 406954
rect 185866 406718 186102 406954
rect 185546 386718 185782 386954
rect 185866 386718 186102 386954
rect 185546 366718 185782 366954
rect 185866 366718 186102 366954
rect 185546 346718 185782 346954
rect 185866 346718 186102 346954
rect 185546 326718 185782 326954
rect 185866 326718 186102 326954
rect 185546 306718 185782 306954
rect 185866 306718 186102 306954
rect 185546 286718 185782 286954
rect 185866 286718 186102 286954
rect 185546 266718 185782 266954
rect 185866 266718 186102 266954
rect 185546 246718 185782 246954
rect 185866 246718 186102 246954
rect 185546 226718 185782 226954
rect 185866 226718 186102 226954
rect 185546 206718 185782 206954
rect 185866 206718 186102 206954
rect 185546 186718 185782 186954
rect 185866 186718 186102 186954
rect 185546 166718 185782 166954
rect 185866 166718 186102 166954
rect 185546 146718 185782 146954
rect 185866 146718 186102 146954
rect 185546 126718 185782 126954
rect 185866 126718 186102 126954
rect 185546 106718 185782 106954
rect 185866 106718 186102 106954
rect 185546 86718 185782 86954
rect 185866 86718 186102 86954
rect 185546 66718 185782 66954
rect 185866 66718 186102 66954
rect 185546 46718 185782 46954
rect 185866 46718 186102 46954
rect 185546 26718 185782 26954
rect 185866 26718 186102 26954
rect 185546 6718 185782 6954
rect 185866 6718 186102 6954
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 690378 189502 690614
rect 189586 690378 189822 690614
rect 189266 670378 189502 670614
rect 189586 670378 189822 670614
rect 189266 650378 189502 650614
rect 189586 650378 189822 650614
rect 189266 630378 189502 630614
rect 189586 630378 189822 630614
rect 189266 610378 189502 610614
rect 189586 610378 189822 610614
rect 189266 590378 189502 590614
rect 189586 590378 189822 590614
rect 189266 570378 189502 570614
rect 189586 570378 189822 570614
rect 189266 550378 189502 550614
rect 189586 550378 189822 550614
rect 189266 530378 189502 530614
rect 189586 530378 189822 530614
rect 189266 510378 189502 510614
rect 189586 510378 189822 510614
rect 189266 490378 189502 490614
rect 189586 490378 189822 490614
rect 189266 470378 189502 470614
rect 189586 470378 189822 470614
rect 189266 450378 189502 450614
rect 189586 450378 189822 450614
rect 189266 430378 189502 430614
rect 189586 430378 189822 430614
rect 189266 410378 189502 410614
rect 189586 410378 189822 410614
rect 189266 390378 189502 390614
rect 189586 390378 189822 390614
rect 189266 370378 189502 370614
rect 189586 370378 189822 370614
rect 189266 350378 189502 350614
rect 189586 350378 189822 350614
rect 189266 330378 189502 330614
rect 189586 330378 189822 330614
rect 189266 310378 189502 310614
rect 189586 310378 189822 310614
rect 189266 290378 189502 290614
rect 189586 290378 189822 290614
rect 189266 270378 189502 270614
rect 189586 270378 189822 270614
rect 189266 250378 189502 250614
rect 189586 250378 189822 250614
rect 189266 230378 189502 230614
rect 189586 230378 189822 230614
rect 189266 210378 189502 210614
rect 189586 210378 189822 210614
rect 189266 190378 189502 190614
rect 189586 190378 189822 190614
rect 189266 170378 189502 170614
rect 189586 170378 189822 170614
rect 189266 150378 189502 150614
rect 189586 150378 189822 150614
rect 189266 130378 189502 130614
rect 189586 130378 189822 130614
rect 189266 110378 189502 110614
rect 189586 110378 189822 110614
rect 189266 90378 189502 90614
rect 189586 90378 189822 90614
rect 189266 70378 189502 70614
rect 189586 70378 189822 70614
rect 189266 50378 189502 50614
rect 189586 50378 189822 50614
rect 189266 30378 189502 30614
rect 189586 30378 189822 30614
rect 189266 10378 189502 10614
rect 189586 10378 189822 10614
rect 191826 705562 192062 705798
rect 192146 705562 192382 705798
rect 191826 705242 192062 705478
rect 192146 705242 192382 705478
rect 191826 693058 192062 693294
rect 192146 693058 192382 693294
rect 191826 673058 192062 673294
rect 192146 673058 192382 673294
rect 191826 653058 192062 653294
rect 192146 653058 192382 653294
rect 191826 633058 192062 633294
rect 192146 633058 192382 633294
rect 191826 613058 192062 613294
rect 192146 613058 192382 613294
rect 191826 593058 192062 593294
rect 192146 593058 192382 593294
rect 191826 573058 192062 573294
rect 192146 573058 192382 573294
rect 191826 553058 192062 553294
rect 192146 553058 192382 553294
rect 191826 533058 192062 533294
rect 192146 533058 192382 533294
rect 191826 513058 192062 513294
rect 192146 513058 192382 513294
rect 191826 493058 192062 493294
rect 192146 493058 192382 493294
rect 191826 473058 192062 473294
rect 192146 473058 192382 473294
rect 191826 453058 192062 453294
rect 192146 453058 192382 453294
rect 191826 433058 192062 433294
rect 192146 433058 192382 433294
rect 191826 413058 192062 413294
rect 192146 413058 192382 413294
rect 191826 393058 192062 393294
rect 192146 393058 192382 393294
rect 191826 373058 192062 373294
rect 192146 373058 192382 373294
rect 191826 353058 192062 353294
rect 192146 353058 192382 353294
rect 191826 333058 192062 333294
rect 192146 333058 192382 333294
rect 191826 313058 192062 313294
rect 192146 313058 192382 313294
rect 191826 293058 192062 293294
rect 192146 293058 192382 293294
rect 191826 273058 192062 273294
rect 192146 273058 192382 273294
rect 191826 253058 192062 253294
rect 192146 253058 192382 253294
rect 191826 233058 192062 233294
rect 192146 233058 192382 233294
rect 191826 213058 192062 213294
rect 192146 213058 192382 213294
rect 191826 193058 192062 193294
rect 192146 193058 192382 193294
rect 191826 173058 192062 173294
rect 192146 173058 192382 173294
rect 191826 153058 192062 153294
rect 192146 153058 192382 153294
rect 191826 133058 192062 133294
rect 192146 133058 192382 133294
rect 191826 113058 192062 113294
rect 192146 113058 192382 113294
rect 191826 93058 192062 93294
rect 192146 93058 192382 93294
rect 191826 73058 192062 73294
rect 192146 73058 192382 73294
rect 191826 53058 192062 53294
rect 192146 53058 192382 53294
rect 191826 33058 192062 33294
rect 192146 33058 192382 33294
rect 191826 13058 192062 13294
rect 192146 13058 192382 13294
rect 191826 -1542 192062 -1306
rect 192146 -1542 192382 -1306
rect 191826 -1862 192062 -1626
rect 192146 -1862 192382 -1626
rect 202986 711322 203222 711558
rect 203306 711322 203542 711558
rect 202986 711002 203222 711238
rect 203306 711002 203542 711238
rect 199266 709402 199502 709638
rect 199586 709402 199822 709638
rect 199266 709082 199502 709318
rect 199586 709082 199822 709318
rect 192986 694038 193222 694274
rect 193306 694038 193542 694274
rect 192986 674038 193222 674274
rect 193306 674038 193542 674274
rect 192986 654038 193222 654274
rect 193306 654038 193542 654274
rect 192986 634038 193222 634274
rect 193306 634038 193542 634274
rect 192986 614038 193222 614274
rect 193306 614038 193542 614274
rect 192986 594038 193222 594274
rect 193306 594038 193542 594274
rect 192986 574038 193222 574274
rect 193306 574038 193542 574274
rect 192986 554038 193222 554274
rect 193306 554038 193542 554274
rect 192986 534038 193222 534274
rect 193306 534038 193542 534274
rect 192986 514038 193222 514274
rect 193306 514038 193542 514274
rect 192986 494038 193222 494274
rect 193306 494038 193542 494274
rect 192986 474038 193222 474274
rect 193306 474038 193542 474274
rect 192986 454038 193222 454274
rect 193306 454038 193542 454274
rect 192986 434038 193222 434274
rect 193306 434038 193542 434274
rect 192986 414038 193222 414274
rect 193306 414038 193542 414274
rect 192986 394038 193222 394274
rect 193306 394038 193542 394274
rect 192986 374038 193222 374274
rect 193306 374038 193542 374274
rect 192986 354038 193222 354274
rect 193306 354038 193542 354274
rect 192986 334038 193222 334274
rect 193306 334038 193542 334274
rect 192986 314038 193222 314274
rect 193306 314038 193542 314274
rect 192986 294038 193222 294274
rect 193306 294038 193542 294274
rect 192986 274038 193222 274274
rect 193306 274038 193542 274274
rect 192986 254038 193222 254274
rect 193306 254038 193542 254274
rect 192986 234038 193222 234274
rect 193306 234038 193542 234274
rect 192986 214038 193222 214274
rect 193306 214038 193542 214274
rect 192986 194038 193222 194274
rect 193306 194038 193542 194274
rect 192986 174038 193222 174274
rect 193306 174038 193542 174274
rect 192986 154038 193222 154274
rect 193306 154038 193542 154274
rect 192986 134038 193222 134274
rect 193306 134038 193542 134274
rect 192986 114038 193222 114274
rect 193306 114038 193542 114274
rect 192986 94038 193222 94274
rect 193306 94038 193542 94274
rect 192986 74038 193222 74274
rect 193306 74038 193542 74274
rect 192986 54038 193222 54274
rect 193306 54038 193542 54274
rect 192986 34038 193222 34274
rect 193306 34038 193542 34274
rect 192986 14038 193222 14274
rect 193306 14038 193542 14274
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 182986 -7302 183222 -7066
rect 183306 -7302 183542 -7066
rect 182986 -7622 183222 -7386
rect 183306 -7622 183542 -7386
rect 195546 707482 195782 707718
rect 195866 707482 196102 707718
rect 195546 707162 195782 707398
rect 195866 707162 196102 707398
rect 195546 696718 195782 696954
rect 195866 696718 196102 696954
rect 195546 676718 195782 676954
rect 195866 676718 196102 676954
rect 195546 656718 195782 656954
rect 195866 656718 196102 656954
rect 195546 636718 195782 636954
rect 195866 636718 196102 636954
rect 195546 616718 195782 616954
rect 195866 616718 196102 616954
rect 195546 596718 195782 596954
rect 195866 596718 196102 596954
rect 195546 576718 195782 576954
rect 195866 576718 196102 576954
rect 195546 556718 195782 556954
rect 195866 556718 196102 556954
rect 195546 536718 195782 536954
rect 195866 536718 196102 536954
rect 195546 516718 195782 516954
rect 195866 516718 196102 516954
rect 195546 496718 195782 496954
rect 195866 496718 196102 496954
rect 195546 476718 195782 476954
rect 195866 476718 196102 476954
rect 195546 456718 195782 456954
rect 195866 456718 196102 456954
rect 195546 436718 195782 436954
rect 195866 436718 196102 436954
rect 199266 700378 199502 700614
rect 199586 700378 199822 700614
rect 199266 680378 199502 680614
rect 199586 680378 199822 680614
rect 199266 660378 199502 660614
rect 199586 660378 199822 660614
rect 199266 640378 199502 640614
rect 199586 640378 199822 640614
rect 199266 620378 199502 620614
rect 199586 620378 199822 620614
rect 199266 600378 199502 600614
rect 199586 600378 199822 600614
rect 199266 580378 199502 580614
rect 199586 580378 199822 580614
rect 199266 560378 199502 560614
rect 199586 560378 199822 560614
rect 199266 540378 199502 540614
rect 199586 540378 199822 540614
rect 195546 416718 195782 416954
rect 195866 416718 196102 416954
rect 195546 396718 195782 396954
rect 195866 396718 196102 396954
rect 195546 376718 195782 376954
rect 195866 376718 196102 376954
rect 195546 356718 195782 356954
rect 195866 356718 196102 356954
rect 195546 336718 195782 336954
rect 195866 336718 196102 336954
rect 195546 316718 195782 316954
rect 195866 316718 196102 316954
rect 195546 296718 195782 296954
rect 195866 296718 196102 296954
rect 195546 276718 195782 276954
rect 195866 276718 196102 276954
rect 195546 256718 195782 256954
rect 195866 256718 196102 256954
rect 201826 704602 202062 704838
rect 202146 704602 202382 704838
rect 201826 704282 202062 704518
rect 202146 704282 202382 704518
rect 201826 683058 202062 683294
rect 202146 683058 202382 683294
rect 201826 663058 202062 663294
rect 202146 663058 202382 663294
rect 201826 643058 202062 643294
rect 202146 643058 202382 643294
rect 201826 623058 202062 623294
rect 202146 623058 202382 623294
rect 201826 603058 202062 603294
rect 202146 603058 202382 603294
rect 201826 583058 202062 583294
rect 202146 583058 202382 583294
rect 201826 563058 202062 563294
rect 202146 563058 202382 563294
rect 201826 543058 202062 543294
rect 202146 543058 202382 543294
rect 212986 710362 213222 710598
rect 213306 710362 213542 710598
rect 212986 710042 213222 710278
rect 213306 710042 213542 710278
rect 209266 708442 209502 708678
rect 209586 708442 209822 708678
rect 209266 708122 209502 708358
rect 209586 708122 209822 708358
rect 202986 684038 203222 684274
rect 203306 684038 203542 684274
rect 202986 664038 203222 664274
rect 203306 664038 203542 664274
rect 202986 644038 203222 644274
rect 203306 644038 203542 644274
rect 202986 624038 203222 624274
rect 203306 624038 203542 624274
rect 202986 604038 203222 604274
rect 203306 604038 203542 604274
rect 202986 584038 203222 584274
rect 203306 584038 203542 584274
rect 202986 564038 203222 564274
rect 203306 564038 203542 564274
rect 202986 544038 203222 544274
rect 203306 544038 203542 544274
rect 205546 706522 205782 706758
rect 205866 706522 206102 706758
rect 205546 706202 205782 706438
rect 205866 706202 206102 706438
rect 205546 686718 205782 686954
rect 205866 686718 206102 686954
rect 205546 666718 205782 666954
rect 205866 666718 206102 666954
rect 205546 646718 205782 646954
rect 205866 646718 206102 646954
rect 205546 626718 205782 626954
rect 205866 626718 206102 626954
rect 205546 606718 205782 606954
rect 205866 606718 206102 606954
rect 205546 586718 205782 586954
rect 205866 586718 206102 586954
rect 205546 566718 205782 566954
rect 205866 566718 206102 566954
rect 205546 546718 205782 546954
rect 205866 546718 206102 546954
rect 209266 690378 209502 690614
rect 209586 690378 209822 690614
rect 209266 670378 209502 670614
rect 209586 670378 209822 670614
rect 209266 650378 209502 650614
rect 209586 650378 209822 650614
rect 209266 630378 209502 630614
rect 209586 630378 209822 630614
rect 209266 610378 209502 610614
rect 209586 610378 209822 610614
rect 209266 590378 209502 590614
rect 209586 590378 209822 590614
rect 209266 570378 209502 570614
rect 209586 570378 209822 570614
rect 209266 550378 209502 550614
rect 209586 550378 209822 550614
rect 211826 705562 212062 705798
rect 212146 705562 212382 705798
rect 211826 705242 212062 705478
rect 212146 705242 212382 705478
rect 211826 693058 212062 693294
rect 212146 693058 212382 693294
rect 211826 673058 212062 673294
rect 212146 673058 212382 673294
rect 211826 653058 212062 653294
rect 212146 653058 212382 653294
rect 211826 633058 212062 633294
rect 212146 633058 212382 633294
rect 211826 613058 212062 613294
rect 212146 613058 212382 613294
rect 211826 593058 212062 593294
rect 212146 593058 212382 593294
rect 211826 573058 212062 573294
rect 212146 573058 212382 573294
rect 211826 553058 212062 553294
rect 212146 553058 212382 553294
rect 222986 711322 223222 711558
rect 223306 711322 223542 711558
rect 222986 711002 223222 711238
rect 223306 711002 223542 711238
rect 219266 709402 219502 709638
rect 219586 709402 219822 709638
rect 219266 709082 219502 709318
rect 219586 709082 219822 709318
rect 212986 694038 213222 694274
rect 213306 694038 213542 694274
rect 212986 674038 213222 674274
rect 213306 674038 213542 674274
rect 212986 654038 213222 654274
rect 213306 654038 213542 654274
rect 212986 634038 213222 634274
rect 213306 634038 213542 634274
rect 212986 614038 213222 614274
rect 213306 614038 213542 614274
rect 212986 594038 213222 594274
rect 213306 594038 213542 594274
rect 212986 574038 213222 574274
rect 213306 574038 213542 574274
rect 212986 554038 213222 554274
rect 213306 554038 213542 554274
rect 215546 707482 215782 707718
rect 215866 707482 216102 707718
rect 215546 707162 215782 707398
rect 215866 707162 216102 707398
rect 215546 696718 215782 696954
rect 215866 696718 216102 696954
rect 215546 676718 215782 676954
rect 215866 676718 216102 676954
rect 215546 656718 215782 656954
rect 215866 656718 216102 656954
rect 215546 636718 215782 636954
rect 215866 636718 216102 636954
rect 215546 616718 215782 616954
rect 215866 616718 216102 616954
rect 215546 596718 215782 596954
rect 215866 596718 216102 596954
rect 215546 576718 215782 576954
rect 215866 576718 216102 576954
rect 215546 556718 215782 556954
rect 215866 556718 216102 556954
rect 219266 700378 219502 700614
rect 219586 700378 219822 700614
rect 219266 680378 219502 680614
rect 219586 680378 219822 680614
rect 219266 660378 219502 660614
rect 219586 660378 219822 660614
rect 219266 640378 219502 640614
rect 219586 640378 219822 640614
rect 219266 620378 219502 620614
rect 219586 620378 219822 620614
rect 219266 600378 219502 600614
rect 219586 600378 219822 600614
rect 219266 580378 219502 580614
rect 219586 580378 219822 580614
rect 219266 560378 219502 560614
rect 219586 560378 219822 560614
rect 219266 540378 219502 540614
rect 219586 540378 219822 540614
rect 221826 704602 222062 704838
rect 222146 704602 222382 704838
rect 221826 704282 222062 704518
rect 222146 704282 222382 704518
rect 221826 683058 222062 683294
rect 222146 683058 222382 683294
rect 221826 663058 222062 663294
rect 222146 663058 222382 663294
rect 221826 643058 222062 643294
rect 222146 643058 222382 643294
rect 221826 623058 222062 623294
rect 222146 623058 222382 623294
rect 221826 603058 222062 603294
rect 222146 603058 222382 603294
rect 221826 583058 222062 583294
rect 222146 583058 222382 583294
rect 221826 563058 222062 563294
rect 222146 563058 222382 563294
rect 221826 543058 222062 543294
rect 222146 543058 222382 543294
rect 232986 710362 233222 710598
rect 233306 710362 233542 710598
rect 232986 710042 233222 710278
rect 233306 710042 233542 710278
rect 229266 708442 229502 708678
rect 229586 708442 229822 708678
rect 229266 708122 229502 708358
rect 229586 708122 229822 708358
rect 222986 684038 223222 684274
rect 223306 684038 223542 684274
rect 222986 664038 223222 664274
rect 223306 664038 223542 664274
rect 222986 644038 223222 644274
rect 223306 644038 223542 644274
rect 222986 624038 223222 624274
rect 223306 624038 223542 624274
rect 222986 604038 223222 604274
rect 223306 604038 223542 604274
rect 222986 584038 223222 584274
rect 223306 584038 223542 584274
rect 222986 564038 223222 564274
rect 223306 564038 223542 564274
rect 222986 544038 223222 544274
rect 223306 544038 223542 544274
rect 225546 706522 225782 706758
rect 225866 706522 226102 706758
rect 225546 706202 225782 706438
rect 225866 706202 226102 706438
rect 225546 686718 225782 686954
rect 225866 686718 226102 686954
rect 225546 666718 225782 666954
rect 225866 666718 226102 666954
rect 225546 646718 225782 646954
rect 225866 646718 226102 646954
rect 225546 626718 225782 626954
rect 225866 626718 226102 626954
rect 225546 606718 225782 606954
rect 225866 606718 226102 606954
rect 225546 586718 225782 586954
rect 225866 586718 226102 586954
rect 225546 566718 225782 566954
rect 225866 566718 226102 566954
rect 225546 546718 225782 546954
rect 225866 546718 226102 546954
rect 229266 690378 229502 690614
rect 229586 690378 229822 690614
rect 229266 670378 229502 670614
rect 229586 670378 229822 670614
rect 229266 650378 229502 650614
rect 229586 650378 229822 650614
rect 229266 630378 229502 630614
rect 229586 630378 229822 630614
rect 229266 610378 229502 610614
rect 229586 610378 229822 610614
rect 229266 590378 229502 590614
rect 229586 590378 229822 590614
rect 229266 570378 229502 570614
rect 229586 570378 229822 570614
rect 229266 550378 229502 550614
rect 229586 550378 229822 550614
rect 231826 705562 232062 705798
rect 232146 705562 232382 705798
rect 231826 705242 232062 705478
rect 232146 705242 232382 705478
rect 231826 693058 232062 693294
rect 232146 693058 232382 693294
rect 231826 673058 232062 673294
rect 232146 673058 232382 673294
rect 231826 653058 232062 653294
rect 232146 653058 232382 653294
rect 231826 633058 232062 633294
rect 232146 633058 232382 633294
rect 231826 613058 232062 613294
rect 232146 613058 232382 613294
rect 231826 593058 232062 593294
rect 232146 593058 232382 593294
rect 231826 573058 232062 573294
rect 232146 573058 232382 573294
rect 231826 553058 232062 553294
rect 232146 553058 232382 553294
rect 242986 711322 243222 711558
rect 243306 711322 243542 711558
rect 242986 711002 243222 711238
rect 243306 711002 243542 711238
rect 239266 709402 239502 709638
rect 239586 709402 239822 709638
rect 239266 709082 239502 709318
rect 239586 709082 239822 709318
rect 232986 694038 233222 694274
rect 233306 694038 233542 694274
rect 232986 674038 233222 674274
rect 233306 674038 233542 674274
rect 232986 654038 233222 654274
rect 233306 654038 233542 654274
rect 232986 634038 233222 634274
rect 233306 634038 233542 634274
rect 232986 614038 233222 614274
rect 233306 614038 233542 614274
rect 232986 594038 233222 594274
rect 233306 594038 233542 594274
rect 232986 574038 233222 574274
rect 233306 574038 233542 574274
rect 232986 554038 233222 554274
rect 233306 554038 233542 554274
rect 235546 707482 235782 707718
rect 235866 707482 236102 707718
rect 235546 707162 235782 707398
rect 235866 707162 236102 707398
rect 235546 696718 235782 696954
rect 235866 696718 236102 696954
rect 235546 676718 235782 676954
rect 235866 676718 236102 676954
rect 239266 700378 239502 700614
rect 239586 700378 239822 700614
rect 239266 680378 239502 680614
rect 239586 680378 239822 680614
rect 239266 660378 239502 660614
rect 239586 660378 239822 660614
rect 241826 704602 242062 704838
rect 242146 704602 242382 704838
rect 241826 704282 242062 704518
rect 242146 704282 242382 704518
rect 241826 683058 242062 683294
rect 242146 683058 242382 683294
rect 241826 663058 242062 663294
rect 242146 663058 242382 663294
rect 252986 710362 253222 710598
rect 253306 710362 253542 710598
rect 252986 710042 253222 710278
rect 253306 710042 253542 710278
rect 249266 708442 249502 708678
rect 249586 708442 249822 708678
rect 249266 708122 249502 708358
rect 249586 708122 249822 708358
rect 242986 684038 243222 684274
rect 243306 684038 243542 684274
rect 242986 664038 243222 664274
rect 243306 664038 243542 664274
rect 245546 706522 245782 706758
rect 245866 706522 246102 706758
rect 245546 706202 245782 706438
rect 245866 706202 246102 706438
rect 245546 686718 245782 686954
rect 245866 686718 246102 686954
rect 245546 666718 245782 666954
rect 245866 666718 246102 666954
rect 249266 690378 249502 690614
rect 249586 690378 249822 690614
rect 249266 670378 249502 670614
rect 249586 670378 249822 670614
rect 251826 705562 252062 705798
rect 252146 705562 252382 705798
rect 251826 705242 252062 705478
rect 252146 705242 252382 705478
rect 251826 693058 252062 693294
rect 252146 693058 252382 693294
rect 251826 673058 252062 673294
rect 252146 673058 252382 673294
rect 262986 711322 263222 711558
rect 263306 711322 263542 711558
rect 262986 711002 263222 711238
rect 263306 711002 263542 711238
rect 259266 709402 259502 709638
rect 259586 709402 259822 709638
rect 259266 709082 259502 709318
rect 259586 709082 259822 709318
rect 252986 694038 253222 694274
rect 253306 694038 253542 694274
rect 252986 674038 253222 674274
rect 253306 674038 253542 674274
rect 255546 707482 255782 707718
rect 255866 707482 256102 707718
rect 255546 707162 255782 707398
rect 255866 707162 256102 707398
rect 255546 696718 255782 696954
rect 255866 696718 256102 696954
rect 255546 676718 255782 676954
rect 255866 676718 256102 676954
rect 259266 700378 259502 700614
rect 259586 700378 259822 700614
rect 259266 680378 259502 680614
rect 259586 680378 259822 680614
rect 259266 660378 259502 660614
rect 259586 660378 259822 660614
rect 261826 704602 262062 704838
rect 262146 704602 262382 704838
rect 261826 704282 262062 704518
rect 262146 704282 262382 704518
rect 261826 683058 262062 683294
rect 262146 683058 262382 683294
rect 261826 663058 262062 663294
rect 262146 663058 262382 663294
rect 272986 710362 273222 710598
rect 273306 710362 273542 710598
rect 272986 710042 273222 710278
rect 273306 710042 273542 710278
rect 269266 708442 269502 708678
rect 269586 708442 269822 708678
rect 269266 708122 269502 708358
rect 269586 708122 269822 708358
rect 262986 684038 263222 684274
rect 263306 684038 263542 684274
rect 262986 664038 263222 664274
rect 263306 664038 263542 664274
rect 265546 706522 265782 706758
rect 265866 706522 266102 706758
rect 265546 706202 265782 706438
rect 265866 706202 266102 706438
rect 265546 686718 265782 686954
rect 265866 686718 266102 686954
rect 265546 666718 265782 666954
rect 265866 666718 266102 666954
rect 269266 690378 269502 690614
rect 269586 690378 269822 690614
rect 269266 670378 269502 670614
rect 269586 670378 269822 670614
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 693058 272062 693294
rect 272146 693058 272382 693294
rect 271826 673058 272062 673294
rect 272146 673058 272382 673294
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 272986 694038 273222 694274
rect 273306 694038 273542 694274
rect 272986 674038 273222 674274
rect 273306 674038 273542 674274
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 275546 696718 275782 696954
rect 275866 696718 276102 696954
rect 275546 676718 275782 676954
rect 275866 676718 276102 676954
rect 279266 700378 279502 700614
rect 279586 700378 279822 700614
rect 279266 680378 279502 680614
rect 279586 680378 279822 680614
rect 279266 660378 279502 660614
rect 279586 660378 279822 660614
rect 281826 704602 282062 704838
rect 282146 704602 282382 704838
rect 281826 704282 282062 704518
rect 282146 704282 282382 704518
rect 281826 683058 282062 683294
rect 282146 683058 282382 683294
rect 281826 663058 282062 663294
rect 282146 663058 282382 663294
rect 292986 710362 293222 710598
rect 293306 710362 293542 710598
rect 292986 710042 293222 710278
rect 293306 710042 293542 710278
rect 289266 708442 289502 708678
rect 289586 708442 289822 708678
rect 289266 708122 289502 708358
rect 289586 708122 289822 708358
rect 282986 684038 283222 684274
rect 283306 684038 283542 684274
rect 282986 664038 283222 664274
rect 283306 664038 283542 664274
rect 285546 706522 285782 706758
rect 285866 706522 286102 706758
rect 285546 706202 285782 706438
rect 285866 706202 286102 706438
rect 285546 686718 285782 686954
rect 285866 686718 286102 686954
rect 285546 666718 285782 666954
rect 285866 666718 286102 666954
rect 289266 690378 289502 690614
rect 289586 690378 289822 690614
rect 289266 670378 289502 670614
rect 289586 670378 289822 670614
rect 291826 705562 292062 705798
rect 292146 705562 292382 705798
rect 291826 705242 292062 705478
rect 292146 705242 292382 705478
rect 291826 693058 292062 693294
rect 292146 693058 292382 693294
rect 291826 673058 292062 673294
rect 292146 673058 292382 673294
rect 302986 711322 303222 711558
rect 303306 711322 303542 711558
rect 302986 711002 303222 711238
rect 303306 711002 303542 711238
rect 299266 709402 299502 709638
rect 299586 709402 299822 709638
rect 299266 709082 299502 709318
rect 299586 709082 299822 709318
rect 292986 694038 293222 694274
rect 293306 694038 293542 694274
rect 292986 674038 293222 674274
rect 293306 674038 293542 674274
rect 295546 707482 295782 707718
rect 295866 707482 296102 707718
rect 295546 707162 295782 707398
rect 295866 707162 296102 707398
rect 295546 696718 295782 696954
rect 295866 696718 296102 696954
rect 295546 676718 295782 676954
rect 295866 676718 296102 676954
rect 299266 700378 299502 700614
rect 299586 700378 299822 700614
rect 299266 680378 299502 680614
rect 299586 680378 299822 680614
rect 299266 660378 299502 660614
rect 299586 660378 299822 660614
rect 301826 704602 302062 704838
rect 302146 704602 302382 704838
rect 301826 704282 302062 704518
rect 302146 704282 302382 704518
rect 301826 683058 302062 683294
rect 302146 683058 302382 683294
rect 301826 663058 302062 663294
rect 302146 663058 302382 663294
rect 312986 710362 313222 710598
rect 313306 710362 313542 710598
rect 312986 710042 313222 710278
rect 313306 710042 313542 710278
rect 309266 708442 309502 708678
rect 309586 708442 309822 708678
rect 309266 708122 309502 708358
rect 309586 708122 309822 708358
rect 302986 684038 303222 684274
rect 303306 684038 303542 684274
rect 302986 664038 303222 664274
rect 303306 664038 303542 664274
rect 305546 706522 305782 706758
rect 305866 706522 306102 706758
rect 305546 706202 305782 706438
rect 305866 706202 306102 706438
rect 305546 686718 305782 686954
rect 305866 686718 306102 686954
rect 305546 666718 305782 666954
rect 305866 666718 306102 666954
rect 309266 690378 309502 690614
rect 309586 690378 309822 690614
rect 309266 670378 309502 670614
rect 309586 670378 309822 670614
rect 311826 705562 312062 705798
rect 312146 705562 312382 705798
rect 311826 705242 312062 705478
rect 312146 705242 312382 705478
rect 311826 693058 312062 693294
rect 312146 693058 312382 693294
rect 311826 673058 312062 673294
rect 312146 673058 312382 673294
rect 322986 711322 323222 711558
rect 323306 711322 323542 711558
rect 322986 711002 323222 711238
rect 323306 711002 323542 711238
rect 319266 709402 319502 709638
rect 319586 709402 319822 709638
rect 319266 709082 319502 709318
rect 319586 709082 319822 709318
rect 312986 694038 313222 694274
rect 313306 694038 313542 694274
rect 312986 674038 313222 674274
rect 313306 674038 313542 674274
rect 315546 707482 315782 707718
rect 315866 707482 316102 707718
rect 315546 707162 315782 707398
rect 315866 707162 316102 707398
rect 315546 696718 315782 696954
rect 315866 696718 316102 696954
rect 315546 676718 315782 676954
rect 315866 676718 316102 676954
rect 319266 700378 319502 700614
rect 319586 700378 319822 700614
rect 319266 680378 319502 680614
rect 319586 680378 319822 680614
rect 319266 660378 319502 660614
rect 319586 660378 319822 660614
rect 321826 704602 322062 704838
rect 322146 704602 322382 704838
rect 321826 704282 322062 704518
rect 322146 704282 322382 704518
rect 321826 683058 322062 683294
rect 322146 683058 322382 683294
rect 321826 663058 322062 663294
rect 322146 663058 322382 663294
rect 332986 710362 333222 710598
rect 333306 710362 333542 710598
rect 332986 710042 333222 710278
rect 333306 710042 333542 710278
rect 329266 708442 329502 708678
rect 329586 708442 329822 708678
rect 329266 708122 329502 708358
rect 329586 708122 329822 708358
rect 322986 684038 323222 684274
rect 323306 684038 323542 684274
rect 322986 664038 323222 664274
rect 323306 664038 323542 664274
rect 325546 706522 325782 706758
rect 325866 706522 326102 706758
rect 325546 706202 325782 706438
rect 325866 706202 326102 706438
rect 325546 686718 325782 686954
rect 325866 686718 326102 686954
rect 325546 666718 325782 666954
rect 325866 666718 326102 666954
rect 329266 690378 329502 690614
rect 329586 690378 329822 690614
rect 329266 670378 329502 670614
rect 329586 670378 329822 670614
rect 331826 705562 332062 705798
rect 332146 705562 332382 705798
rect 331826 705242 332062 705478
rect 332146 705242 332382 705478
rect 331826 693058 332062 693294
rect 332146 693058 332382 693294
rect 331826 673058 332062 673294
rect 332146 673058 332382 673294
rect 342986 711322 343222 711558
rect 343306 711322 343542 711558
rect 342986 711002 343222 711238
rect 343306 711002 343542 711238
rect 339266 709402 339502 709638
rect 339586 709402 339822 709638
rect 339266 709082 339502 709318
rect 339586 709082 339822 709318
rect 332986 694038 333222 694274
rect 333306 694038 333542 694274
rect 332986 674038 333222 674274
rect 333306 674038 333542 674274
rect 335546 707482 335782 707718
rect 335866 707482 336102 707718
rect 335546 707162 335782 707398
rect 335866 707162 336102 707398
rect 335546 696718 335782 696954
rect 335866 696718 336102 696954
rect 335546 676718 335782 676954
rect 335866 676718 336102 676954
rect 339266 700378 339502 700614
rect 339586 700378 339822 700614
rect 339266 680378 339502 680614
rect 339586 680378 339822 680614
rect 339266 660378 339502 660614
rect 339586 660378 339822 660614
rect 235546 656718 235782 656954
rect 235866 656718 236102 656954
rect 240328 653058 240564 653294
rect 335392 653058 335628 653294
rect 241008 643058 241244 643294
rect 334712 643058 334948 643294
rect 235546 636718 235782 636954
rect 235866 636718 236102 636954
rect 341826 704602 342062 704838
rect 342146 704602 342382 704838
rect 341826 704282 342062 704518
rect 342146 704282 342382 704518
rect 341826 683058 342062 683294
rect 342146 683058 342382 683294
rect 341826 663058 342062 663294
rect 342146 663058 342382 663294
rect 339266 640378 339502 640614
rect 339586 640378 339822 640614
rect 240328 633058 240564 633294
rect 335392 633058 335628 633294
rect 241008 623058 241244 623294
rect 334712 623058 334948 623294
rect 235546 616718 235782 616954
rect 235866 616718 236102 616954
rect 339266 620378 339502 620614
rect 339586 620378 339822 620614
rect 240328 613058 240564 613294
rect 335392 613058 335628 613294
rect 241008 603058 241244 603294
rect 334712 603058 334948 603294
rect 235546 596718 235782 596954
rect 235866 596718 236102 596954
rect 240328 593058 240564 593294
rect 335392 593058 335628 593294
rect 241008 583058 241244 583294
rect 334712 583058 334948 583294
rect 235546 576718 235782 576954
rect 235866 576718 236102 576954
rect 235546 556718 235782 556954
rect 235866 556718 236102 556954
rect 239266 560378 239502 560614
rect 239586 560378 239822 560614
rect 239266 540378 239502 540614
rect 239586 540378 239822 540614
rect 241826 563058 242062 563294
rect 242146 563058 242382 563294
rect 241826 543058 242062 543294
rect 242146 543058 242382 543294
rect 242986 564038 243222 564274
rect 243306 564038 243542 564274
rect 242986 544038 243222 544274
rect 243306 544038 243542 544274
rect 245546 566718 245782 566954
rect 245866 566718 246102 566954
rect 245546 546718 245782 546954
rect 245866 546718 246102 546954
rect 249266 570378 249502 570614
rect 249586 570378 249822 570614
rect 249266 550378 249502 550614
rect 249586 550378 249822 550614
rect 251826 573058 252062 573294
rect 252146 573058 252382 573294
rect 251826 553058 252062 553294
rect 252146 553058 252382 553294
rect 252986 574038 253222 574274
rect 253306 574038 253542 574274
rect 252986 554038 253222 554274
rect 253306 554038 253542 554274
rect 255546 556718 255782 556954
rect 255866 556718 256102 556954
rect 259266 560378 259502 560614
rect 259586 560378 259822 560614
rect 259266 540378 259502 540614
rect 259586 540378 259822 540614
rect 261826 563058 262062 563294
rect 262146 563058 262382 563294
rect 261826 543058 262062 543294
rect 262146 543058 262382 543294
rect 262986 564038 263222 564274
rect 263306 564038 263542 564274
rect 262986 544038 263222 544274
rect 263306 544038 263542 544274
rect 265546 566718 265782 566954
rect 265866 566718 266102 566954
rect 265546 546718 265782 546954
rect 265866 546718 266102 546954
rect 269266 570378 269502 570614
rect 269586 570378 269822 570614
rect 269266 550378 269502 550614
rect 269586 550378 269822 550614
rect 271826 573058 272062 573294
rect 272146 573058 272382 573294
rect 271826 553058 272062 553294
rect 272146 553058 272382 553294
rect 272986 574038 273222 574274
rect 273306 574038 273542 574274
rect 272986 554038 273222 554274
rect 273306 554038 273542 554274
rect 275546 556718 275782 556954
rect 275866 556718 276102 556954
rect 279266 560378 279502 560614
rect 279586 560378 279822 560614
rect 279266 540378 279502 540614
rect 279586 540378 279822 540614
rect 281826 563058 282062 563294
rect 282146 563058 282382 563294
rect 281826 543058 282062 543294
rect 282146 543058 282382 543294
rect 282986 564038 283222 564274
rect 283306 564038 283542 564274
rect 282986 544038 283222 544274
rect 283306 544038 283542 544274
rect 285546 566718 285782 566954
rect 285866 566718 286102 566954
rect 285546 546718 285782 546954
rect 285866 546718 286102 546954
rect 289266 570378 289502 570614
rect 289586 570378 289822 570614
rect 289266 550378 289502 550614
rect 289586 550378 289822 550614
rect 291826 573058 292062 573294
rect 292146 573058 292382 573294
rect 291826 553058 292062 553294
rect 292146 553058 292382 553294
rect 292986 574038 293222 574274
rect 293306 574038 293542 574274
rect 292986 554038 293222 554274
rect 293306 554038 293542 554274
rect 295546 556718 295782 556954
rect 295866 556718 296102 556954
rect 299266 560378 299502 560614
rect 299586 560378 299822 560614
rect 299266 540378 299502 540614
rect 299586 540378 299822 540614
rect 301826 563058 302062 563294
rect 302146 563058 302382 563294
rect 301826 543058 302062 543294
rect 302146 543058 302382 543294
rect 302986 564038 303222 564274
rect 303306 564038 303542 564274
rect 302986 544038 303222 544274
rect 303306 544038 303542 544274
rect 305546 566718 305782 566954
rect 305866 566718 306102 566954
rect 305546 546718 305782 546954
rect 305866 546718 306102 546954
rect 309266 570378 309502 570614
rect 309586 570378 309822 570614
rect 309266 550378 309502 550614
rect 309586 550378 309822 550614
rect 311826 573058 312062 573294
rect 312146 573058 312382 573294
rect 311826 553058 312062 553294
rect 312146 553058 312382 553294
rect 312986 574038 313222 574274
rect 313306 574038 313542 574274
rect 312986 554038 313222 554274
rect 313306 554038 313542 554274
rect 315546 556718 315782 556954
rect 315866 556718 316102 556954
rect 319266 560378 319502 560614
rect 319586 560378 319822 560614
rect 319266 540378 319502 540614
rect 319586 540378 319822 540614
rect 321826 563058 322062 563294
rect 322146 563058 322382 563294
rect 321826 543058 322062 543294
rect 322146 543058 322382 543294
rect 322986 564038 323222 564274
rect 323306 564038 323542 564274
rect 322986 544038 323222 544274
rect 323306 544038 323542 544274
rect 325546 566718 325782 566954
rect 325866 566718 326102 566954
rect 325546 546718 325782 546954
rect 325866 546718 326102 546954
rect 329266 570378 329502 570614
rect 329586 570378 329822 570614
rect 329266 550378 329502 550614
rect 329586 550378 329822 550614
rect 331826 573058 332062 573294
rect 332146 573058 332382 573294
rect 331826 553058 332062 553294
rect 332146 553058 332382 553294
rect 332986 574038 333222 574274
rect 333306 574038 333542 574274
rect 332986 554038 333222 554274
rect 333306 554038 333542 554274
rect 335546 556718 335782 556954
rect 335866 556718 336102 556954
rect 200328 533058 200564 533294
rect 336056 533058 336292 533294
rect 201008 523058 201244 523294
rect 335376 523058 335612 523294
rect 200328 513058 200564 513294
rect 336056 513058 336292 513294
rect 201008 503058 201244 503294
rect 335376 503058 335612 503294
rect 200328 493058 200564 493294
rect 336056 493058 336292 493294
rect 201008 483058 201244 483294
rect 335376 483058 335612 483294
rect 200328 473058 200564 473294
rect 336056 473058 336292 473294
rect 201008 463058 201244 463294
rect 335376 463058 335612 463294
rect 199266 440378 199502 440614
rect 199586 440378 199822 440614
rect 201826 443058 202062 443294
rect 202146 443058 202382 443294
rect 201826 423058 202062 423294
rect 202146 423058 202382 423294
rect 202986 444038 203222 444274
rect 203306 444038 203542 444274
rect 202986 424038 203222 424274
rect 203306 424038 203542 424274
rect 205546 446718 205782 446954
rect 205866 446718 206102 446954
rect 205546 426718 205782 426954
rect 205866 426718 206102 426954
rect 209266 450378 209502 450614
rect 209586 450378 209822 450614
rect 209266 430378 209502 430614
rect 209586 430378 209822 430614
rect 211826 433058 212062 433294
rect 212146 433058 212382 433294
rect 212986 434038 213222 434274
rect 213306 434038 213542 434274
rect 215546 436718 215782 436954
rect 215866 436718 216102 436954
rect 219266 440378 219502 440614
rect 219586 440378 219822 440614
rect 221826 443058 222062 443294
rect 222146 443058 222382 443294
rect 221826 423058 222062 423294
rect 222146 423058 222382 423294
rect 222986 444038 223222 444274
rect 223306 444038 223542 444274
rect 222986 424038 223222 424274
rect 223306 424038 223542 424274
rect 225546 446718 225782 446954
rect 225866 446718 226102 446954
rect 225546 426718 225782 426954
rect 225866 426718 226102 426954
rect 229266 450378 229502 450614
rect 229586 450378 229822 450614
rect 229266 430378 229502 430614
rect 229586 430378 229822 430614
rect 231826 433058 232062 433294
rect 232146 433058 232382 433294
rect 232986 434038 233222 434274
rect 233306 434038 233542 434274
rect 235546 436718 235782 436954
rect 235866 436718 236102 436954
rect 239266 440378 239502 440614
rect 239586 440378 239822 440614
rect 241826 443058 242062 443294
rect 242146 443058 242382 443294
rect 241826 423058 242062 423294
rect 242146 423058 242382 423294
rect 242986 444038 243222 444274
rect 243306 444038 243542 444274
rect 242986 424038 243222 424274
rect 243306 424038 243542 424274
rect 245546 446718 245782 446954
rect 245866 446718 246102 446954
rect 245546 426718 245782 426954
rect 245866 426718 246102 426954
rect 249266 450378 249502 450614
rect 249586 450378 249822 450614
rect 249266 430378 249502 430614
rect 249586 430378 249822 430614
rect 251826 433058 252062 433294
rect 252146 433058 252382 433294
rect 252986 434038 253222 434274
rect 253306 434038 253542 434274
rect 255546 436718 255782 436954
rect 255866 436718 256102 436954
rect 259266 440378 259502 440614
rect 259586 440378 259822 440614
rect 261826 443058 262062 443294
rect 262146 443058 262382 443294
rect 261826 423058 262062 423294
rect 262146 423058 262382 423294
rect 262986 444038 263222 444274
rect 263306 444038 263542 444274
rect 262986 424038 263222 424274
rect 263306 424038 263542 424274
rect 265546 446718 265782 446954
rect 265866 446718 266102 446954
rect 265546 426718 265782 426954
rect 265866 426718 266102 426954
rect 269266 450378 269502 450614
rect 269586 450378 269822 450614
rect 269266 430378 269502 430614
rect 269586 430378 269822 430614
rect 271826 433058 272062 433294
rect 272146 433058 272382 433294
rect 272986 434038 273222 434274
rect 273306 434038 273542 434274
rect 275546 436718 275782 436954
rect 275866 436718 276102 436954
rect 279266 440378 279502 440614
rect 279586 440378 279822 440614
rect 281826 443058 282062 443294
rect 282146 443058 282382 443294
rect 281826 423058 282062 423294
rect 282146 423058 282382 423294
rect 282986 444038 283222 444274
rect 283306 444038 283542 444274
rect 282986 424038 283222 424274
rect 283306 424038 283542 424274
rect 285546 446718 285782 446954
rect 285866 446718 286102 446954
rect 285546 426718 285782 426954
rect 285866 426718 286102 426954
rect 289266 450378 289502 450614
rect 289586 450378 289822 450614
rect 289266 430378 289502 430614
rect 289586 430378 289822 430614
rect 291826 433058 292062 433294
rect 292146 433058 292382 433294
rect 292986 434038 293222 434274
rect 293306 434038 293542 434274
rect 295546 436718 295782 436954
rect 295866 436718 296102 436954
rect 299266 440378 299502 440614
rect 299586 440378 299822 440614
rect 301826 443058 302062 443294
rect 302146 443058 302382 443294
rect 301826 423058 302062 423294
rect 302146 423058 302382 423294
rect 302986 444038 303222 444274
rect 303306 444038 303542 444274
rect 302986 424038 303222 424274
rect 303306 424038 303542 424274
rect 305546 446718 305782 446954
rect 305866 446718 306102 446954
rect 305546 426718 305782 426954
rect 305866 426718 306102 426954
rect 309266 450378 309502 450614
rect 309586 450378 309822 450614
rect 309266 430378 309502 430614
rect 309586 430378 309822 430614
rect 311826 433058 312062 433294
rect 312146 433058 312382 433294
rect 312986 434038 313222 434274
rect 313306 434038 313542 434274
rect 315546 436718 315782 436954
rect 315866 436718 316102 436954
rect 319266 440378 319502 440614
rect 319586 440378 319822 440614
rect 321826 443058 322062 443294
rect 322146 443058 322382 443294
rect 321826 423058 322062 423294
rect 322146 423058 322382 423294
rect 322986 444038 323222 444274
rect 323306 444038 323542 444274
rect 322986 424038 323222 424274
rect 323306 424038 323542 424274
rect 325546 446718 325782 446954
rect 325866 446718 326102 446954
rect 325546 426718 325782 426954
rect 325866 426718 326102 426954
rect 329266 450378 329502 450614
rect 329586 450378 329822 450614
rect 329266 430378 329502 430614
rect 329586 430378 329822 430614
rect 331826 433058 332062 433294
rect 332146 433058 332382 433294
rect 332986 434038 333222 434274
rect 333306 434038 333542 434274
rect 335546 436718 335782 436954
rect 335866 436718 336102 436954
rect 339266 600378 339502 600614
rect 339586 600378 339822 600614
rect 339266 580378 339502 580614
rect 339586 580378 339822 580614
rect 339266 560378 339502 560614
rect 339586 560378 339822 560614
rect 339266 540378 339502 540614
rect 339586 540378 339822 540614
rect 339266 520378 339502 520614
rect 339586 520378 339822 520614
rect 339266 500378 339502 500614
rect 339586 500378 339822 500614
rect 339266 480378 339502 480614
rect 339586 480378 339822 480614
rect 339266 460378 339502 460614
rect 339586 460378 339822 460614
rect 339266 440378 339502 440614
rect 339586 440378 339822 440614
rect 341826 643058 342062 643294
rect 342146 643058 342382 643294
rect 341826 623058 342062 623294
rect 342146 623058 342382 623294
rect 341826 603058 342062 603294
rect 342146 603058 342382 603294
rect 341826 583058 342062 583294
rect 342146 583058 342382 583294
rect 341826 563058 342062 563294
rect 342146 563058 342382 563294
rect 341826 543058 342062 543294
rect 342146 543058 342382 543294
rect 341826 523058 342062 523294
rect 342146 523058 342382 523294
rect 341826 503058 342062 503294
rect 342146 503058 342382 503294
rect 341826 483058 342062 483294
rect 342146 483058 342382 483294
rect 341826 463058 342062 463294
rect 342146 463058 342382 463294
rect 341826 443058 342062 443294
rect 342146 443058 342382 443294
rect 341826 423058 342062 423294
rect 342146 423058 342382 423294
rect 352986 710362 353222 710598
rect 353306 710362 353542 710598
rect 352986 710042 353222 710278
rect 353306 710042 353542 710278
rect 349266 708442 349502 708678
rect 349586 708442 349822 708678
rect 349266 708122 349502 708358
rect 349586 708122 349822 708358
rect 342986 684038 343222 684274
rect 343306 684038 343542 684274
rect 342986 664038 343222 664274
rect 343306 664038 343542 664274
rect 342986 644038 343222 644274
rect 343306 644038 343542 644274
rect 342986 624038 343222 624274
rect 343306 624038 343542 624274
rect 342986 604038 343222 604274
rect 343306 604038 343542 604274
rect 342986 584038 343222 584274
rect 343306 584038 343542 584274
rect 342986 564038 343222 564274
rect 343306 564038 343542 564274
rect 342986 544038 343222 544274
rect 343306 544038 343542 544274
rect 342986 524038 343222 524274
rect 343306 524038 343542 524274
rect 342986 504038 343222 504274
rect 343306 504038 343542 504274
rect 342986 484038 343222 484274
rect 343306 484038 343542 484274
rect 342986 464038 343222 464274
rect 343306 464038 343542 464274
rect 342986 444038 343222 444274
rect 343306 444038 343542 444274
rect 342986 424038 343222 424274
rect 343306 424038 343542 424274
rect 345546 706522 345782 706758
rect 345866 706522 346102 706758
rect 345546 706202 345782 706438
rect 345866 706202 346102 706438
rect 345546 686718 345782 686954
rect 345866 686718 346102 686954
rect 345546 666718 345782 666954
rect 345866 666718 346102 666954
rect 345546 646718 345782 646954
rect 345866 646718 346102 646954
rect 345546 626718 345782 626954
rect 345866 626718 346102 626954
rect 345546 606718 345782 606954
rect 345866 606718 346102 606954
rect 345546 586718 345782 586954
rect 345866 586718 346102 586954
rect 345546 566718 345782 566954
rect 345866 566718 346102 566954
rect 345546 546718 345782 546954
rect 345866 546718 346102 546954
rect 345546 526718 345782 526954
rect 345866 526718 346102 526954
rect 345546 506718 345782 506954
rect 345866 506718 346102 506954
rect 345546 486718 345782 486954
rect 345866 486718 346102 486954
rect 345546 466718 345782 466954
rect 345866 466718 346102 466954
rect 345546 446718 345782 446954
rect 345866 446718 346102 446954
rect 345546 426718 345782 426954
rect 345866 426718 346102 426954
rect 349266 690378 349502 690614
rect 349586 690378 349822 690614
rect 349266 670378 349502 670614
rect 349586 670378 349822 670614
rect 349266 650378 349502 650614
rect 349586 650378 349822 650614
rect 349266 630378 349502 630614
rect 349586 630378 349822 630614
rect 349266 610378 349502 610614
rect 349586 610378 349822 610614
rect 349266 590378 349502 590614
rect 349586 590378 349822 590614
rect 349266 570378 349502 570614
rect 349586 570378 349822 570614
rect 349266 550378 349502 550614
rect 349586 550378 349822 550614
rect 349266 530378 349502 530614
rect 349586 530378 349822 530614
rect 349266 510378 349502 510614
rect 349586 510378 349822 510614
rect 349266 490378 349502 490614
rect 349586 490378 349822 490614
rect 349266 470378 349502 470614
rect 349586 470378 349822 470614
rect 349266 450378 349502 450614
rect 349586 450378 349822 450614
rect 349266 430378 349502 430614
rect 349586 430378 349822 430614
rect 351826 705562 352062 705798
rect 352146 705562 352382 705798
rect 351826 705242 352062 705478
rect 352146 705242 352382 705478
rect 351826 693058 352062 693294
rect 352146 693058 352382 693294
rect 351826 673058 352062 673294
rect 352146 673058 352382 673294
rect 351826 653058 352062 653294
rect 352146 653058 352382 653294
rect 351826 633058 352062 633294
rect 352146 633058 352382 633294
rect 351826 613058 352062 613294
rect 352146 613058 352382 613294
rect 351826 593058 352062 593294
rect 352146 593058 352382 593294
rect 351826 573058 352062 573294
rect 352146 573058 352382 573294
rect 351826 553058 352062 553294
rect 352146 553058 352382 553294
rect 351826 533058 352062 533294
rect 352146 533058 352382 533294
rect 351826 513058 352062 513294
rect 352146 513058 352382 513294
rect 351826 493058 352062 493294
rect 352146 493058 352382 493294
rect 351826 473058 352062 473294
rect 352146 473058 352382 473294
rect 351826 453058 352062 453294
rect 352146 453058 352382 453294
rect 351826 433058 352062 433294
rect 352146 433058 352382 433294
rect 362986 711322 363222 711558
rect 363306 711322 363542 711558
rect 362986 711002 363222 711238
rect 363306 711002 363542 711238
rect 359266 709402 359502 709638
rect 359586 709402 359822 709638
rect 359266 709082 359502 709318
rect 359586 709082 359822 709318
rect 352986 694038 353222 694274
rect 353306 694038 353542 694274
rect 352986 674038 353222 674274
rect 353306 674038 353542 674274
rect 352986 654038 353222 654274
rect 353306 654038 353542 654274
rect 352986 634038 353222 634274
rect 353306 634038 353542 634274
rect 352986 614038 353222 614274
rect 353306 614038 353542 614274
rect 352986 594038 353222 594274
rect 353306 594038 353542 594274
rect 352986 574038 353222 574274
rect 353306 574038 353542 574274
rect 352986 554038 353222 554274
rect 353306 554038 353542 554274
rect 352986 534038 353222 534274
rect 353306 534038 353542 534274
rect 352986 514038 353222 514274
rect 353306 514038 353542 514274
rect 352986 494038 353222 494274
rect 353306 494038 353542 494274
rect 352986 474038 353222 474274
rect 353306 474038 353542 474274
rect 352986 454038 353222 454274
rect 353306 454038 353542 454274
rect 352986 434038 353222 434274
rect 353306 434038 353542 434274
rect 355546 707482 355782 707718
rect 355866 707482 356102 707718
rect 355546 707162 355782 707398
rect 355866 707162 356102 707398
rect 355546 696718 355782 696954
rect 355866 696718 356102 696954
rect 355546 676718 355782 676954
rect 355866 676718 356102 676954
rect 355546 656718 355782 656954
rect 355866 656718 356102 656954
rect 355546 636718 355782 636954
rect 355866 636718 356102 636954
rect 355546 616718 355782 616954
rect 355866 616718 356102 616954
rect 355546 596718 355782 596954
rect 355866 596718 356102 596954
rect 355546 576718 355782 576954
rect 355866 576718 356102 576954
rect 355546 556718 355782 556954
rect 355866 556718 356102 556954
rect 355546 536718 355782 536954
rect 355866 536718 356102 536954
rect 355546 516718 355782 516954
rect 355866 516718 356102 516954
rect 355546 496718 355782 496954
rect 355866 496718 356102 496954
rect 355546 476718 355782 476954
rect 355866 476718 356102 476954
rect 355546 456718 355782 456954
rect 355866 456718 356102 456954
rect 355546 436718 355782 436954
rect 355866 436718 356102 436954
rect 359266 700378 359502 700614
rect 359586 700378 359822 700614
rect 359266 680378 359502 680614
rect 359586 680378 359822 680614
rect 359266 660378 359502 660614
rect 359586 660378 359822 660614
rect 359266 640378 359502 640614
rect 359586 640378 359822 640614
rect 359266 620378 359502 620614
rect 359586 620378 359822 620614
rect 359266 600378 359502 600614
rect 359586 600378 359822 600614
rect 359266 580378 359502 580614
rect 359586 580378 359822 580614
rect 359266 560378 359502 560614
rect 359586 560378 359822 560614
rect 359266 540378 359502 540614
rect 359586 540378 359822 540614
rect 359266 520378 359502 520614
rect 359586 520378 359822 520614
rect 359266 500378 359502 500614
rect 359586 500378 359822 500614
rect 359266 480378 359502 480614
rect 359586 480378 359822 480614
rect 359266 460378 359502 460614
rect 359586 460378 359822 460614
rect 359266 440378 359502 440614
rect 359586 440378 359822 440614
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 683058 362062 683294
rect 362146 683058 362382 683294
rect 361826 663058 362062 663294
rect 362146 663058 362382 663294
rect 361826 643058 362062 643294
rect 362146 643058 362382 643294
rect 361826 623058 362062 623294
rect 362146 623058 362382 623294
rect 361826 603058 362062 603294
rect 362146 603058 362382 603294
rect 361826 583058 362062 583294
rect 362146 583058 362382 583294
rect 361826 563058 362062 563294
rect 362146 563058 362382 563294
rect 361826 543058 362062 543294
rect 362146 543058 362382 543294
rect 361826 523058 362062 523294
rect 362146 523058 362382 523294
rect 361826 503058 362062 503294
rect 362146 503058 362382 503294
rect 361826 483058 362062 483294
rect 362146 483058 362382 483294
rect 361826 463058 362062 463294
rect 362146 463058 362382 463294
rect 361826 443058 362062 443294
rect 362146 443058 362382 443294
rect 361826 423058 362062 423294
rect 362146 423058 362382 423294
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 362986 684038 363222 684274
rect 363306 684038 363542 684274
rect 362986 664038 363222 664274
rect 363306 664038 363542 664274
rect 362986 644038 363222 644274
rect 363306 644038 363542 644274
rect 362986 624038 363222 624274
rect 363306 624038 363542 624274
rect 362986 604038 363222 604274
rect 363306 604038 363542 604274
rect 362986 584038 363222 584274
rect 363306 584038 363542 584274
rect 362986 564038 363222 564274
rect 363306 564038 363542 564274
rect 362986 544038 363222 544274
rect 363306 544038 363542 544274
rect 362986 524038 363222 524274
rect 363306 524038 363542 524274
rect 362986 504038 363222 504274
rect 363306 504038 363542 504274
rect 362986 484038 363222 484274
rect 363306 484038 363542 484274
rect 362986 464038 363222 464274
rect 363306 464038 363542 464274
rect 362986 444038 363222 444274
rect 363306 444038 363542 444274
rect 362986 424038 363222 424274
rect 363306 424038 363542 424274
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 365546 686718 365782 686954
rect 365866 686718 366102 686954
rect 365546 666718 365782 666954
rect 365866 666718 366102 666954
rect 365546 646718 365782 646954
rect 365866 646718 366102 646954
rect 365546 626718 365782 626954
rect 365866 626718 366102 626954
rect 365546 606718 365782 606954
rect 365866 606718 366102 606954
rect 365546 586718 365782 586954
rect 365866 586718 366102 586954
rect 365546 566718 365782 566954
rect 365866 566718 366102 566954
rect 365546 546718 365782 546954
rect 365866 546718 366102 546954
rect 365546 526718 365782 526954
rect 365866 526718 366102 526954
rect 365546 506718 365782 506954
rect 365866 506718 366102 506954
rect 365546 486718 365782 486954
rect 365866 486718 366102 486954
rect 365546 466718 365782 466954
rect 365866 466718 366102 466954
rect 365546 446718 365782 446954
rect 365866 446718 366102 446954
rect 365546 426718 365782 426954
rect 365866 426718 366102 426954
rect 369266 690378 369502 690614
rect 369586 690378 369822 690614
rect 369266 670378 369502 670614
rect 369586 670378 369822 670614
rect 369266 650378 369502 650614
rect 369586 650378 369822 650614
rect 369266 630378 369502 630614
rect 369586 630378 369822 630614
rect 369266 610378 369502 610614
rect 369586 610378 369822 610614
rect 369266 590378 369502 590614
rect 369586 590378 369822 590614
rect 369266 570378 369502 570614
rect 369586 570378 369822 570614
rect 369266 550378 369502 550614
rect 369586 550378 369822 550614
rect 369266 530378 369502 530614
rect 369586 530378 369822 530614
rect 369266 510378 369502 510614
rect 369586 510378 369822 510614
rect 369266 490378 369502 490614
rect 369586 490378 369822 490614
rect 369266 470378 369502 470614
rect 369586 470378 369822 470614
rect 369266 450378 369502 450614
rect 369586 450378 369822 450614
rect 369266 430378 369502 430614
rect 369586 430378 369822 430614
rect 371826 705562 372062 705798
rect 372146 705562 372382 705798
rect 371826 705242 372062 705478
rect 372146 705242 372382 705478
rect 371826 693058 372062 693294
rect 372146 693058 372382 693294
rect 371826 673058 372062 673294
rect 372146 673058 372382 673294
rect 371826 653058 372062 653294
rect 372146 653058 372382 653294
rect 371826 633058 372062 633294
rect 372146 633058 372382 633294
rect 371826 613058 372062 613294
rect 372146 613058 372382 613294
rect 371826 593058 372062 593294
rect 372146 593058 372382 593294
rect 371826 573058 372062 573294
rect 372146 573058 372382 573294
rect 371826 553058 372062 553294
rect 372146 553058 372382 553294
rect 371826 533058 372062 533294
rect 372146 533058 372382 533294
rect 371826 513058 372062 513294
rect 372146 513058 372382 513294
rect 371826 493058 372062 493294
rect 372146 493058 372382 493294
rect 371826 473058 372062 473294
rect 372146 473058 372382 473294
rect 371826 453058 372062 453294
rect 372146 453058 372382 453294
rect 371826 433058 372062 433294
rect 372146 433058 372382 433294
rect 382986 711322 383222 711558
rect 383306 711322 383542 711558
rect 382986 711002 383222 711238
rect 383306 711002 383542 711238
rect 379266 709402 379502 709638
rect 379586 709402 379822 709638
rect 379266 709082 379502 709318
rect 379586 709082 379822 709318
rect 372986 694038 373222 694274
rect 373306 694038 373542 694274
rect 372986 674038 373222 674274
rect 373306 674038 373542 674274
rect 372986 654038 373222 654274
rect 373306 654038 373542 654274
rect 372986 634038 373222 634274
rect 373306 634038 373542 634274
rect 372986 614038 373222 614274
rect 373306 614038 373542 614274
rect 372986 594038 373222 594274
rect 373306 594038 373542 594274
rect 372986 574038 373222 574274
rect 373306 574038 373542 574274
rect 372986 554038 373222 554274
rect 373306 554038 373542 554274
rect 372986 534038 373222 534274
rect 373306 534038 373542 534274
rect 372986 514038 373222 514274
rect 373306 514038 373542 514274
rect 372986 494038 373222 494274
rect 373306 494038 373542 494274
rect 372986 474038 373222 474274
rect 373306 474038 373542 474274
rect 372986 454038 373222 454274
rect 373306 454038 373542 454274
rect 372986 434038 373222 434274
rect 373306 434038 373542 434274
rect 375546 707482 375782 707718
rect 375866 707482 376102 707718
rect 375546 707162 375782 707398
rect 375866 707162 376102 707398
rect 375546 696718 375782 696954
rect 375866 696718 376102 696954
rect 375546 676718 375782 676954
rect 375866 676718 376102 676954
rect 375546 656718 375782 656954
rect 375866 656718 376102 656954
rect 375546 636718 375782 636954
rect 375866 636718 376102 636954
rect 375546 616718 375782 616954
rect 375866 616718 376102 616954
rect 375546 596718 375782 596954
rect 375866 596718 376102 596954
rect 375546 576718 375782 576954
rect 375866 576718 376102 576954
rect 375546 556718 375782 556954
rect 375866 556718 376102 556954
rect 375546 536718 375782 536954
rect 375866 536718 376102 536954
rect 375546 516718 375782 516954
rect 375866 516718 376102 516954
rect 375546 496718 375782 496954
rect 375866 496718 376102 496954
rect 375546 476718 375782 476954
rect 375866 476718 376102 476954
rect 375546 456718 375782 456954
rect 375866 456718 376102 456954
rect 375546 436718 375782 436954
rect 375866 436718 376102 436954
rect 379266 700378 379502 700614
rect 379586 700378 379822 700614
rect 379266 680378 379502 680614
rect 379586 680378 379822 680614
rect 379266 660378 379502 660614
rect 379586 660378 379822 660614
rect 379266 640378 379502 640614
rect 379586 640378 379822 640614
rect 379266 620378 379502 620614
rect 379586 620378 379822 620614
rect 379266 600378 379502 600614
rect 379586 600378 379822 600614
rect 379266 580378 379502 580614
rect 379586 580378 379822 580614
rect 379266 560378 379502 560614
rect 379586 560378 379822 560614
rect 379266 540378 379502 540614
rect 379586 540378 379822 540614
rect 379266 520378 379502 520614
rect 379586 520378 379822 520614
rect 379266 500378 379502 500614
rect 379586 500378 379822 500614
rect 379266 480378 379502 480614
rect 379586 480378 379822 480614
rect 379266 460378 379502 460614
rect 379586 460378 379822 460614
rect 379266 440378 379502 440614
rect 379586 440378 379822 440614
rect 381826 704602 382062 704838
rect 382146 704602 382382 704838
rect 381826 704282 382062 704518
rect 382146 704282 382382 704518
rect 381826 683058 382062 683294
rect 382146 683058 382382 683294
rect 381826 663058 382062 663294
rect 382146 663058 382382 663294
rect 381826 643058 382062 643294
rect 382146 643058 382382 643294
rect 381826 623058 382062 623294
rect 382146 623058 382382 623294
rect 381826 603058 382062 603294
rect 382146 603058 382382 603294
rect 381826 583058 382062 583294
rect 382146 583058 382382 583294
rect 381826 563058 382062 563294
rect 382146 563058 382382 563294
rect 381826 543058 382062 543294
rect 382146 543058 382382 543294
rect 381826 523058 382062 523294
rect 382146 523058 382382 523294
rect 381826 503058 382062 503294
rect 382146 503058 382382 503294
rect 381826 483058 382062 483294
rect 382146 483058 382382 483294
rect 381826 463058 382062 463294
rect 382146 463058 382382 463294
rect 381826 443058 382062 443294
rect 382146 443058 382382 443294
rect 381826 423058 382062 423294
rect 382146 423058 382382 423294
rect 392986 710362 393222 710598
rect 393306 710362 393542 710598
rect 392986 710042 393222 710278
rect 393306 710042 393542 710278
rect 389266 708442 389502 708678
rect 389586 708442 389822 708678
rect 389266 708122 389502 708358
rect 389586 708122 389822 708358
rect 382986 684038 383222 684274
rect 383306 684038 383542 684274
rect 382986 664038 383222 664274
rect 383306 664038 383542 664274
rect 382986 644038 383222 644274
rect 383306 644038 383542 644274
rect 382986 624038 383222 624274
rect 383306 624038 383542 624274
rect 382986 604038 383222 604274
rect 383306 604038 383542 604274
rect 382986 584038 383222 584274
rect 383306 584038 383542 584274
rect 382986 564038 383222 564274
rect 383306 564038 383542 564274
rect 382986 544038 383222 544274
rect 383306 544038 383542 544274
rect 382986 524038 383222 524274
rect 383306 524038 383542 524274
rect 382986 504038 383222 504274
rect 383306 504038 383542 504274
rect 382986 484038 383222 484274
rect 383306 484038 383542 484274
rect 382986 464038 383222 464274
rect 383306 464038 383542 464274
rect 382986 444038 383222 444274
rect 383306 444038 383542 444274
rect 382986 424038 383222 424274
rect 383306 424038 383542 424274
rect 385546 706522 385782 706758
rect 385866 706522 386102 706758
rect 385546 706202 385782 706438
rect 385866 706202 386102 706438
rect 385546 686718 385782 686954
rect 385866 686718 386102 686954
rect 385546 666718 385782 666954
rect 385866 666718 386102 666954
rect 385546 646718 385782 646954
rect 385866 646718 386102 646954
rect 385546 626718 385782 626954
rect 385866 626718 386102 626954
rect 385546 606718 385782 606954
rect 385866 606718 386102 606954
rect 385546 586718 385782 586954
rect 385866 586718 386102 586954
rect 385546 566718 385782 566954
rect 385866 566718 386102 566954
rect 385546 546718 385782 546954
rect 385866 546718 386102 546954
rect 385546 526718 385782 526954
rect 385866 526718 386102 526954
rect 385546 506718 385782 506954
rect 385866 506718 386102 506954
rect 385546 486718 385782 486954
rect 385866 486718 386102 486954
rect 385546 466718 385782 466954
rect 385866 466718 386102 466954
rect 385546 446718 385782 446954
rect 385866 446718 386102 446954
rect 385546 426718 385782 426954
rect 385866 426718 386102 426954
rect 389266 690378 389502 690614
rect 389586 690378 389822 690614
rect 389266 670378 389502 670614
rect 389586 670378 389822 670614
rect 389266 650378 389502 650614
rect 389586 650378 389822 650614
rect 389266 630378 389502 630614
rect 389586 630378 389822 630614
rect 389266 610378 389502 610614
rect 389586 610378 389822 610614
rect 389266 590378 389502 590614
rect 389586 590378 389822 590614
rect 389266 570378 389502 570614
rect 389586 570378 389822 570614
rect 389266 550378 389502 550614
rect 389586 550378 389822 550614
rect 389266 530378 389502 530614
rect 389586 530378 389822 530614
rect 389266 510378 389502 510614
rect 389586 510378 389822 510614
rect 389266 490378 389502 490614
rect 389586 490378 389822 490614
rect 389266 470378 389502 470614
rect 389586 470378 389822 470614
rect 389266 450378 389502 450614
rect 389586 450378 389822 450614
rect 389266 430378 389502 430614
rect 389586 430378 389822 430614
rect 391826 705562 392062 705798
rect 392146 705562 392382 705798
rect 391826 705242 392062 705478
rect 392146 705242 392382 705478
rect 391826 693058 392062 693294
rect 392146 693058 392382 693294
rect 391826 673058 392062 673294
rect 392146 673058 392382 673294
rect 391826 653058 392062 653294
rect 392146 653058 392382 653294
rect 391826 633058 392062 633294
rect 392146 633058 392382 633294
rect 391826 613058 392062 613294
rect 392146 613058 392382 613294
rect 391826 593058 392062 593294
rect 392146 593058 392382 593294
rect 391826 573058 392062 573294
rect 392146 573058 392382 573294
rect 391826 553058 392062 553294
rect 392146 553058 392382 553294
rect 391826 533058 392062 533294
rect 392146 533058 392382 533294
rect 391826 513058 392062 513294
rect 392146 513058 392382 513294
rect 391826 493058 392062 493294
rect 392146 493058 392382 493294
rect 391826 473058 392062 473294
rect 392146 473058 392382 473294
rect 391826 453058 392062 453294
rect 392146 453058 392382 453294
rect 391826 433058 392062 433294
rect 392146 433058 392382 433294
rect 402986 711322 403222 711558
rect 403306 711322 403542 711558
rect 402986 711002 403222 711238
rect 403306 711002 403542 711238
rect 399266 709402 399502 709638
rect 399586 709402 399822 709638
rect 399266 709082 399502 709318
rect 399586 709082 399822 709318
rect 392986 694038 393222 694274
rect 393306 694038 393542 694274
rect 392986 674038 393222 674274
rect 393306 674038 393542 674274
rect 392986 654038 393222 654274
rect 393306 654038 393542 654274
rect 392986 634038 393222 634274
rect 393306 634038 393542 634274
rect 392986 614038 393222 614274
rect 393306 614038 393542 614274
rect 392986 594038 393222 594274
rect 393306 594038 393542 594274
rect 392986 574038 393222 574274
rect 393306 574038 393542 574274
rect 392986 554038 393222 554274
rect 393306 554038 393542 554274
rect 392986 534038 393222 534274
rect 393306 534038 393542 534274
rect 392986 514038 393222 514274
rect 393306 514038 393542 514274
rect 392986 494038 393222 494274
rect 393306 494038 393542 494274
rect 392986 474038 393222 474274
rect 393306 474038 393542 474274
rect 392986 454038 393222 454274
rect 393306 454038 393542 454274
rect 392986 434038 393222 434274
rect 393306 434038 393542 434274
rect 395546 707482 395782 707718
rect 395866 707482 396102 707718
rect 395546 707162 395782 707398
rect 395866 707162 396102 707398
rect 395546 696718 395782 696954
rect 395866 696718 396102 696954
rect 395546 676718 395782 676954
rect 395866 676718 396102 676954
rect 395546 656718 395782 656954
rect 395866 656718 396102 656954
rect 395546 636718 395782 636954
rect 395866 636718 396102 636954
rect 395546 616718 395782 616954
rect 395866 616718 396102 616954
rect 395546 596718 395782 596954
rect 395866 596718 396102 596954
rect 395546 576718 395782 576954
rect 395866 576718 396102 576954
rect 395546 556718 395782 556954
rect 395866 556718 396102 556954
rect 395546 536718 395782 536954
rect 395866 536718 396102 536954
rect 395546 516718 395782 516954
rect 395866 516718 396102 516954
rect 395546 496718 395782 496954
rect 395866 496718 396102 496954
rect 395546 476718 395782 476954
rect 395866 476718 396102 476954
rect 395546 456718 395782 456954
rect 395866 456718 396102 456954
rect 395546 436718 395782 436954
rect 395866 436718 396102 436954
rect 399266 700378 399502 700614
rect 399586 700378 399822 700614
rect 399266 680378 399502 680614
rect 399586 680378 399822 680614
rect 399266 660378 399502 660614
rect 399586 660378 399822 660614
rect 399266 640378 399502 640614
rect 399586 640378 399822 640614
rect 399266 620378 399502 620614
rect 399586 620378 399822 620614
rect 399266 600378 399502 600614
rect 399586 600378 399822 600614
rect 399266 580378 399502 580614
rect 399586 580378 399822 580614
rect 399266 560378 399502 560614
rect 399586 560378 399822 560614
rect 399266 540378 399502 540614
rect 399586 540378 399822 540614
rect 399266 520378 399502 520614
rect 399586 520378 399822 520614
rect 399266 500378 399502 500614
rect 399586 500378 399822 500614
rect 399266 480378 399502 480614
rect 399586 480378 399822 480614
rect 399266 460378 399502 460614
rect 399586 460378 399822 460614
rect 399266 440378 399502 440614
rect 399586 440378 399822 440614
rect 401826 704602 402062 704838
rect 402146 704602 402382 704838
rect 401826 704282 402062 704518
rect 402146 704282 402382 704518
rect 401826 683058 402062 683294
rect 402146 683058 402382 683294
rect 401826 663058 402062 663294
rect 402146 663058 402382 663294
rect 401826 643058 402062 643294
rect 402146 643058 402382 643294
rect 401826 623058 402062 623294
rect 402146 623058 402382 623294
rect 401826 603058 402062 603294
rect 402146 603058 402382 603294
rect 401826 583058 402062 583294
rect 402146 583058 402382 583294
rect 401826 563058 402062 563294
rect 402146 563058 402382 563294
rect 401826 543058 402062 543294
rect 402146 543058 402382 543294
rect 401826 523058 402062 523294
rect 402146 523058 402382 523294
rect 401826 503058 402062 503294
rect 402146 503058 402382 503294
rect 401826 483058 402062 483294
rect 402146 483058 402382 483294
rect 401826 463058 402062 463294
rect 402146 463058 402382 463294
rect 401826 443058 402062 443294
rect 402146 443058 402382 443294
rect 401826 423058 402062 423294
rect 402146 423058 402382 423294
rect 412986 710362 413222 710598
rect 413306 710362 413542 710598
rect 412986 710042 413222 710278
rect 413306 710042 413542 710278
rect 409266 708442 409502 708678
rect 409586 708442 409822 708678
rect 409266 708122 409502 708358
rect 409586 708122 409822 708358
rect 402986 684038 403222 684274
rect 403306 684038 403542 684274
rect 402986 664038 403222 664274
rect 403306 664038 403542 664274
rect 402986 644038 403222 644274
rect 403306 644038 403542 644274
rect 402986 624038 403222 624274
rect 403306 624038 403542 624274
rect 402986 604038 403222 604274
rect 403306 604038 403542 604274
rect 402986 584038 403222 584274
rect 403306 584038 403542 584274
rect 402986 564038 403222 564274
rect 403306 564038 403542 564274
rect 402986 544038 403222 544274
rect 403306 544038 403542 544274
rect 402986 524038 403222 524274
rect 403306 524038 403542 524274
rect 402986 504038 403222 504274
rect 403306 504038 403542 504274
rect 402986 484038 403222 484274
rect 403306 484038 403542 484274
rect 402986 464038 403222 464274
rect 403306 464038 403542 464274
rect 402986 444038 403222 444274
rect 403306 444038 403542 444274
rect 402986 424038 403222 424274
rect 403306 424038 403542 424274
rect 405546 706522 405782 706758
rect 405866 706522 406102 706758
rect 405546 706202 405782 706438
rect 405866 706202 406102 706438
rect 405546 686718 405782 686954
rect 405866 686718 406102 686954
rect 405546 666718 405782 666954
rect 405866 666718 406102 666954
rect 409266 690378 409502 690614
rect 409586 690378 409822 690614
rect 409266 670378 409502 670614
rect 409586 670378 409822 670614
rect 411826 705562 412062 705798
rect 412146 705562 412382 705798
rect 411826 705242 412062 705478
rect 412146 705242 412382 705478
rect 411826 693058 412062 693294
rect 412146 693058 412382 693294
rect 411826 673058 412062 673294
rect 412146 673058 412382 673294
rect 422986 711322 423222 711558
rect 423306 711322 423542 711558
rect 422986 711002 423222 711238
rect 423306 711002 423542 711238
rect 419266 709402 419502 709638
rect 419586 709402 419822 709638
rect 419266 709082 419502 709318
rect 419586 709082 419822 709318
rect 412986 694038 413222 694274
rect 413306 694038 413542 694274
rect 412986 674038 413222 674274
rect 413306 674038 413542 674274
rect 415546 707482 415782 707718
rect 415866 707482 416102 707718
rect 415546 707162 415782 707398
rect 415866 707162 416102 707398
rect 415546 696718 415782 696954
rect 415866 696718 416102 696954
rect 415546 676718 415782 676954
rect 415866 676718 416102 676954
rect 419266 700378 419502 700614
rect 419586 700378 419822 700614
rect 419266 680378 419502 680614
rect 419586 680378 419822 680614
rect 419266 660378 419502 660614
rect 419586 660378 419822 660614
rect 421826 704602 422062 704838
rect 422146 704602 422382 704838
rect 421826 704282 422062 704518
rect 422146 704282 422382 704518
rect 421826 683058 422062 683294
rect 422146 683058 422382 683294
rect 421826 663058 422062 663294
rect 422146 663058 422382 663294
rect 432986 710362 433222 710598
rect 433306 710362 433542 710598
rect 432986 710042 433222 710278
rect 433306 710042 433542 710278
rect 429266 708442 429502 708678
rect 429586 708442 429822 708678
rect 429266 708122 429502 708358
rect 429586 708122 429822 708358
rect 422986 684038 423222 684274
rect 423306 684038 423542 684274
rect 422986 664038 423222 664274
rect 423306 664038 423542 664274
rect 425546 706522 425782 706758
rect 425866 706522 426102 706758
rect 425546 706202 425782 706438
rect 425866 706202 426102 706438
rect 425546 686718 425782 686954
rect 425866 686718 426102 686954
rect 425546 666718 425782 666954
rect 425866 666718 426102 666954
rect 429266 690378 429502 690614
rect 429586 690378 429822 690614
rect 429266 670378 429502 670614
rect 429586 670378 429822 670614
rect 431826 705562 432062 705798
rect 432146 705562 432382 705798
rect 431826 705242 432062 705478
rect 432146 705242 432382 705478
rect 431826 693058 432062 693294
rect 432146 693058 432382 693294
rect 431826 673058 432062 673294
rect 432146 673058 432382 673294
rect 442986 711322 443222 711558
rect 443306 711322 443542 711558
rect 442986 711002 443222 711238
rect 443306 711002 443542 711238
rect 439266 709402 439502 709638
rect 439586 709402 439822 709638
rect 439266 709082 439502 709318
rect 439586 709082 439822 709318
rect 432986 694038 433222 694274
rect 433306 694038 433542 694274
rect 432986 674038 433222 674274
rect 433306 674038 433542 674274
rect 435546 707482 435782 707718
rect 435866 707482 436102 707718
rect 435546 707162 435782 707398
rect 435866 707162 436102 707398
rect 435546 696718 435782 696954
rect 435866 696718 436102 696954
rect 435546 676718 435782 676954
rect 435866 676718 436102 676954
rect 439266 700378 439502 700614
rect 439586 700378 439822 700614
rect 439266 680378 439502 680614
rect 439586 680378 439822 680614
rect 439266 660378 439502 660614
rect 439586 660378 439822 660614
rect 441826 704602 442062 704838
rect 442146 704602 442382 704838
rect 441826 704282 442062 704518
rect 442146 704282 442382 704518
rect 441826 683058 442062 683294
rect 442146 683058 442382 683294
rect 441826 663058 442062 663294
rect 442146 663058 442382 663294
rect 452986 710362 453222 710598
rect 453306 710362 453542 710598
rect 452986 710042 453222 710278
rect 453306 710042 453542 710278
rect 449266 708442 449502 708678
rect 449586 708442 449822 708678
rect 449266 708122 449502 708358
rect 449586 708122 449822 708358
rect 442986 684038 443222 684274
rect 443306 684038 443542 684274
rect 442986 664038 443222 664274
rect 443306 664038 443542 664274
rect 445546 706522 445782 706758
rect 445866 706522 446102 706758
rect 445546 706202 445782 706438
rect 445866 706202 446102 706438
rect 445546 686718 445782 686954
rect 445866 686718 446102 686954
rect 445546 666718 445782 666954
rect 445866 666718 446102 666954
rect 449266 690378 449502 690614
rect 449586 690378 449822 690614
rect 449266 670378 449502 670614
rect 449586 670378 449822 670614
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 693058 452062 693294
rect 452146 693058 452382 693294
rect 451826 673058 452062 673294
rect 452146 673058 452382 673294
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 452986 694038 453222 694274
rect 453306 694038 453542 694274
rect 452986 674038 453222 674274
rect 453306 674038 453542 674274
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 455546 696718 455782 696954
rect 455866 696718 456102 696954
rect 455546 676718 455782 676954
rect 455866 676718 456102 676954
rect 459266 700378 459502 700614
rect 459586 700378 459822 700614
rect 459266 680378 459502 680614
rect 459586 680378 459822 680614
rect 459266 660378 459502 660614
rect 459586 660378 459822 660614
rect 461826 704602 462062 704838
rect 462146 704602 462382 704838
rect 461826 704282 462062 704518
rect 462146 704282 462382 704518
rect 461826 683058 462062 683294
rect 462146 683058 462382 683294
rect 461826 663058 462062 663294
rect 462146 663058 462382 663294
rect 472986 710362 473222 710598
rect 473306 710362 473542 710598
rect 472986 710042 473222 710278
rect 473306 710042 473542 710278
rect 469266 708442 469502 708678
rect 469586 708442 469822 708678
rect 469266 708122 469502 708358
rect 469586 708122 469822 708358
rect 462986 684038 463222 684274
rect 463306 684038 463542 684274
rect 462986 664038 463222 664274
rect 463306 664038 463542 664274
rect 465546 706522 465782 706758
rect 465866 706522 466102 706758
rect 465546 706202 465782 706438
rect 465866 706202 466102 706438
rect 465546 686718 465782 686954
rect 465866 686718 466102 686954
rect 465546 666718 465782 666954
rect 465866 666718 466102 666954
rect 469266 690378 469502 690614
rect 469586 690378 469822 690614
rect 469266 670378 469502 670614
rect 469586 670378 469822 670614
rect 471826 705562 472062 705798
rect 472146 705562 472382 705798
rect 471826 705242 472062 705478
rect 472146 705242 472382 705478
rect 471826 693058 472062 693294
rect 472146 693058 472382 693294
rect 471826 673058 472062 673294
rect 472146 673058 472382 673294
rect 482986 711322 483222 711558
rect 483306 711322 483542 711558
rect 482986 711002 483222 711238
rect 483306 711002 483542 711238
rect 479266 709402 479502 709638
rect 479586 709402 479822 709638
rect 479266 709082 479502 709318
rect 479586 709082 479822 709318
rect 472986 694038 473222 694274
rect 473306 694038 473542 694274
rect 472986 674038 473222 674274
rect 473306 674038 473542 674274
rect 475546 707482 475782 707718
rect 475866 707482 476102 707718
rect 475546 707162 475782 707398
rect 475866 707162 476102 707398
rect 475546 696718 475782 696954
rect 475866 696718 476102 696954
rect 475546 676718 475782 676954
rect 475866 676718 476102 676954
rect 479266 700378 479502 700614
rect 479586 700378 479822 700614
rect 479266 680378 479502 680614
rect 479586 680378 479822 680614
rect 479266 660378 479502 660614
rect 479586 660378 479822 660614
rect 481826 704602 482062 704838
rect 482146 704602 482382 704838
rect 481826 704282 482062 704518
rect 482146 704282 482382 704518
rect 481826 683058 482062 683294
rect 482146 683058 482382 683294
rect 481826 663058 482062 663294
rect 482146 663058 482382 663294
rect 492986 710362 493222 710598
rect 493306 710362 493542 710598
rect 492986 710042 493222 710278
rect 493306 710042 493542 710278
rect 489266 708442 489502 708678
rect 489586 708442 489822 708678
rect 489266 708122 489502 708358
rect 489586 708122 489822 708358
rect 482986 684038 483222 684274
rect 483306 684038 483542 684274
rect 482986 664038 483222 664274
rect 483306 664038 483542 664274
rect 485546 706522 485782 706758
rect 485866 706522 486102 706758
rect 485546 706202 485782 706438
rect 485866 706202 486102 706438
rect 485546 686718 485782 686954
rect 485866 686718 486102 686954
rect 485546 666718 485782 666954
rect 485866 666718 486102 666954
rect 489266 690378 489502 690614
rect 489586 690378 489822 690614
rect 489266 670378 489502 670614
rect 489586 670378 489822 670614
rect 491826 705562 492062 705798
rect 492146 705562 492382 705798
rect 491826 705242 492062 705478
rect 492146 705242 492382 705478
rect 491826 693058 492062 693294
rect 492146 693058 492382 693294
rect 491826 673058 492062 673294
rect 492146 673058 492382 673294
rect 502986 711322 503222 711558
rect 503306 711322 503542 711558
rect 502986 711002 503222 711238
rect 503306 711002 503542 711238
rect 499266 709402 499502 709638
rect 499586 709402 499822 709638
rect 499266 709082 499502 709318
rect 499586 709082 499822 709318
rect 492986 694038 493222 694274
rect 493306 694038 493542 694274
rect 492986 674038 493222 674274
rect 493306 674038 493542 674274
rect 495546 707482 495782 707718
rect 495866 707482 496102 707718
rect 495546 707162 495782 707398
rect 495866 707162 496102 707398
rect 495546 696718 495782 696954
rect 495866 696718 496102 696954
rect 495546 676718 495782 676954
rect 495866 676718 496102 676954
rect 499266 700378 499502 700614
rect 499586 700378 499822 700614
rect 499266 680378 499502 680614
rect 499586 680378 499822 680614
rect 499266 660378 499502 660614
rect 499586 660378 499822 660614
rect 501826 704602 502062 704838
rect 502146 704602 502382 704838
rect 501826 704282 502062 704518
rect 502146 704282 502382 704518
rect 501826 683058 502062 683294
rect 502146 683058 502382 683294
rect 501826 663058 502062 663294
rect 502146 663058 502382 663294
rect 512986 710362 513222 710598
rect 513306 710362 513542 710598
rect 512986 710042 513222 710278
rect 513306 710042 513542 710278
rect 509266 708442 509502 708678
rect 509586 708442 509822 708678
rect 509266 708122 509502 708358
rect 509586 708122 509822 708358
rect 502986 684038 503222 684274
rect 503306 684038 503542 684274
rect 502986 664038 503222 664274
rect 503306 664038 503542 664274
rect 505546 706522 505782 706758
rect 505866 706522 506102 706758
rect 505546 706202 505782 706438
rect 505866 706202 506102 706438
rect 505546 686718 505782 686954
rect 505866 686718 506102 686954
rect 505546 666718 505782 666954
rect 505866 666718 506102 666954
rect 509266 690378 509502 690614
rect 509586 690378 509822 690614
rect 509266 670378 509502 670614
rect 509586 670378 509822 670614
rect 410328 653058 410564 653294
rect 505392 653058 505628 653294
rect 405546 646718 405782 646954
rect 405866 646718 406102 646954
rect 509266 650378 509502 650614
rect 509586 650378 509822 650614
rect 411008 643058 411244 643294
rect 504712 643058 504948 643294
rect 410328 633058 410564 633294
rect 505392 633058 505628 633294
rect 405546 626718 405782 626954
rect 405866 626718 406102 626954
rect 509266 630378 509502 630614
rect 509586 630378 509822 630614
rect 411008 623058 411244 623294
rect 504712 623058 504948 623294
rect 410328 613058 410564 613294
rect 505392 613058 505628 613294
rect 405546 606718 405782 606954
rect 405866 606718 406102 606954
rect 509266 610378 509502 610614
rect 509586 610378 509822 610614
rect 411008 603058 411244 603294
rect 504712 603058 504948 603294
rect 410328 593058 410564 593294
rect 505392 593058 505628 593294
rect 405546 586718 405782 586954
rect 405866 586718 406102 586954
rect 509266 590378 509502 590614
rect 509586 590378 509822 590614
rect 411008 583058 411244 583294
rect 504712 583058 504948 583294
rect 405546 566718 405782 566954
rect 405866 566718 406102 566954
rect 405546 546718 405782 546954
rect 405866 546718 406102 546954
rect 409266 570378 409502 570614
rect 409586 570378 409822 570614
rect 409266 550378 409502 550614
rect 409586 550378 409822 550614
rect 411826 573058 412062 573294
rect 412146 573058 412382 573294
rect 411826 553058 412062 553294
rect 412146 553058 412382 553294
rect 412986 574038 413222 574274
rect 413306 574038 413542 574274
rect 412986 554038 413222 554274
rect 413306 554038 413542 554274
rect 415546 556718 415782 556954
rect 415866 556718 416102 556954
rect 419266 560378 419502 560614
rect 419586 560378 419822 560614
rect 419266 540378 419502 540614
rect 419586 540378 419822 540614
rect 421826 563058 422062 563294
rect 422146 563058 422382 563294
rect 421826 543058 422062 543294
rect 422146 543058 422382 543294
rect 422986 564038 423222 564274
rect 423306 564038 423542 564274
rect 422986 544038 423222 544274
rect 423306 544038 423542 544274
rect 425546 566718 425782 566954
rect 425866 566718 426102 566954
rect 425546 546718 425782 546954
rect 425866 546718 426102 546954
rect 429266 570378 429502 570614
rect 429586 570378 429822 570614
rect 429266 550378 429502 550614
rect 429586 550378 429822 550614
rect 431826 573058 432062 573294
rect 432146 573058 432382 573294
rect 431826 553058 432062 553294
rect 432146 553058 432382 553294
rect 432986 574038 433222 574274
rect 433306 574038 433542 574274
rect 432986 554038 433222 554274
rect 433306 554038 433542 554274
rect 435546 556718 435782 556954
rect 435866 556718 436102 556954
rect 439266 560378 439502 560614
rect 439586 560378 439822 560614
rect 439266 540378 439502 540614
rect 439586 540378 439822 540614
rect 441826 563058 442062 563294
rect 442146 563058 442382 563294
rect 441826 543058 442062 543294
rect 442146 543058 442382 543294
rect 442986 564038 443222 564274
rect 443306 564038 443542 564274
rect 442986 544038 443222 544274
rect 443306 544038 443542 544274
rect 445546 566718 445782 566954
rect 445866 566718 446102 566954
rect 445546 546718 445782 546954
rect 445866 546718 446102 546954
rect 449266 570378 449502 570614
rect 449586 570378 449822 570614
rect 449266 550378 449502 550614
rect 449586 550378 449822 550614
rect 451826 573058 452062 573294
rect 452146 573058 452382 573294
rect 451826 553058 452062 553294
rect 452146 553058 452382 553294
rect 452986 574038 453222 574274
rect 453306 574038 453542 574274
rect 452986 554038 453222 554274
rect 453306 554038 453542 554274
rect 455546 556718 455782 556954
rect 455866 556718 456102 556954
rect 459266 560378 459502 560614
rect 459586 560378 459822 560614
rect 459266 540378 459502 540614
rect 459586 540378 459822 540614
rect 461826 563058 462062 563294
rect 462146 563058 462382 563294
rect 461826 543058 462062 543294
rect 462146 543058 462382 543294
rect 462986 564038 463222 564274
rect 463306 564038 463542 564274
rect 462986 544038 463222 544274
rect 463306 544038 463542 544274
rect 465546 566718 465782 566954
rect 465866 566718 466102 566954
rect 465546 546718 465782 546954
rect 465866 546718 466102 546954
rect 469266 570378 469502 570614
rect 469586 570378 469822 570614
rect 469266 550378 469502 550614
rect 469586 550378 469822 550614
rect 471826 573058 472062 573294
rect 472146 573058 472382 573294
rect 471826 553058 472062 553294
rect 472146 553058 472382 553294
rect 472986 574038 473222 574274
rect 473306 574038 473542 574274
rect 472986 554038 473222 554274
rect 473306 554038 473542 554274
rect 475546 556718 475782 556954
rect 475866 556718 476102 556954
rect 479266 560378 479502 560614
rect 479586 560378 479822 560614
rect 479266 540378 479502 540614
rect 479586 540378 479822 540614
rect 481826 563058 482062 563294
rect 482146 563058 482382 563294
rect 481826 543058 482062 543294
rect 482146 543058 482382 543294
rect 482986 564038 483222 564274
rect 483306 564038 483542 564274
rect 482986 544038 483222 544274
rect 483306 544038 483542 544274
rect 485546 566718 485782 566954
rect 485866 566718 486102 566954
rect 485546 546718 485782 546954
rect 485866 546718 486102 546954
rect 489266 570378 489502 570614
rect 489586 570378 489822 570614
rect 489266 550378 489502 550614
rect 489586 550378 489822 550614
rect 491826 573058 492062 573294
rect 492146 573058 492382 573294
rect 491826 553058 492062 553294
rect 492146 553058 492382 553294
rect 492986 574038 493222 574274
rect 493306 574038 493542 574274
rect 492986 554038 493222 554274
rect 493306 554038 493542 554274
rect 495546 556718 495782 556954
rect 495866 556718 496102 556954
rect 499266 560378 499502 560614
rect 499586 560378 499822 560614
rect 499266 540378 499502 540614
rect 499586 540378 499822 540614
rect 501826 563058 502062 563294
rect 502146 563058 502382 563294
rect 501826 543058 502062 543294
rect 502146 543058 502382 543294
rect 502986 564038 503222 564274
rect 503306 564038 503542 564274
rect 502986 544038 503222 544274
rect 503306 544038 503542 544274
rect 505546 566718 505782 566954
rect 505866 566718 506102 566954
rect 505546 546718 505782 546954
rect 505866 546718 506102 546954
rect 509266 570378 509502 570614
rect 509586 570378 509822 570614
rect 509266 550378 509502 550614
rect 509586 550378 509822 550614
rect 511826 705562 512062 705798
rect 512146 705562 512382 705798
rect 511826 705242 512062 705478
rect 512146 705242 512382 705478
rect 511826 693058 512062 693294
rect 512146 693058 512382 693294
rect 511826 673058 512062 673294
rect 512146 673058 512382 673294
rect 511826 653058 512062 653294
rect 512146 653058 512382 653294
rect 511826 633058 512062 633294
rect 512146 633058 512382 633294
rect 511826 613058 512062 613294
rect 512146 613058 512382 613294
rect 511826 593058 512062 593294
rect 512146 593058 512382 593294
rect 511826 573058 512062 573294
rect 512146 573058 512382 573294
rect 511826 553058 512062 553294
rect 512146 553058 512382 553294
rect 522986 711322 523222 711558
rect 523306 711322 523542 711558
rect 522986 711002 523222 711238
rect 523306 711002 523542 711238
rect 519266 709402 519502 709638
rect 519586 709402 519822 709638
rect 519266 709082 519502 709318
rect 519586 709082 519822 709318
rect 512986 694038 513222 694274
rect 513306 694038 513542 694274
rect 512986 674038 513222 674274
rect 513306 674038 513542 674274
rect 512986 654038 513222 654274
rect 513306 654038 513542 654274
rect 512986 634038 513222 634274
rect 513306 634038 513542 634274
rect 512986 614038 513222 614274
rect 513306 614038 513542 614274
rect 512986 594038 513222 594274
rect 513306 594038 513542 594274
rect 512986 574038 513222 574274
rect 513306 574038 513542 574274
rect 512986 554038 513222 554274
rect 513306 554038 513542 554274
rect 515546 707482 515782 707718
rect 515866 707482 516102 707718
rect 515546 707162 515782 707398
rect 515866 707162 516102 707398
rect 515546 696718 515782 696954
rect 515866 696718 516102 696954
rect 515546 676718 515782 676954
rect 515866 676718 516102 676954
rect 515546 656718 515782 656954
rect 515866 656718 516102 656954
rect 515546 636718 515782 636954
rect 515866 636718 516102 636954
rect 515546 616718 515782 616954
rect 515866 616718 516102 616954
rect 515546 596718 515782 596954
rect 515866 596718 516102 596954
rect 515546 576718 515782 576954
rect 515866 576718 516102 576954
rect 515546 556718 515782 556954
rect 515866 556718 516102 556954
rect 519266 700378 519502 700614
rect 519586 700378 519822 700614
rect 519266 680378 519502 680614
rect 519586 680378 519822 680614
rect 519266 660378 519502 660614
rect 519586 660378 519822 660614
rect 519266 640378 519502 640614
rect 519586 640378 519822 640614
rect 519266 620378 519502 620614
rect 519586 620378 519822 620614
rect 519266 600378 519502 600614
rect 519586 600378 519822 600614
rect 519266 580378 519502 580614
rect 519586 580378 519822 580614
rect 519266 560378 519502 560614
rect 519586 560378 519822 560614
rect 519266 540378 519502 540614
rect 519586 540378 519822 540614
rect 521826 704602 522062 704838
rect 522146 704602 522382 704838
rect 521826 704282 522062 704518
rect 522146 704282 522382 704518
rect 521826 683058 522062 683294
rect 522146 683058 522382 683294
rect 521826 663058 522062 663294
rect 522146 663058 522382 663294
rect 521826 643058 522062 643294
rect 522146 643058 522382 643294
rect 521826 623058 522062 623294
rect 522146 623058 522382 623294
rect 521826 603058 522062 603294
rect 522146 603058 522382 603294
rect 521826 583058 522062 583294
rect 522146 583058 522382 583294
rect 521826 563058 522062 563294
rect 522146 563058 522382 563294
rect 521826 543058 522062 543294
rect 522146 543058 522382 543294
rect 532986 710362 533222 710598
rect 533306 710362 533542 710598
rect 532986 710042 533222 710278
rect 533306 710042 533542 710278
rect 529266 708442 529502 708678
rect 529586 708442 529822 708678
rect 529266 708122 529502 708358
rect 529586 708122 529822 708358
rect 522986 684038 523222 684274
rect 523306 684038 523542 684274
rect 522986 664038 523222 664274
rect 523306 664038 523542 664274
rect 522986 644038 523222 644274
rect 523306 644038 523542 644274
rect 522986 624038 523222 624274
rect 523306 624038 523542 624274
rect 522986 604038 523222 604274
rect 523306 604038 523542 604274
rect 522986 584038 523222 584274
rect 523306 584038 523542 584274
rect 522986 564038 523222 564274
rect 523306 564038 523542 564274
rect 522986 544038 523222 544274
rect 523306 544038 523542 544274
rect 525546 706522 525782 706758
rect 525866 706522 526102 706758
rect 525546 706202 525782 706438
rect 525866 706202 526102 706438
rect 525546 686718 525782 686954
rect 525866 686718 526102 686954
rect 525546 666718 525782 666954
rect 525866 666718 526102 666954
rect 525546 646718 525782 646954
rect 525866 646718 526102 646954
rect 525546 626718 525782 626954
rect 525866 626718 526102 626954
rect 525546 606718 525782 606954
rect 525866 606718 526102 606954
rect 525546 586718 525782 586954
rect 525866 586718 526102 586954
rect 525546 566718 525782 566954
rect 525866 566718 526102 566954
rect 525546 546718 525782 546954
rect 525866 546718 526102 546954
rect 529266 690378 529502 690614
rect 529586 690378 529822 690614
rect 529266 670378 529502 670614
rect 529586 670378 529822 670614
rect 529266 650378 529502 650614
rect 529586 650378 529822 650614
rect 529266 630378 529502 630614
rect 529586 630378 529822 630614
rect 529266 610378 529502 610614
rect 529586 610378 529822 610614
rect 529266 590378 529502 590614
rect 529586 590378 529822 590614
rect 529266 570378 529502 570614
rect 529586 570378 529822 570614
rect 529266 550378 529502 550614
rect 529586 550378 529822 550614
rect 531826 705562 532062 705798
rect 532146 705562 532382 705798
rect 531826 705242 532062 705478
rect 532146 705242 532382 705478
rect 531826 693058 532062 693294
rect 532146 693058 532382 693294
rect 531826 673058 532062 673294
rect 532146 673058 532382 673294
rect 531826 653058 532062 653294
rect 532146 653058 532382 653294
rect 531826 633058 532062 633294
rect 532146 633058 532382 633294
rect 531826 613058 532062 613294
rect 532146 613058 532382 613294
rect 531826 593058 532062 593294
rect 532146 593058 532382 593294
rect 531826 573058 532062 573294
rect 532146 573058 532382 573294
rect 531826 553058 532062 553294
rect 532146 553058 532382 553294
rect 542986 711322 543222 711558
rect 543306 711322 543542 711558
rect 542986 711002 543222 711238
rect 543306 711002 543542 711238
rect 539266 709402 539502 709638
rect 539586 709402 539822 709638
rect 539266 709082 539502 709318
rect 539586 709082 539822 709318
rect 532986 694038 533222 694274
rect 533306 694038 533542 694274
rect 532986 674038 533222 674274
rect 533306 674038 533542 674274
rect 532986 654038 533222 654274
rect 533306 654038 533542 654274
rect 532986 634038 533222 634274
rect 533306 634038 533542 634274
rect 532986 614038 533222 614274
rect 533306 614038 533542 614274
rect 532986 594038 533222 594274
rect 533306 594038 533542 594274
rect 532986 574038 533222 574274
rect 533306 574038 533542 574274
rect 532986 554038 533222 554274
rect 533306 554038 533542 554274
rect 535546 707482 535782 707718
rect 535866 707482 536102 707718
rect 535546 707162 535782 707398
rect 535866 707162 536102 707398
rect 535546 696718 535782 696954
rect 535866 696718 536102 696954
rect 535546 676718 535782 676954
rect 535866 676718 536102 676954
rect 535546 656718 535782 656954
rect 535866 656718 536102 656954
rect 535546 636718 535782 636954
rect 535866 636718 536102 636954
rect 535546 616718 535782 616954
rect 535866 616718 536102 616954
rect 535546 596718 535782 596954
rect 535866 596718 536102 596954
rect 535546 576718 535782 576954
rect 535866 576718 536102 576954
rect 535546 556718 535782 556954
rect 535866 556718 536102 556954
rect 539266 700378 539502 700614
rect 539586 700378 539822 700614
rect 539266 680378 539502 680614
rect 539586 680378 539822 680614
rect 539266 660378 539502 660614
rect 539586 660378 539822 660614
rect 539266 640378 539502 640614
rect 539586 640378 539822 640614
rect 539266 620378 539502 620614
rect 539586 620378 539822 620614
rect 539266 600378 539502 600614
rect 539586 600378 539822 600614
rect 539266 580378 539502 580614
rect 539586 580378 539822 580614
rect 539266 560378 539502 560614
rect 539586 560378 539822 560614
rect 539266 540378 539502 540614
rect 539586 540378 539822 540614
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 683058 542062 683294
rect 542146 683058 542382 683294
rect 541826 663058 542062 663294
rect 542146 663058 542382 663294
rect 541826 643058 542062 643294
rect 542146 643058 542382 643294
rect 541826 623058 542062 623294
rect 542146 623058 542382 623294
rect 541826 603058 542062 603294
rect 542146 603058 542382 603294
rect 541826 583058 542062 583294
rect 542146 583058 542382 583294
rect 541826 563058 542062 563294
rect 542146 563058 542382 563294
rect 541826 543058 542062 543294
rect 542146 543058 542382 543294
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 542986 684038 543222 684274
rect 543306 684038 543542 684274
rect 542986 664038 543222 664274
rect 543306 664038 543542 664274
rect 542986 644038 543222 644274
rect 543306 644038 543542 644274
rect 542986 624038 543222 624274
rect 543306 624038 543542 624274
rect 542986 604038 543222 604274
rect 543306 604038 543542 604274
rect 542986 584038 543222 584274
rect 543306 584038 543542 584274
rect 542986 564038 543222 564274
rect 543306 564038 543542 564274
rect 542986 544038 543222 544274
rect 543306 544038 543542 544274
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 545546 686718 545782 686954
rect 545866 686718 546102 686954
rect 545546 666718 545782 666954
rect 545866 666718 546102 666954
rect 545546 646718 545782 646954
rect 545866 646718 546102 646954
rect 545546 626718 545782 626954
rect 545866 626718 546102 626954
rect 545546 606718 545782 606954
rect 545866 606718 546102 606954
rect 545546 586718 545782 586954
rect 545866 586718 546102 586954
rect 545546 566718 545782 566954
rect 545866 566718 546102 566954
rect 545546 546718 545782 546954
rect 545866 546718 546102 546954
rect 549266 690378 549502 690614
rect 549586 690378 549822 690614
rect 549266 670378 549502 670614
rect 549586 670378 549822 670614
rect 549266 650378 549502 650614
rect 549586 650378 549822 650614
rect 549266 630378 549502 630614
rect 549586 630378 549822 630614
rect 549266 610378 549502 610614
rect 549586 610378 549822 610614
rect 549266 590378 549502 590614
rect 549586 590378 549822 590614
rect 549266 570378 549502 570614
rect 549586 570378 549822 570614
rect 549266 550378 549502 550614
rect 549586 550378 549822 550614
rect 410328 533058 410564 533294
rect 546056 533058 546292 533294
rect 405546 526718 405782 526954
rect 405866 526718 406102 526954
rect 549266 530378 549502 530614
rect 549586 530378 549822 530614
rect 411008 523058 411244 523294
rect 545376 523058 545612 523294
rect 410328 513058 410564 513294
rect 546056 513058 546292 513294
rect 405546 506718 405782 506954
rect 405866 506718 406102 506954
rect 549266 510378 549502 510614
rect 549586 510378 549822 510614
rect 411008 503058 411244 503294
rect 545376 503058 545612 503294
rect 410328 493058 410564 493294
rect 546056 493058 546292 493294
rect 405546 486718 405782 486954
rect 405866 486718 406102 486954
rect 549266 490378 549502 490614
rect 549586 490378 549822 490614
rect 411008 483058 411244 483294
rect 545376 483058 545612 483294
rect 410328 473058 410564 473294
rect 546056 473058 546292 473294
rect 405546 466718 405782 466954
rect 405866 466718 406102 466954
rect 549266 470378 549502 470614
rect 549586 470378 549822 470614
rect 411008 463058 411244 463294
rect 545376 463058 545612 463294
rect 405546 446718 405782 446954
rect 405866 446718 406102 446954
rect 405546 426718 405782 426954
rect 405866 426718 406102 426954
rect 409266 450378 409502 450614
rect 409586 450378 409822 450614
rect 409266 430378 409502 430614
rect 409586 430378 409822 430614
rect 411826 433058 412062 433294
rect 412146 433058 412382 433294
rect 412986 434038 413222 434274
rect 413306 434038 413542 434274
rect 415546 436718 415782 436954
rect 415866 436718 416102 436954
rect 419266 440378 419502 440614
rect 419586 440378 419822 440614
rect 421826 443058 422062 443294
rect 422146 443058 422382 443294
rect 421826 423058 422062 423294
rect 422146 423058 422382 423294
rect 422986 444038 423222 444274
rect 423306 444038 423542 444274
rect 422986 424038 423222 424274
rect 423306 424038 423542 424274
rect 425546 446718 425782 446954
rect 425866 446718 426102 446954
rect 425546 426718 425782 426954
rect 425866 426718 426102 426954
rect 429266 450378 429502 450614
rect 429586 450378 429822 450614
rect 429266 430378 429502 430614
rect 429586 430378 429822 430614
rect 431826 433058 432062 433294
rect 432146 433058 432382 433294
rect 432986 434038 433222 434274
rect 433306 434038 433542 434274
rect 435546 436718 435782 436954
rect 435866 436718 436102 436954
rect 439266 440378 439502 440614
rect 439586 440378 439822 440614
rect 441826 443058 442062 443294
rect 442146 443058 442382 443294
rect 441826 423058 442062 423294
rect 442146 423058 442382 423294
rect 442986 444038 443222 444274
rect 443306 444038 443542 444274
rect 442986 424038 443222 424274
rect 443306 424038 443542 424274
rect 445546 446718 445782 446954
rect 445866 446718 446102 446954
rect 445546 426718 445782 426954
rect 445866 426718 446102 426954
rect 449266 450378 449502 450614
rect 449586 450378 449822 450614
rect 449266 430378 449502 430614
rect 449586 430378 449822 430614
rect 451826 433058 452062 433294
rect 452146 433058 452382 433294
rect 452986 434038 453222 434274
rect 453306 434038 453542 434274
rect 455546 436718 455782 436954
rect 455866 436718 456102 436954
rect 459266 440378 459502 440614
rect 459586 440378 459822 440614
rect 461826 443058 462062 443294
rect 462146 443058 462382 443294
rect 461826 423058 462062 423294
rect 462146 423058 462382 423294
rect 462986 444038 463222 444274
rect 463306 444038 463542 444274
rect 462986 424038 463222 424274
rect 463306 424038 463542 424274
rect 465546 446718 465782 446954
rect 465866 446718 466102 446954
rect 465546 426718 465782 426954
rect 465866 426718 466102 426954
rect 469266 450378 469502 450614
rect 469586 450378 469822 450614
rect 469266 430378 469502 430614
rect 469586 430378 469822 430614
rect 471826 433058 472062 433294
rect 472146 433058 472382 433294
rect 472986 434038 473222 434274
rect 473306 434038 473542 434274
rect 475546 436718 475782 436954
rect 475866 436718 476102 436954
rect 479266 440378 479502 440614
rect 479586 440378 479822 440614
rect 481826 443058 482062 443294
rect 482146 443058 482382 443294
rect 481826 423058 482062 423294
rect 482146 423058 482382 423294
rect 482986 444038 483222 444274
rect 483306 444038 483542 444274
rect 482986 424038 483222 424274
rect 483306 424038 483542 424274
rect 485546 446718 485782 446954
rect 485866 446718 486102 446954
rect 485546 426718 485782 426954
rect 485866 426718 486102 426954
rect 489266 450378 489502 450614
rect 489586 450378 489822 450614
rect 489266 430378 489502 430614
rect 489586 430378 489822 430614
rect 491826 433058 492062 433294
rect 492146 433058 492382 433294
rect 492986 434038 493222 434274
rect 493306 434038 493542 434274
rect 495546 436718 495782 436954
rect 495866 436718 496102 436954
rect 499266 440378 499502 440614
rect 499586 440378 499822 440614
rect 501826 443058 502062 443294
rect 502146 443058 502382 443294
rect 501826 423058 502062 423294
rect 502146 423058 502382 423294
rect 502986 444038 503222 444274
rect 503306 444038 503542 444274
rect 502986 424038 503222 424274
rect 503306 424038 503542 424274
rect 505546 446718 505782 446954
rect 505866 446718 506102 446954
rect 505546 426718 505782 426954
rect 505866 426718 506102 426954
rect 509266 450378 509502 450614
rect 509586 450378 509822 450614
rect 509266 430378 509502 430614
rect 509586 430378 509822 430614
rect 511826 433058 512062 433294
rect 512146 433058 512382 433294
rect 512986 434038 513222 434274
rect 513306 434038 513542 434274
rect 515546 436718 515782 436954
rect 515866 436718 516102 436954
rect 519266 440378 519502 440614
rect 519586 440378 519822 440614
rect 521826 443058 522062 443294
rect 522146 443058 522382 443294
rect 521826 423058 522062 423294
rect 522146 423058 522382 423294
rect 522986 444038 523222 444274
rect 523306 444038 523542 444274
rect 522986 424038 523222 424274
rect 523306 424038 523542 424274
rect 525546 446718 525782 446954
rect 525866 446718 526102 446954
rect 525546 426718 525782 426954
rect 525866 426718 526102 426954
rect 529266 450378 529502 450614
rect 529586 450378 529822 450614
rect 529266 430378 529502 430614
rect 529586 430378 529822 430614
rect 531826 433058 532062 433294
rect 532146 433058 532382 433294
rect 532986 434038 533222 434274
rect 533306 434038 533542 434274
rect 535546 436718 535782 436954
rect 535866 436718 536102 436954
rect 539266 440378 539502 440614
rect 539586 440378 539822 440614
rect 541826 443058 542062 443294
rect 542146 443058 542382 443294
rect 541826 423058 542062 423294
rect 542146 423058 542382 423294
rect 542986 444038 543222 444274
rect 543306 444038 543542 444274
rect 542986 424038 543222 424274
rect 543306 424038 543542 424274
rect 545546 446718 545782 446954
rect 545866 446718 546102 446954
rect 545546 426718 545782 426954
rect 545866 426718 546102 426954
rect 549266 450378 549502 450614
rect 549586 450378 549822 450614
rect 549266 430378 549502 430614
rect 549586 430378 549822 430614
rect 551826 705562 552062 705798
rect 552146 705562 552382 705798
rect 551826 705242 552062 705478
rect 552146 705242 552382 705478
rect 551826 693058 552062 693294
rect 552146 693058 552382 693294
rect 551826 673058 552062 673294
rect 552146 673058 552382 673294
rect 551826 653058 552062 653294
rect 552146 653058 552382 653294
rect 551826 633058 552062 633294
rect 552146 633058 552382 633294
rect 551826 613058 552062 613294
rect 552146 613058 552382 613294
rect 551826 593058 552062 593294
rect 552146 593058 552382 593294
rect 551826 573058 552062 573294
rect 552146 573058 552382 573294
rect 551826 553058 552062 553294
rect 552146 553058 552382 553294
rect 551826 533058 552062 533294
rect 552146 533058 552382 533294
rect 551826 513058 552062 513294
rect 552146 513058 552382 513294
rect 551826 493058 552062 493294
rect 552146 493058 552382 493294
rect 551826 473058 552062 473294
rect 552146 473058 552382 473294
rect 551826 453058 552062 453294
rect 552146 453058 552382 453294
rect 551826 433058 552062 433294
rect 552146 433058 552382 433294
rect 562986 711322 563222 711558
rect 563306 711322 563542 711558
rect 562986 711002 563222 711238
rect 563306 711002 563542 711238
rect 559266 709402 559502 709638
rect 559586 709402 559822 709638
rect 559266 709082 559502 709318
rect 559586 709082 559822 709318
rect 552986 694038 553222 694274
rect 553306 694038 553542 694274
rect 552986 674038 553222 674274
rect 553306 674038 553542 674274
rect 552986 654038 553222 654274
rect 553306 654038 553542 654274
rect 552986 634038 553222 634274
rect 553306 634038 553542 634274
rect 552986 614038 553222 614274
rect 553306 614038 553542 614274
rect 552986 594038 553222 594274
rect 553306 594038 553542 594274
rect 552986 574038 553222 574274
rect 553306 574038 553542 574274
rect 552986 554038 553222 554274
rect 553306 554038 553542 554274
rect 552986 534038 553222 534274
rect 553306 534038 553542 534274
rect 552986 514038 553222 514274
rect 553306 514038 553542 514274
rect 552986 494038 553222 494274
rect 553306 494038 553542 494274
rect 552986 474038 553222 474274
rect 553306 474038 553542 474274
rect 552986 454038 553222 454274
rect 553306 454038 553542 454274
rect 552986 434038 553222 434274
rect 553306 434038 553542 434274
rect 555546 707482 555782 707718
rect 555866 707482 556102 707718
rect 555546 707162 555782 707398
rect 555866 707162 556102 707398
rect 555546 696718 555782 696954
rect 555866 696718 556102 696954
rect 555546 676718 555782 676954
rect 555866 676718 556102 676954
rect 555546 656718 555782 656954
rect 555866 656718 556102 656954
rect 555546 636718 555782 636954
rect 555866 636718 556102 636954
rect 555546 616718 555782 616954
rect 555866 616718 556102 616954
rect 555546 596718 555782 596954
rect 555866 596718 556102 596954
rect 555546 576718 555782 576954
rect 555866 576718 556102 576954
rect 555546 556718 555782 556954
rect 555866 556718 556102 556954
rect 555546 536718 555782 536954
rect 555866 536718 556102 536954
rect 555546 516718 555782 516954
rect 555866 516718 556102 516954
rect 555546 496718 555782 496954
rect 555866 496718 556102 496954
rect 555546 476718 555782 476954
rect 555866 476718 556102 476954
rect 555546 456718 555782 456954
rect 555866 456718 556102 456954
rect 555546 436718 555782 436954
rect 555866 436718 556102 436954
rect 559266 700378 559502 700614
rect 559586 700378 559822 700614
rect 559266 680378 559502 680614
rect 559586 680378 559822 680614
rect 559266 660378 559502 660614
rect 559586 660378 559822 660614
rect 559266 640378 559502 640614
rect 559586 640378 559822 640614
rect 559266 620378 559502 620614
rect 559586 620378 559822 620614
rect 559266 600378 559502 600614
rect 559586 600378 559822 600614
rect 559266 580378 559502 580614
rect 559586 580378 559822 580614
rect 559266 560378 559502 560614
rect 559586 560378 559822 560614
rect 559266 540378 559502 540614
rect 559586 540378 559822 540614
rect 559266 520378 559502 520614
rect 559586 520378 559822 520614
rect 559266 500378 559502 500614
rect 559586 500378 559822 500614
rect 559266 480378 559502 480614
rect 559586 480378 559822 480614
rect 559266 460378 559502 460614
rect 559586 460378 559822 460614
rect 559266 440378 559502 440614
rect 559586 440378 559822 440614
rect 559266 420378 559502 420614
rect 559586 420378 559822 420614
rect 219610 413058 219846 413294
rect 250330 413058 250566 413294
rect 281050 413058 281286 413294
rect 311770 413058 312006 413294
rect 342490 413058 342726 413294
rect 373210 413058 373446 413294
rect 403930 413058 404166 413294
rect 434650 413058 434886 413294
rect 465370 413058 465606 413294
rect 496090 413058 496326 413294
rect 526810 413058 527046 413294
rect 204250 403058 204486 403294
rect 234970 403058 235206 403294
rect 265690 403058 265926 403294
rect 296410 403058 296646 403294
rect 327130 403058 327366 403294
rect 357850 403058 358086 403294
rect 388570 403058 388806 403294
rect 419290 403058 419526 403294
rect 450010 403058 450246 403294
rect 480730 403058 480966 403294
rect 511450 403058 511686 403294
rect 542170 403058 542406 403294
rect 559266 400378 559502 400614
rect 559586 400378 559822 400614
rect 219610 393058 219846 393294
rect 250330 393058 250566 393294
rect 281050 393058 281286 393294
rect 311770 393058 312006 393294
rect 342490 393058 342726 393294
rect 373210 393058 373446 393294
rect 403930 393058 404166 393294
rect 434650 393058 434886 393294
rect 465370 393058 465606 393294
rect 496090 393058 496326 393294
rect 526810 393058 527046 393294
rect 204250 383058 204486 383294
rect 234970 383058 235206 383294
rect 265690 383058 265926 383294
rect 296410 383058 296646 383294
rect 327130 383058 327366 383294
rect 357850 383058 358086 383294
rect 388570 383058 388806 383294
rect 419290 383058 419526 383294
rect 450010 383058 450246 383294
rect 480730 383058 480966 383294
rect 511450 383058 511686 383294
rect 542170 383058 542406 383294
rect 559266 380378 559502 380614
rect 559586 380378 559822 380614
rect 219610 373058 219846 373294
rect 250330 373058 250566 373294
rect 281050 373058 281286 373294
rect 311770 373058 312006 373294
rect 342490 373058 342726 373294
rect 373210 373058 373446 373294
rect 403930 373058 404166 373294
rect 434650 373058 434886 373294
rect 465370 373058 465606 373294
rect 496090 373058 496326 373294
rect 526810 373058 527046 373294
rect 204250 363058 204486 363294
rect 234970 363058 235206 363294
rect 265690 363058 265926 363294
rect 296410 363058 296646 363294
rect 327130 363058 327366 363294
rect 357850 363058 358086 363294
rect 388570 363058 388806 363294
rect 419290 363058 419526 363294
rect 450010 363058 450246 363294
rect 480730 363058 480966 363294
rect 511450 363058 511686 363294
rect 542170 363058 542406 363294
rect 559266 360378 559502 360614
rect 559586 360378 559822 360614
rect 219610 353058 219846 353294
rect 250330 353058 250566 353294
rect 281050 353058 281286 353294
rect 311770 353058 312006 353294
rect 342490 353058 342726 353294
rect 373210 353058 373446 353294
rect 403930 353058 404166 353294
rect 434650 353058 434886 353294
rect 465370 353058 465606 353294
rect 496090 353058 496326 353294
rect 526810 353058 527046 353294
rect 204250 343058 204486 343294
rect 234970 343058 235206 343294
rect 265690 343058 265926 343294
rect 296410 343058 296646 343294
rect 327130 343058 327366 343294
rect 357850 343058 358086 343294
rect 388570 343058 388806 343294
rect 419290 343058 419526 343294
rect 450010 343058 450246 343294
rect 480730 343058 480966 343294
rect 511450 343058 511686 343294
rect 542170 343058 542406 343294
rect 559266 340378 559502 340614
rect 559586 340378 559822 340614
rect 219610 333058 219846 333294
rect 250330 333058 250566 333294
rect 281050 333058 281286 333294
rect 311770 333058 312006 333294
rect 342490 333058 342726 333294
rect 373210 333058 373446 333294
rect 403930 333058 404166 333294
rect 434650 333058 434886 333294
rect 465370 333058 465606 333294
rect 496090 333058 496326 333294
rect 526810 333058 527046 333294
rect 204250 323058 204486 323294
rect 234970 323058 235206 323294
rect 265690 323058 265926 323294
rect 296410 323058 296646 323294
rect 327130 323058 327366 323294
rect 357850 323058 358086 323294
rect 388570 323058 388806 323294
rect 419290 323058 419526 323294
rect 450010 323058 450246 323294
rect 480730 323058 480966 323294
rect 511450 323058 511686 323294
rect 542170 323058 542406 323294
rect 559266 320378 559502 320614
rect 559586 320378 559822 320614
rect 219610 313058 219846 313294
rect 250330 313058 250566 313294
rect 281050 313058 281286 313294
rect 311770 313058 312006 313294
rect 342490 313058 342726 313294
rect 373210 313058 373446 313294
rect 403930 313058 404166 313294
rect 434650 313058 434886 313294
rect 465370 313058 465606 313294
rect 496090 313058 496326 313294
rect 526810 313058 527046 313294
rect 204250 303058 204486 303294
rect 234970 303058 235206 303294
rect 265690 303058 265926 303294
rect 296410 303058 296646 303294
rect 327130 303058 327366 303294
rect 357850 303058 358086 303294
rect 388570 303058 388806 303294
rect 419290 303058 419526 303294
rect 450010 303058 450246 303294
rect 480730 303058 480966 303294
rect 511450 303058 511686 303294
rect 542170 303058 542406 303294
rect 559266 300378 559502 300614
rect 559586 300378 559822 300614
rect 219610 293058 219846 293294
rect 250330 293058 250566 293294
rect 281050 293058 281286 293294
rect 311770 293058 312006 293294
rect 342490 293058 342726 293294
rect 373210 293058 373446 293294
rect 403930 293058 404166 293294
rect 434650 293058 434886 293294
rect 465370 293058 465606 293294
rect 496090 293058 496326 293294
rect 526810 293058 527046 293294
rect 204250 283058 204486 283294
rect 234970 283058 235206 283294
rect 265690 283058 265926 283294
rect 296410 283058 296646 283294
rect 327130 283058 327366 283294
rect 357850 283058 358086 283294
rect 388570 283058 388806 283294
rect 419290 283058 419526 283294
rect 450010 283058 450246 283294
rect 480730 283058 480966 283294
rect 511450 283058 511686 283294
rect 542170 283058 542406 283294
rect 559266 280378 559502 280614
rect 559586 280378 559822 280614
rect 219610 273058 219846 273294
rect 250330 273058 250566 273294
rect 281050 273058 281286 273294
rect 311770 273058 312006 273294
rect 342490 273058 342726 273294
rect 373210 273058 373446 273294
rect 403930 273058 404166 273294
rect 434650 273058 434886 273294
rect 465370 273058 465606 273294
rect 496090 273058 496326 273294
rect 526810 273058 527046 273294
rect 204250 263058 204486 263294
rect 234970 263058 235206 263294
rect 265690 263058 265926 263294
rect 296410 263058 296646 263294
rect 327130 263058 327366 263294
rect 357850 263058 358086 263294
rect 388570 263058 388806 263294
rect 419290 263058 419526 263294
rect 450010 263058 450246 263294
rect 480730 263058 480966 263294
rect 511450 263058 511686 263294
rect 542170 263058 542406 263294
rect 559266 260378 559502 260614
rect 559586 260378 559822 260614
rect 219610 253058 219846 253294
rect 250330 253058 250566 253294
rect 281050 253058 281286 253294
rect 311770 253058 312006 253294
rect 342490 253058 342726 253294
rect 373210 253058 373446 253294
rect 403930 253058 404166 253294
rect 434650 253058 434886 253294
rect 465370 253058 465606 253294
rect 496090 253058 496326 253294
rect 526810 253058 527046 253294
rect 204250 243058 204486 243294
rect 234970 243058 235206 243294
rect 265690 243058 265926 243294
rect 296410 243058 296646 243294
rect 327130 243058 327366 243294
rect 357850 243058 358086 243294
rect 388570 243058 388806 243294
rect 419290 243058 419526 243294
rect 450010 243058 450246 243294
rect 480730 243058 480966 243294
rect 511450 243058 511686 243294
rect 542170 243058 542406 243294
rect 195546 236718 195782 236954
rect 195866 236718 196102 236954
rect 559266 240378 559502 240614
rect 559586 240378 559822 240614
rect 219610 233058 219846 233294
rect 250330 233058 250566 233294
rect 281050 233058 281286 233294
rect 311770 233058 312006 233294
rect 342490 233058 342726 233294
rect 373210 233058 373446 233294
rect 403930 233058 404166 233294
rect 434650 233058 434886 233294
rect 465370 233058 465606 233294
rect 496090 233058 496326 233294
rect 526810 233058 527046 233294
rect 204250 223058 204486 223294
rect 234970 223058 235206 223294
rect 265690 223058 265926 223294
rect 296410 223058 296646 223294
rect 327130 223058 327366 223294
rect 357850 223058 358086 223294
rect 388570 223058 388806 223294
rect 419290 223058 419526 223294
rect 450010 223058 450246 223294
rect 480730 223058 480966 223294
rect 511450 223058 511686 223294
rect 542170 223058 542406 223294
rect 195546 216718 195782 216954
rect 195866 216718 196102 216954
rect 559266 220378 559502 220614
rect 559586 220378 559822 220614
rect 219610 213058 219846 213294
rect 250330 213058 250566 213294
rect 281050 213058 281286 213294
rect 311770 213058 312006 213294
rect 342490 213058 342726 213294
rect 373210 213058 373446 213294
rect 403930 213058 404166 213294
rect 434650 213058 434886 213294
rect 465370 213058 465606 213294
rect 496090 213058 496326 213294
rect 526810 213058 527046 213294
rect 204250 203058 204486 203294
rect 234970 203058 235206 203294
rect 265690 203058 265926 203294
rect 296410 203058 296646 203294
rect 327130 203058 327366 203294
rect 357850 203058 358086 203294
rect 388570 203058 388806 203294
rect 419290 203058 419526 203294
rect 450010 203058 450246 203294
rect 480730 203058 480966 203294
rect 511450 203058 511686 203294
rect 542170 203058 542406 203294
rect 195546 196718 195782 196954
rect 195866 196718 196102 196954
rect 559266 200378 559502 200614
rect 559586 200378 559822 200614
rect 219610 193058 219846 193294
rect 250330 193058 250566 193294
rect 281050 193058 281286 193294
rect 311770 193058 312006 193294
rect 342490 193058 342726 193294
rect 373210 193058 373446 193294
rect 403930 193058 404166 193294
rect 434650 193058 434886 193294
rect 465370 193058 465606 193294
rect 496090 193058 496326 193294
rect 526810 193058 527046 193294
rect 204250 183058 204486 183294
rect 234970 183058 235206 183294
rect 265690 183058 265926 183294
rect 296410 183058 296646 183294
rect 327130 183058 327366 183294
rect 357850 183058 358086 183294
rect 388570 183058 388806 183294
rect 419290 183058 419526 183294
rect 450010 183058 450246 183294
rect 480730 183058 480966 183294
rect 511450 183058 511686 183294
rect 542170 183058 542406 183294
rect 195546 176718 195782 176954
rect 195866 176718 196102 176954
rect 559266 180378 559502 180614
rect 559586 180378 559822 180614
rect 219610 173058 219846 173294
rect 250330 173058 250566 173294
rect 281050 173058 281286 173294
rect 311770 173058 312006 173294
rect 342490 173058 342726 173294
rect 373210 173058 373446 173294
rect 403930 173058 404166 173294
rect 434650 173058 434886 173294
rect 465370 173058 465606 173294
rect 496090 173058 496326 173294
rect 526810 173058 527046 173294
rect 204250 163058 204486 163294
rect 234970 163058 235206 163294
rect 265690 163058 265926 163294
rect 296410 163058 296646 163294
rect 327130 163058 327366 163294
rect 357850 163058 358086 163294
rect 388570 163058 388806 163294
rect 419290 163058 419526 163294
rect 450010 163058 450246 163294
rect 480730 163058 480966 163294
rect 511450 163058 511686 163294
rect 542170 163058 542406 163294
rect 195546 156718 195782 156954
rect 195866 156718 196102 156954
rect 559266 160378 559502 160614
rect 559586 160378 559822 160614
rect 219610 153058 219846 153294
rect 250330 153058 250566 153294
rect 281050 153058 281286 153294
rect 311770 153058 312006 153294
rect 342490 153058 342726 153294
rect 373210 153058 373446 153294
rect 403930 153058 404166 153294
rect 434650 153058 434886 153294
rect 465370 153058 465606 153294
rect 496090 153058 496326 153294
rect 526810 153058 527046 153294
rect 204250 143058 204486 143294
rect 234970 143058 235206 143294
rect 265690 143058 265926 143294
rect 296410 143058 296646 143294
rect 327130 143058 327366 143294
rect 357850 143058 358086 143294
rect 388570 143058 388806 143294
rect 419290 143058 419526 143294
rect 450010 143058 450246 143294
rect 480730 143058 480966 143294
rect 511450 143058 511686 143294
rect 542170 143058 542406 143294
rect 195546 136718 195782 136954
rect 195866 136718 196102 136954
rect 559266 140378 559502 140614
rect 559586 140378 559822 140614
rect 219610 133058 219846 133294
rect 250330 133058 250566 133294
rect 281050 133058 281286 133294
rect 311770 133058 312006 133294
rect 342490 133058 342726 133294
rect 373210 133058 373446 133294
rect 403930 133058 404166 133294
rect 434650 133058 434886 133294
rect 465370 133058 465606 133294
rect 496090 133058 496326 133294
rect 526810 133058 527046 133294
rect 204250 123058 204486 123294
rect 234970 123058 235206 123294
rect 265690 123058 265926 123294
rect 296410 123058 296646 123294
rect 327130 123058 327366 123294
rect 357850 123058 358086 123294
rect 388570 123058 388806 123294
rect 419290 123058 419526 123294
rect 450010 123058 450246 123294
rect 480730 123058 480966 123294
rect 511450 123058 511686 123294
rect 542170 123058 542406 123294
rect 195546 116718 195782 116954
rect 195866 116718 196102 116954
rect 559266 120378 559502 120614
rect 559586 120378 559822 120614
rect 219610 113058 219846 113294
rect 250330 113058 250566 113294
rect 281050 113058 281286 113294
rect 311770 113058 312006 113294
rect 342490 113058 342726 113294
rect 373210 113058 373446 113294
rect 403930 113058 404166 113294
rect 434650 113058 434886 113294
rect 465370 113058 465606 113294
rect 496090 113058 496326 113294
rect 526810 113058 527046 113294
rect 204250 103058 204486 103294
rect 234970 103058 235206 103294
rect 265690 103058 265926 103294
rect 296410 103058 296646 103294
rect 327130 103058 327366 103294
rect 357850 103058 358086 103294
rect 388570 103058 388806 103294
rect 419290 103058 419526 103294
rect 450010 103058 450246 103294
rect 480730 103058 480966 103294
rect 511450 103058 511686 103294
rect 542170 103058 542406 103294
rect 195546 96718 195782 96954
rect 195866 96718 196102 96954
rect 559266 100378 559502 100614
rect 559586 100378 559822 100614
rect 219610 93058 219846 93294
rect 250330 93058 250566 93294
rect 281050 93058 281286 93294
rect 311770 93058 312006 93294
rect 342490 93058 342726 93294
rect 373210 93058 373446 93294
rect 403930 93058 404166 93294
rect 434650 93058 434886 93294
rect 465370 93058 465606 93294
rect 496090 93058 496326 93294
rect 526810 93058 527046 93294
rect 204250 83058 204486 83294
rect 234970 83058 235206 83294
rect 265690 83058 265926 83294
rect 296410 83058 296646 83294
rect 327130 83058 327366 83294
rect 357850 83058 358086 83294
rect 388570 83058 388806 83294
rect 419290 83058 419526 83294
rect 450010 83058 450246 83294
rect 480730 83058 480966 83294
rect 511450 83058 511686 83294
rect 542170 83058 542406 83294
rect 195546 76718 195782 76954
rect 195866 76718 196102 76954
rect 559266 80378 559502 80614
rect 559586 80378 559822 80614
rect 219610 73058 219846 73294
rect 250330 73058 250566 73294
rect 281050 73058 281286 73294
rect 311770 73058 312006 73294
rect 342490 73058 342726 73294
rect 373210 73058 373446 73294
rect 403930 73058 404166 73294
rect 434650 73058 434886 73294
rect 465370 73058 465606 73294
rect 496090 73058 496326 73294
rect 526810 73058 527046 73294
rect 204250 63058 204486 63294
rect 234970 63058 235206 63294
rect 265690 63058 265926 63294
rect 296410 63058 296646 63294
rect 327130 63058 327366 63294
rect 357850 63058 358086 63294
rect 388570 63058 388806 63294
rect 419290 63058 419526 63294
rect 450010 63058 450246 63294
rect 480730 63058 480966 63294
rect 511450 63058 511686 63294
rect 542170 63058 542406 63294
rect 559266 60378 559502 60614
rect 559586 60378 559822 60614
rect 195546 56718 195782 56954
rect 195866 56718 196102 56954
rect 195546 36718 195782 36954
rect 195866 36718 196102 36954
rect 195546 16718 195782 16954
rect 195866 16718 196102 16954
rect 195546 -3462 195782 -3226
rect 195866 -3462 196102 -3226
rect 195546 -3782 195782 -3546
rect 195866 -3782 196102 -3546
rect 199266 40378 199502 40614
rect 199586 40378 199822 40614
rect 199266 20378 199502 20614
rect 199586 20378 199822 20614
rect 201826 43058 202062 43294
rect 202146 43058 202382 43294
rect 201826 23058 202062 23294
rect 202146 23058 202382 23294
rect 201826 3058 202062 3294
rect 202146 3058 202382 3294
rect 201826 -582 202062 -346
rect 202146 -582 202382 -346
rect 201826 -902 202062 -666
rect 202146 -902 202382 -666
rect 202986 44038 203222 44274
rect 203306 44038 203542 44274
rect 202986 24038 203222 24274
rect 203306 24038 203542 24274
rect 199266 -5382 199502 -5146
rect 199586 -5382 199822 -5146
rect 199266 -5702 199502 -5466
rect 199586 -5702 199822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 205546 46718 205782 46954
rect 205866 46718 206102 46954
rect 205546 26718 205782 26954
rect 205866 26718 206102 26954
rect 205546 6718 205782 6954
rect 205866 6718 206102 6954
rect 205546 -2502 205782 -2266
rect 205866 -2502 206102 -2266
rect 205546 -2822 205782 -2586
rect 205866 -2822 206102 -2586
rect 209266 50378 209502 50614
rect 209586 50378 209822 50614
rect 209266 30378 209502 30614
rect 209586 30378 209822 30614
rect 209266 10378 209502 10614
rect 209586 10378 209822 10614
rect 211826 53058 212062 53294
rect 212146 53058 212382 53294
rect 211826 33058 212062 33294
rect 212146 33058 212382 33294
rect 211826 13058 212062 13294
rect 212146 13058 212382 13294
rect 211826 -1542 212062 -1306
rect 212146 -1542 212382 -1306
rect 211826 -1862 212062 -1626
rect 212146 -1862 212382 -1626
rect 212986 54038 213222 54274
rect 213306 54038 213542 54274
rect 212986 34038 213222 34274
rect 213306 34038 213542 34274
rect 212986 14038 213222 14274
rect 213306 14038 213542 14274
rect 209266 -4422 209502 -4186
rect 209586 -4422 209822 -4186
rect 209266 -4742 209502 -4506
rect 209586 -4742 209822 -4506
rect 202986 -7302 203222 -7066
rect 203306 -7302 203542 -7066
rect 202986 -7622 203222 -7386
rect 203306 -7622 203542 -7386
rect 215546 56718 215782 56954
rect 215866 56718 216102 56954
rect 215546 36718 215782 36954
rect 215866 36718 216102 36954
rect 215546 16718 215782 16954
rect 215866 16718 216102 16954
rect 215546 -3462 215782 -3226
rect 215866 -3462 216102 -3226
rect 215546 -3782 215782 -3546
rect 215866 -3782 216102 -3546
rect 219266 40378 219502 40614
rect 219586 40378 219822 40614
rect 219266 20378 219502 20614
rect 219586 20378 219822 20614
rect 221826 43058 222062 43294
rect 222146 43058 222382 43294
rect 221826 23058 222062 23294
rect 222146 23058 222382 23294
rect 221826 3058 222062 3294
rect 222146 3058 222382 3294
rect 221826 -582 222062 -346
rect 222146 -582 222382 -346
rect 221826 -902 222062 -666
rect 222146 -902 222382 -666
rect 222986 44038 223222 44274
rect 223306 44038 223542 44274
rect 222986 24038 223222 24274
rect 223306 24038 223542 24274
rect 219266 -5382 219502 -5146
rect 219586 -5382 219822 -5146
rect 219266 -5702 219502 -5466
rect 219586 -5702 219822 -5466
rect 212986 -6342 213222 -6106
rect 213306 -6342 213542 -6106
rect 212986 -6662 213222 -6426
rect 213306 -6662 213542 -6426
rect 225546 46718 225782 46954
rect 225866 46718 226102 46954
rect 225546 26718 225782 26954
rect 225866 26718 226102 26954
rect 225546 6718 225782 6954
rect 225866 6718 226102 6954
rect 225546 -2502 225782 -2266
rect 225866 -2502 226102 -2266
rect 225546 -2822 225782 -2586
rect 225866 -2822 226102 -2586
rect 229266 50378 229502 50614
rect 229586 50378 229822 50614
rect 229266 30378 229502 30614
rect 229586 30378 229822 30614
rect 229266 10378 229502 10614
rect 229586 10378 229822 10614
rect 231826 53058 232062 53294
rect 232146 53058 232382 53294
rect 231826 33058 232062 33294
rect 232146 33058 232382 33294
rect 231826 13058 232062 13294
rect 232146 13058 232382 13294
rect 231826 -1542 232062 -1306
rect 232146 -1542 232382 -1306
rect 231826 -1862 232062 -1626
rect 232146 -1862 232382 -1626
rect 232986 54038 233222 54274
rect 233306 54038 233542 54274
rect 232986 34038 233222 34274
rect 233306 34038 233542 34274
rect 232986 14038 233222 14274
rect 233306 14038 233542 14274
rect 229266 -4422 229502 -4186
rect 229586 -4422 229822 -4186
rect 229266 -4742 229502 -4506
rect 229586 -4742 229822 -4506
rect 222986 -7302 223222 -7066
rect 223306 -7302 223542 -7066
rect 222986 -7622 223222 -7386
rect 223306 -7622 223542 -7386
rect 235546 56718 235782 56954
rect 235866 56718 236102 56954
rect 235546 36718 235782 36954
rect 235866 36718 236102 36954
rect 235546 16718 235782 16954
rect 235866 16718 236102 16954
rect 235546 -3462 235782 -3226
rect 235866 -3462 236102 -3226
rect 235546 -3782 235782 -3546
rect 235866 -3782 236102 -3546
rect 239266 40378 239502 40614
rect 239586 40378 239822 40614
rect 239266 20378 239502 20614
rect 239586 20378 239822 20614
rect 241826 43058 242062 43294
rect 242146 43058 242382 43294
rect 241826 23058 242062 23294
rect 242146 23058 242382 23294
rect 241826 3058 242062 3294
rect 242146 3058 242382 3294
rect 241826 -582 242062 -346
rect 242146 -582 242382 -346
rect 241826 -902 242062 -666
rect 242146 -902 242382 -666
rect 242986 44038 243222 44274
rect 243306 44038 243542 44274
rect 242986 24038 243222 24274
rect 243306 24038 243542 24274
rect 239266 -5382 239502 -5146
rect 239586 -5382 239822 -5146
rect 239266 -5702 239502 -5466
rect 239586 -5702 239822 -5466
rect 232986 -6342 233222 -6106
rect 233306 -6342 233542 -6106
rect 232986 -6662 233222 -6426
rect 233306 -6662 233542 -6426
rect 245546 46718 245782 46954
rect 245866 46718 246102 46954
rect 245546 26718 245782 26954
rect 245866 26718 246102 26954
rect 245546 6718 245782 6954
rect 245866 6718 246102 6954
rect 245546 -2502 245782 -2266
rect 245866 -2502 246102 -2266
rect 245546 -2822 245782 -2586
rect 245866 -2822 246102 -2586
rect 249266 50378 249502 50614
rect 249586 50378 249822 50614
rect 249266 30378 249502 30614
rect 249586 30378 249822 30614
rect 249266 10378 249502 10614
rect 249586 10378 249822 10614
rect 251826 53058 252062 53294
rect 252146 53058 252382 53294
rect 251826 33058 252062 33294
rect 252146 33058 252382 33294
rect 251826 13058 252062 13294
rect 252146 13058 252382 13294
rect 251826 -1542 252062 -1306
rect 252146 -1542 252382 -1306
rect 251826 -1862 252062 -1626
rect 252146 -1862 252382 -1626
rect 252986 54038 253222 54274
rect 253306 54038 253542 54274
rect 252986 34038 253222 34274
rect 253306 34038 253542 34274
rect 252986 14038 253222 14274
rect 253306 14038 253542 14274
rect 249266 -4422 249502 -4186
rect 249586 -4422 249822 -4186
rect 249266 -4742 249502 -4506
rect 249586 -4742 249822 -4506
rect 242986 -7302 243222 -7066
rect 243306 -7302 243542 -7066
rect 242986 -7622 243222 -7386
rect 243306 -7622 243542 -7386
rect 255546 56718 255782 56954
rect 255866 56718 256102 56954
rect 255546 36718 255782 36954
rect 255866 36718 256102 36954
rect 255546 16718 255782 16954
rect 255866 16718 256102 16954
rect 255546 -3462 255782 -3226
rect 255866 -3462 256102 -3226
rect 255546 -3782 255782 -3546
rect 255866 -3782 256102 -3546
rect 259266 40378 259502 40614
rect 259586 40378 259822 40614
rect 259266 20378 259502 20614
rect 259586 20378 259822 20614
rect 261826 43058 262062 43294
rect 262146 43058 262382 43294
rect 261826 23058 262062 23294
rect 262146 23058 262382 23294
rect 261826 3058 262062 3294
rect 262146 3058 262382 3294
rect 261826 -582 262062 -346
rect 262146 -582 262382 -346
rect 261826 -902 262062 -666
rect 262146 -902 262382 -666
rect 262986 44038 263222 44274
rect 263306 44038 263542 44274
rect 262986 24038 263222 24274
rect 263306 24038 263542 24274
rect 259266 -5382 259502 -5146
rect 259586 -5382 259822 -5146
rect 259266 -5702 259502 -5466
rect 259586 -5702 259822 -5466
rect 252986 -6342 253222 -6106
rect 253306 -6342 253542 -6106
rect 252986 -6662 253222 -6426
rect 253306 -6662 253542 -6426
rect 265546 46718 265782 46954
rect 265866 46718 266102 46954
rect 265546 26718 265782 26954
rect 265866 26718 266102 26954
rect 265546 6718 265782 6954
rect 265866 6718 266102 6954
rect 265546 -2502 265782 -2266
rect 265866 -2502 266102 -2266
rect 265546 -2822 265782 -2586
rect 265866 -2822 266102 -2586
rect 269266 50378 269502 50614
rect 269586 50378 269822 50614
rect 269266 30378 269502 30614
rect 269586 30378 269822 30614
rect 269266 10378 269502 10614
rect 269586 10378 269822 10614
rect 271826 53058 272062 53294
rect 272146 53058 272382 53294
rect 271826 33058 272062 33294
rect 272146 33058 272382 33294
rect 271826 13058 272062 13294
rect 272146 13058 272382 13294
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 272986 54038 273222 54274
rect 273306 54038 273542 54274
rect 272986 34038 273222 34274
rect 273306 34038 273542 34274
rect 272986 14038 273222 14274
rect 273306 14038 273542 14274
rect 269266 -4422 269502 -4186
rect 269586 -4422 269822 -4186
rect 269266 -4742 269502 -4506
rect 269586 -4742 269822 -4506
rect 262986 -7302 263222 -7066
rect 263306 -7302 263542 -7066
rect 262986 -7622 263222 -7386
rect 263306 -7622 263542 -7386
rect 275546 56718 275782 56954
rect 275866 56718 276102 56954
rect 275546 36718 275782 36954
rect 275866 36718 276102 36954
rect 275546 16718 275782 16954
rect 275866 16718 276102 16954
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 40378 279502 40614
rect 279586 40378 279822 40614
rect 279266 20378 279502 20614
rect 279586 20378 279822 20614
rect 281826 43058 282062 43294
rect 282146 43058 282382 43294
rect 281826 23058 282062 23294
rect 282146 23058 282382 23294
rect 281826 3058 282062 3294
rect 282146 3058 282382 3294
rect 281826 -582 282062 -346
rect 282146 -582 282382 -346
rect 281826 -902 282062 -666
rect 282146 -902 282382 -666
rect 282986 44038 283222 44274
rect 283306 44038 283542 44274
rect 282986 24038 283222 24274
rect 283306 24038 283542 24274
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 272986 -6342 273222 -6106
rect 273306 -6342 273542 -6106
rect 272986 -6662 273222 -6426
rect 273306 -6662 273542 -6426
rect 285546 46718 285782 46954
rect 285866 46718 286102 46954
rect 285546 26718 285782 26954
rect 285866 26718 286102 26954
rect 285546 6718 285782 6954
rect 285866 6718 286102 6954
rect 285546 -2502 285782 -2266
rect 285866 -2502 286102 -2266
rect 285546 -2822 285782 -2586
rect 285866 -2822 286102 -2586
rect 289266 50378 289502 50614
rect 289586 50378 289822 50614
rect 289266 30378 289502 30614
rect 289586 30378 289822 30614
rect 289266 10378 289502 10614
rect 289586 10378 289822 10614
rect 291826 53058 292062 53294
rect 292146 53058 292382 53294
rect 291826 33058 292062 33294
rect 292146 33058 292382 33294
rect 291826 13058 292062 13294
rect 292146 13058 292382 13294
rect 291826 -1542 292062 -1306
rect 292146 -1542 292382 -1306
rect 291826 -1862 292062 -1626
rect 292146 -1862 292382 -1626
rect 292986 54038 293222 54274
rect 293306 54038 293542 54274
rect 292986 34038 293222 34274
rect 293306 34038 293542 34274
rect 292986 14038 293222 14274
rect 293306 14038 293542 14274
rect 289266 -4422 289502 -4186
rect 289586 -4422 289822 -4186
rect 289266 -4742 289502 -4506
rect 289586 -4742 289822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 295546 56718 295782 56954
rect 295866 56718 296102 56954
rect 295546 36718 295782 36954
rect 295866 36718 296102 36954
rect 295546 16718 295782 16954
rect 295866 16718 296102 16954
rect 295546 -3462 295782 -3226
rect 295866 -3462 296102 -3226
rect 295546 -3782 295782 -3546
rect 295866 -3782 296102 -3546
rect 299266 40378 299502 40614
rect 299586 40378 299822 40614
rect 299266 20378 299502 20614
rect 299586 20378 299822 20614
rect 301826 43058 302062 43294
rect 302146 43058 302382 43294
rect 301826 23058 302062 23294
rect 302146 23058 302382 23294
rect 301826 3058 302062 3294
rect 302146 3058 302382 3294
rect 301826 -582 302062 -346
rect 302146 -582 302382 -346
rect 301826 -902 302062 -666
rect 302146 -902 302382 -666
rect 302986 44038 303222 44274
rect 303306 44038 303542 44274
rect 302986 24038 303222 24274
rect 303306 24038 303542 24274
rect 299266 -5382 299502 -5146
rect 299586 -5382 299822 -5146
rect 299266 -5702 299502 -5466
rect 299586 -5702 299822 -5466
rect 292986 -6342 293222 -6106
rect 293306 -6342 293542 -6106
rect 292986 -6662 293222 -6426
rect 293306 -6662 293542 -6426
rect 305546 46718 305782 46954
rect 305866 46718 306102 46954
rect 305546 26718 305782 26954
rect 305866 26718 306102 26954
rect 305546 6718 305782 6954
rect 305866 6718 306102 6954
rect 305546 -2502 305782 -2266
rect 305866 -2502 306102 -2266
rect 305546 -2822 305782 -2586
rect 305866 -2822 306102 -2586
rect 309266 50378 309502 50614
rect 309586 50378 309822 50614
rect 309266 30378 309502 30614
rect 309586 30378 309822 30614
rect 309266 10378 309502 10614
rect 309586 10378 309822 10614
rect 311826 53058 312062 53294
rect 312146 53058 312382 53294
rect 311826 33058 312062 33294
rect 312146 33058 312382 33294
rect 311826 13058 312062 13294
rect 312146 13058 312382 13294
rect 311826 -1542 312062 -1306
rect 312146 -1542 312382 -1306
rect 311826 -1862 312062 -1626
rect 312146 -1862 312382 -1626
rect 312986 54038 313222 54274
rect 313306 54038 313542 54274
rect 312986 34038 313222 34274
rect 313306 34038 313542 34274
rect 312986 14038 313222 14274
rect 313306 14038 313542 14274
rect 309266 -4422 309502 -4186
rect 309586 -4422 309822 -4186
rect 309266 -4742 309502 -4506
rect 309586 -4742 309822 -4506
rect 302986 -7302 303222 -7066
rect 303306 -7302 303542 -7066
rect 302986 -7622 303222 -7386
rect 303306 -7622 303542 -7386
rect 315546 56718 315782 56954
rect 315866 56718 316102 56954
rect 315546 36718 315782 36954
rect 315866 36718 316102 36954
rect 315546 16718 315782 16954
rect 315866 16718 316102 16954
rect 315546 -3462 315782 -3226
rect 315866 -3462 316102 -3226
rect 315546 -3782 315782 -3546
rect 315866 -3782 316102 -3546
rect 319266 40378 319502 40614
rect 319586 40378 319822 40614
rect 319266 20378 319502 20614
rect 319586 20378 319822 20614
rect 321826 43058 322062 43294
rect 322146 43058 322382 43294
rect 321826 23058 322062 23294
rect 322146 23058 322382 23294
rect 321826 3058 322062 3294
rect 322146 3058 322382 3294
rect 321826 -582 322062 -346
rect 322146 -582 322382 -346
rect 321826 -902 322062 -666
rect 322146 -902 322382 -666
rect 322986 44038 323222 44274
rect 323306 44038 323542 44274
rect 322986 24038 323222 24274
rect 323306 24038 323542 24274
rect 319266 -5382 319502 -5146
rect 319586 -5382 319822 -5146
rect 319266 -5702 319502 -5466
rect 319586 -5702 319822 -5466
rect 312986 -6342 313222 -6106
rect 313306 -6342 313542 -6106
rect 312986 -6662 313222 -6426
rect 313306 -6662 313542 -6426
rect 325546 46718 325782 46954
rect 325866 46718 326102 46954
rect 325546 26718 325782 26954
rect 325866 26718 326102 26954
rect 325546 6718 325782 6954
rect 325866 6718 326102 6954
rect 325546 -2502 325782 -2266
rect 325866 -2502 326102 -2266
rect 325546 -2822 325782 -2586
rect 325866 -2822 326102 -2586
rect 329266 50378 329502 50614
rect 329586 50378 329822 50614
rect 329266 30378 329502 30614
rect 329586 30378 329822 30614
rect 329266 10378 329502 10614
rect 329586 10378 329822 10614
rect 331826 53058 332062 53294
rect 332146 53058 332382 53294
rect 331826 33058 332062 33294
rect 332146 33058 332382 33294
rect 331826 13058 332062 13294
rect 332146 13058 332382 13294
rect 331826 -1542 332062 -1306
rect 332146 -1542 332382 -1306
rect 331826 -1862 332062 -1626
rect 332146 -1862 332382 -1626
rect 332986 54038 333222 54274
rect 333306 54038 333542 54274
rect 332986 34038 333222 34274
rect 333306 34038 333542 34274
rect 332986 14038 333222 14274
rect 333306 14038 333542 14274
rect 329266 -4422 329502 -4186
rect 329586 -4422 329822 -4186
rect 329266 -4742 329502 -4506
rect 329586 -4742 329822 -4506
rect 322986 -7302 323222 -7066
rect 323306 -7302 323542 -7066
rect 322986 -7622 323222 -7386
rect 323306 -7622 323542 -7386
rect 335546 56718 335782 56954
rect 335866 56718 336102 56954
rect 335546 36718 335782 36954
rect 335866 36718 336102 36954
rect 335546 16718 335782 16954
rect 335866 16718 336102 16954
rect 335546 -3462 335782 -3226
rect 335866 -3462 336102 -3226
rect 335546 -3782 335782 -3546
rect 335866 -3782 336102 -3546
rect 339266 40378 339502 40614
rect 339586 40378 339822 40614
rect 339266 20378 339502 20614
rect 339586 20378 339822 20614
rect 341826 43058 342062 43294
rect 342146 43058 342382 43294
rect 341826 23058 342062 23294
rect 342146 23058 342382 23294
rect 341826 3058 342062 3294
rect 342146 3058 342382 3294
rect 341826 -582 342062 -346
rect 342146 -582 342382 -346
rect 341826 -902 342062 -666
rect 342146 -902 342382 -666
rect 342986 44038 343222 44274
rect 343306 44038 343542 44274
rect 342986 24038 343222 24274
rect 343306 24038 343542 24274
rect 339266 -5382 339502 -5146
rect 339586 -5382 339822 -5146
rect 339266 -5702 339502 -5466
rect 339586 -5702 339822 -5466
rect 332986 -6342 333222 -6106
rect 333306 -6342 333542 -6106
rect 332986 -6662 333222 -6426
rect 333306 -6662 333542 -6426
rect 345546 46718 345782 46954
rect 345866 46718 346102 46954
rect 345546 26718 345782 26954
rect 345866 26718 346102 26954
rect 345546 6718 345782 6954
rect 345866 6718 346102 6954
rect 345546 -2502 345782 -2266
rect 345866 -2502 346102 -2266
rect 345546 -2822 345782 -2586
rect 345866 -2822 346102 -2586
rect 349266 50378 349502 50614
rect 349586 50378 349822 50614
rect 349266 30378 349502 30614
rect 349586 30378 349822 30614
rect 349266 10378 349502 10614
rect 349586 10378 349822 10614
rect 351826 53058 352062 53294
rect 352146 53058 352382 53294
rect 351826 33058 352062 33294
rect 352146 33058 352382 33294
rect 351826 13058 352062 13294
rect 352146 13058 352382 13294
rect 351826 -1542 352062 -1306
rect 352146 -1542 352382 -1306
rect 351826 -1862 352062 -1626
rect 352146 -1862 352382 -1626
rect 352986 54038 353222 54274
rect 353306 54038 353542 54274
rect 352986 34038 353222 34274
rect 353306 34038 353542 34274
rect 352986 14038 353222 14274
rect 353306 14038 353542 14274
rect 349266 -4422 349502 -4186
rect 349586 -4422 349822 -4186
rect 349266 -4742 349502 -4506
rect 349586 -4742 349822 -4506
rect 342986 -7302 343222 -7066
rect 343306 -7302 343542 -7066
rect 342986 -7622 343222 -7386
rect 343306 -7622 343542 -7386
rect 355546 56718 355782 56954
rect 355866 56718 356102 56954
rect 355546 36718 355782 36954
rect 355866 36718 356102 36954
rect 355546 16718 355782 16954
rect 355866 16718 356102 16954
rect 355546 -3462 355782 -3226
rect 355866 -3462 356102 -3226
rect 355546 -3782 355782 -3546
rect 355866 -3782 356102 -3546
rect 359266 40378 359502 40614
rect 359586 40378 359822 40614
rect 359266 20378 359502 20614
rect 359586 20378 359822 20614
rect 361826 43058 362062 43294
rect 362146 43058 362382 43294
rect 361826 23058 362062 23294
rect 362146 23058 362382 23294
rect 361826 3058 362062 3294
rect 362146 3058 362382 3294
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 362986 44038 363222 44274
rect 363306 44038 363542 44274
rect 362986 24038 363222 24274
rect 363306 24038 363542 24274
rect 359266 -5382 359502 -5146
rect 359586 -5382 359822 -5146
rect 359266 -5702 359502 -5466
rect 359586 -5702 359822 -5466
rect 352986 -6342 353222 -6106
rect 353306 -6342 353542 -6106
rect 352986 -6662 353222 -6426
rect 353306 -6662 353542 -6426
rect 365546 46718 365782 46954
rect 365866 46718 366102 46954
rect 365546 26718 365782 26954
rect 365866 26718 366102 26954
rect 365546 6718 365782 6954
rect 365866 6718 366102 6954
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 50378 369502 50614
rect 369586 50378 369822 50614
rect 369266 30378 369502 30614
rect 369586 30378 369822 30614
rect 369266 10378 369502 10614
rect 369586 10378 369822 10614
rect 371826 53058 372062 53294
rect 372146 53058 372382 53294
rect 371826 33058 372062 33294
rect 372146 33058 372382 33294
rect 371826 13058 372062 13294
rect 372146 13058 372382 13294
rect 371826 -1542 372062 -1306
rect 372146 -1542 372382 -1306
rect 371826 -1862 372062 -1626
rect 372146 -1862 372382 -1626
rect 372986 54038 373222 54274
rect 373306 54038 373542 54274
rect 372986 34038 373222 34274
rect 373306 34038 373542 34274
rect 372986 14038 373222 14274
rect 373306 14038 373542 14274
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 362986 -7302 363222 -7066
rect 363306 -7302 363542 -7066
rect 362986 -7622 363222 -7386
rect 363306 -7622 363542 -7386
rect 375546 56718 375782 56954
rect 375866 56718 376102 56954
rect 375546 36718 375782 36954
rect 375866 36718 376102 36954
rect 375546 16718 375782 16954
rect 375866 16718 376102 16954
rect 375546 -3462 375782 -3226
rect 375866 -3462 376102 -3226
rect 375546 -3782 375782 -3546
rect 375866 -3782 376102 -3546
rect 379266 40378 379502 40614
rect 379586 40378 379822 40614
rect 379266 20378 379502 20614
rect 379586 20378 379822 20614
rect 381826 43058 382062 43294
rect 382146 43058 382382 43294
rect 381826 23058 382062 23294
rect 382146 23058 382382 23294
rect 381826 3058 382062 3294
rect 382146 3058 382382 3294
rect 381826 -582 382062 -346
rect 382146 -582 382382 -346
rect 381826 -902 382062 -666
rect 382146 -902 382382 -666
rect 382986 44038 383222 44274
rect 383306 44038 383542 44274
rect 382986 24038 383222 24274
rect 383306 24038 383542 24274
rect 379266 -5382 379502 -5146
rect 379586 -5382 379822 -5146
rect 379266 -5702 379502 -5466
rect 379586 -5702 379822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 385546 46718 385782 46954
rect 385866 46718 386102 46954
rect 385546 26718 385782 26954
rect 385866 26718 386102 26954
rect 385546 6718 385782 6954
rect 385866 6718 386102 6954
rect 385546 -2502 385782 -2266
rect 385866 -2502 386102 -2266
rect 385546 -2822 385782 -2586
rect 385866 -2822 386102 -2586
rect 389266 50378 389502 50614
rect 389586 50378 389822 50614
rect 389266 30378 389502 30614
rect 389586 30378 389822 30614
rect 389266 10378 389502 10614
rect 389586 10378 389822 10614
rect 391826 53058 392062 53294
rect 392146 53058 392382 53294
rect 391826 33058 392062 33294
rect 392146 33058 392382 33294
rect 391826 13058 392062 13294
rect 392146 13058 392382 13294
rect 391826 -1542 392062 -1306
rect 392146 -1542 392382 -1306
rect 391826 -1862 392062 -1626
rect 392146 -1862 392382 -1626
rect 392986 54038 393222 54274
rect 393306 54038 393542 54274
rect 392986 34038 393222 34274
rect 393306 34038 393542 34274
rect 392986 14038 393222 14274
rect 393306 14038 393542 14274
rect 389266 -4422 389502 -4186
rect 389586 -4422 389822 -4186
rect 389266 -4742 389502 -4506
rect 389586 -4742 389822 -4506
rect 382986 -7302 383222 -7066
rect 383306 -7302 383542 -7066
rect 382986 -7622 383222 -7386
rect 383306 -7622 383542 -7386
rect 395546 56718 395782 56954
rect 395866 56718 396102 56954
rect 395546 36718 395782 36954
rect 395866 36718 396102 36954
rect 395546 16718 395782 16954
rect 395866 16718 396102 16954
rect 395546 -3462 395782 -3226
rect 395866 -3462 396102 -3226
rect 395546 -3782 395782 -3546
rect 395866 -3782 396102 -3546
rect 399266 40378 399502 40614
rect 399586 40378 399822 40614
rect 399266 20378 399502 20614
rect 399586 20378 399822 20614
rect 401826 43058 402062 43294
rect 402146 43058 402382 43294
rect 401826 23058 402062 23294
rect 402146 23058 402382 23294
rect 401826 3058 402062 3294
rect 402146 3058 402382 3294
rect 401826 -582 402062 -346
rect 402146 -582 402382 -346
rect 401826 -902 402062 -666
rect 402146 -902 402382 -666
rect 402986 44038 403222 44274
rect 403306 44038 403542 44274
rect 402986 24038 403222 24274
rect 403306 24038 403542 24274
rect 399266 -5382 399502 -5146
rect 399586 -5382 399822 -5146
rect 399266 -5702 399502 -5466
rect 399586 -5702 399822 -5466
rect 392986 -6342 393222 -6106
rect 393306 -6342 393542 -6106
rect 392986 -6662 393222 -6426
rect 393306 -6662 393542 -6426
rect 405546 46718 405782 46954
rect 405866 46718 406102 46954
rect 405546 26718 405782 26954
rect 405866 26718 406102 26954
rect 405546 6718 405782 6954
rect 405866 6718 406102 6954
rect 405546 -2502 405782 -2266
rect 405866 -2502 406102 -2266
rect 405546 -2822 405782 -2586
rect 405866 -2822 406102 -2586
rect 409266 50378 409502 50614
rect 409586 50378 409822 50614
rect 409266 30378 409502 30614
rect 409586 30378 409822 30614
rect 409266 10378 409502 10614
rect 409586 10378 409822 10614
rect 411826 53058 412062 53294
rect 412146 53058 412382 53294
rect 411826 33058 412062 33294
rect 412146 33058 412382 33294
rect 411826 13058 412062 13294
rect 412146 13058 412382 13294
rect 411826 -1542 412062 -1306
rect 412146 -1542 412382 -1306
rect 411826 -1862 412062 -1626
rect 412146 -1862 412382 -1626
rect 412986 54038 413222 54274
rect 413306 54038 413542 54274
rect 412986 34038 413222 34274
rect 413306 34038 413542 34274
rect 412986 14038 413222 14274
rect 413306 14038 413542 14274
rect 409266 -4422 409502 -4186
rect 409586 -4422 409822 -4186
rect 409266 -4742 409502 -4506
rect 409586 -4742 409822 -4506
rect 402986 -7302 403222 -7066
rect 403306 -7302 403542 -7066
rect 402986 -7622 403222 -7386
rect 403306 -7622 403542 -7386
rect 415546 56718 415782 56954
rect 415866 56718 416102 56954
rect 415546 36718 415782 36954
rect 415866 36718 416102 36954
rect 415546 16718 415782 16954
rect 415866 16718 416102 16954
rect 415546 -3462 415782 -3226
rect 415866 -3462 416102 -3226
rect 415546 -3782 415782 -3546
rect 415866 -3782 416102 -3546
rect 419266 40378 419502 40614
rect 419586 40378 419822 40614
rect 419266 20378 419502 20614
rect 419586 20378 419822 20614
rect 421826 43058 422062 43294
rect 422146 43058 422382 43294
rect 421826 23058 422062 23294
rect 422146 23058 422382 23294
rect 421826 3058 422062 3294
rect 422146 3058 422382 3294
rect 421826 -582 422062 -346
rect 422146 -582 422382 -346
rect 421826 -902 422062 -666
rect 422146 -902 422382 -666
rect 422986 44038 423222 44274
rect 423306 44038 423542 44274
rect 422986 24038 423222 24274
rect 423306 24038 423542 24274
rect 419266 -5382 419502 -5146
rect 419586 -5382 419822 -5146
rect 419266 -5702 419502 -5466
rect 419586 -5702 419822 -5466
rect 412986 -6342 413222 -6106
rect 413306 -6342 413542 -6106
rect 412986 -6662 413222 -6426
rect 413306 -6662 413542 -6426
rect 425546 46718 425782 46954
rect 425866 46718 426102 46954
rect 425546 26718 425782 26954
rect 425866 26718 426102 26954
rect 425546 6718 425782 6954
rect 425866 6718 426102 6954
rect 425546 -2502 425782 -2266
rect 425866 -2502 426102 -2266
rect 425546 -2822 425782 -2586
rect 425866 -2822 426102 -2586
rect 429266 50378 429502 50614
rect 429586 50378 429822 50614
rect 429266 30378 429502 30614
rect 429586 30378 429822 30614
rect 429266 10378 429502 10614
rect 429586 10378 429822 10614
rect 431826 53058 432062 53294
rect 432146 53058 432382 53294
rect 431826 33058 432062 33294
rect 432146 33058 432382 33294
rect 431826 13058 432062 13294
rect 432146 13058 432382 13294
rect 431826 -1542 432062 -1306
rect 432146 -1542 432382 -1306
rect 431826 -1862 432062 -1626
rect 432146 -1862 432382 -1626
rect 432986 54038 433222 54274
rect 433306 54038 433542 54274
rect 432986 34038 433222 34274
rect 433306 34038 433542 34274
rect 432986 14038 433222 14274
rect 433306 14038 433542 14274
rect 429266 -4422 429502 -4186
rect 429586 -4422 429822 -4186
rect 429266 -4742 429502 -4506
rect 429586 -4742 429822 -4506
rect 422986 -7302 423222 -7066
rect 423306 -7302 423542 -7066
rect 422986 -7622 423222 -7386
rect 423306 -7622 423542 -7386
rect 435546 56718 435782 56954
rect 435866 56718 436102 56954
rect 435546 36718 435782 36954
rect 435866 36718 436102 36954
rect 435546 16718 435782 16954
rect 435866 16718 436102 16954
rect 435546 -3462 435782 -3226
rect 435866 -3462 436102 -3226
rect 435546 -3782 435782 -3546
rect 435866 -3782 436102 -3546
rect 439266 40378 439502 40614
rect 439586 40378 439822 40614
rect 439266 20378 439502 20614
rect 439586 20378 439822 20614
rect 441826 43058 442062 43294
rect 442146 43058 442382 43294
rect 441826 23058 442062 23294
rect 442146 23058 442382 23294
rect 441826 3058 442062 3294
rect 442146 3058 442382 3294
rect 441826 -582 442062 -346
rect 442146 -582 442382 -346
rect 441826 -902 442062 -666
rect 442146 -902 442382 -666
rect 442986 44038 443222 44274
rect 443306 44038 443542 44274
rect 442986 24038 443222 24274
rect 443306 24038 443542 24274
rect 439266 -5382 439502 -5146
rect 439586 -5382 439822 -5146
rect 439266 -5702 439502 -5466
rect 439586 -5702 439822 -5466
rect 432986 -6342 433222 -6106
rect 433306 -6342 433542 -6106
rect 432986 -6662 433222 -6426
rect 433306 -6662 433542 -6426
rect 445546 46718 445782 46954
rect 445866 46718 446102 46954
rect 445546 26718 445782 26954
rect 445866 26718 446102 26954
rect 445546 6718 445782 6954
rect 445866 6718 446102 6954
rect 445546 -2502 445782 -2266
rect 445866 -2502 446102 -2266
rect 445546 -2822 445782 -2586
rect 445866 -2822 446102 -2586
rect 449266 50378 449502 50614
rect 449586 50378 449822 50614
rect 449266 30378 449502 30614
rect 449586 30378 449822 30614
rect 449266 10378 449502 10614
rect 449586 10378 449822 10614
rect 451826 53058 452062 53294
rect 452146 53058 452382 53294
rect 451826 33058 452062 33294
rect 452146 33058 452382 33294
rect 451826 13058 452062 13294
rect 452146 13058 452382 13294
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 452986 54038 453222 54274
rect 453306 54038 453542 54274
rect 452986 34038 453222 34274
rect 453306 34038 453542 34274
rect 452986 14038 453222 14274
rect 453306 14038 453542 14274
rect 449266 -4422 449502 -4186
rect 449586 -4422 449822 -4186
rect 449266 -4742 449502 -4506
rect 449586 -4742 449822 -4506
rect 442986 -7302 443222 -7066
rect 443306 -7302 443542 -7066
rect 442986 -7622 443222 -7386
rect 443306 -7622 443542 -7386
rect 455546 56718 455782 56954
rect 455866 56718 456102 56954
rect 455546 36718 455782 36954
rect 455866 36718 456102 36954
rect 455546 16718 455782 16954
rect 455866 16718 456102 16954
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 40378 459502 40614
rect 459586 40378 459822 40614
rect 459266 20378 459502 20614
rect 459586 20378 459822 20614
rect 461826 43058 462062 43294
rect 462146 43058 462382 43294
rect 461826 23058 462062 23294
rect 462146 23058 462382 23294
rect 461826 3058 462062 3294
rect 462146 3058 462382 3294
rect 461826 -582 462062 -346
rect 462146 -582 462382 -346
rect 461826 -902 462062 -666
rect 462146 -902 462382 -666
rect 462986 44038 463222 44274
rect 463306 44038 463542 44274
rect 462986 24038 463222 24274
rect 463306 24038 463542 24274
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 452986 -6342 453222 -6106
rect 453306 -6342 453542 -6106
rect 452986 -6662 453222 -6426
rect 453306 -6662 453542 -6426
rect 465546 46718 465782 46954
rect 465866 46718 466102 46954
rect 465546 26718 465782 26954
rect 465866 26718 466102 26954
rect 465546 6718 465782 6954
rect 465866 6718 466102 6954
rect 465546 -2502 465782 -2266
rect 465866 -2502 466102 -2266
rect 465546 -2822 465782 -2586
rect 465866 -2822 466102 -2586
rect 469266 50378 469502 50614
rect 469586 50378 469822 50614
rect 469266 30378 469502 30614
rect 469586 30378 469822 30614
rect 469266 10378 469502 10614
rect 469586 10378 469822 10614
rect 471826 53058 472062 53294
rect 472146 53058 472382 53294
rect 471826 33058 472062 33294
rect 472146 33058 472382 33294
rect 471826 13058 472062 13294
rect 472146 13058 472382 13294
rect 471826 -1542 472062 -1306
rect 472146 -1542 472382 -1306
rect 471826 -1862 472062 -1626
rect 472146 -1862 472382 -1626
rect 472986 54038 473222 54274
rect 473306 54038 473542 54274
rect 472986 34038 473222 34274
rect 473306 34038 473542 34274
rect 472986 14038 473222 14274
rect 473306 14038 473542 14274
rect 469266 -4422 469502 -4186
rect 469586 -4422 469822 -4186
rect 469266 -4742 469502 -4506
rect 469586 -4742 469822 -4506
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 475546 56718 475782 56954
rect 475866 56718 476102 56954
rect 475546 36718 475782 36954
rect 475866 36718 476102 36954
rect 475546 16718 475782 16954
rect 475866 16718 476102 16954
rect 475546 -3462 475782 -3226
rect 475866 -3462 476102 -3226
rect 475546 -3782 475782 -3546
rect 475866 -3782 476102 -3546
rect 479266 40378 479502 40614
rect 479586 40378 479822 40614
rect 479266 20378 479502 20614
rect 479586 20378 479822 20614
rect 481826 43058 482062 43294
rect 482146 43058 482382 43294
rect 481826 23058 482062 23294
rect 482146 23058 482382 23294
rect 481826 3058 482062 3294
rect 482146 3058 482382 3294
rect 481826 -582 482062 -346
rect 482146 -582 482382 -346
rect 481826 -902 482062 -666
rect 482146 -902 482382 -666
rect 482986 44038 483222 44274
rect 483306 44038 483542 44274
rect 482986 24038 483222 24274
rect 483306 24038 483542 24274
rect 479266 -5382 479502 -5146
rect 479586 -5382 479822 -5146
rect 479266 -5702 479502 -5466
rect 479586 -5702 479822 -5466
rect 472986 -6342 473222 -6106
rect 473306 -6342 473542 -6106
rect 472986 -6662 473222 -6426
rect 473306 -6662 473542 -6426
rect 485546 46718 485782 46954
rect 485866 46718 486102 46954
rect 485546 26718 485782 26954
rect 485866 26718 486102 26954
rect 485546 6718 485782 6954
rect 485866 6718 486102 6954
rect 485546 -2502 485782 -2266
rect 485866 -2502 486102 -2266
rect 485546 -2822 485782 -2586
rect 485866 -2822 486102 -2586
rect 489266 50378 489502 50614
rect 489586 50378 489822 50614
rect 489266 30378 489502 30614
rect 489586 30378 489822 30614
rect 489266 10378 489502 10614
rect 489586 10378 489822 10614
rect 491826 53058 492062 53294
rect 492146 53058 492382 53294
rect 491826 33058 492062 33294
rect 492146 33058 492382 33294
rect 491826 13058 492062 13294
rect 492146 13058 492382 13294
rect 491826 -1542 492062 -1306
rect 492146 -1542 492382 -1306
rect 491826 -1862 492062 -1626
rect 492146 -1862 492382 -1626
rect 492986 54038 493222 54274
rect 493306 54038 493542 54274
rect 492986 34038 493222 34274
rect 493306 34038 493542 34274
rect 492986 14038 493222 14274
rect 493306 14038 493542 14274
rect 489266 -4422 489502 -4186
rect 489586 -4422 489822 -4186
rect 489266 -4742 489502 -4506
rect 489586 -4742 489822 -4506
rect 482986 -7302 483222 -7066
rect 483306 -7302 483542 -7066
rect 482986 -7622 483222 -7386
rect 483306 -7622 483542 -7386
rect 495546 56718 495782 56954
rect 495866 56718 496102 56954
rect 495546 36718 495782 36954
rect 495866 36718 496102 36954
rect 495546 16718 495782 16954
rect 495866 16718 496102 16954
rect 495546 -3462 495782 -3226
rect 495866 -3462 496102 -3226
rect 495546 -3782 495782 -3546
rect 495866 -3782 496102 -3546
rect 499266 40378 499502 40614
rect 499586 40378 499822 40614
rect 499266 20378 499502 20614
rect 499586 20378 499822 20614
rect 501826 43058 502062 43294
rect 502146 43058 502382 43294
rect 501826 23058 502062 23294
rect 502146 23058 502382 23294
rect 501826 3058 502062 3294
rect 502146 3058 502382 3294
rect 501826 -582 502062 -346
rect 502146 -582 502382 -346
rect 501826 -902 502062 -666
rect 502146 -902 502382 -666
rect 502986 44038 503222 44274
rect 503306 44038 503542 44274
rect 502986 24038 503222 24274
rect 503306 24038 503542 24274
rect 499266 -5382 499502 -5146
rect 499586 -5382 499822 -5146
rect 499266 -5702 499502 -5466
rect 499586 -5702 499822 -5466
rect 492986 -6342 493222 -6106
rect 493306 -6342 493542 -6106
rect 492986 -6662 493222 -6426
rect 493306 -6662 493542 -6426
rect 505546 46718 505782 46954
rect 505866 46718 506102 46954
rect 505546 26718 505782 26954
rect 505866 26718 506102 26954
rect 505546 6718 505782 6954
rect 505866 6718 506102 6954
rect 505546 -2502 505782 -2266
rect 505866 -2502 506102 -2266
rect 505546 -2822 505782 -2586
rect 505866 -2822 506102 -2586
rect 509266 50378 509502 50614
rect 509586 50378 509822 50614
rect 509266 30378 509502 30614
rect 509586 30378 509822 30614
rect 509266 10378 509502 10614
rect 509586 10378 509822 10614
rect 511826 53058 512062 53294
rect 512146 53058 512382 53294
rect 511826 33058 512062 33294
rect 512146 33058 512382 33294
rect 511826 13058 512062 13294
rect 512146 13058 512382 13294
rect 511826 -1542 512062 -1306
rect 512146 -1542 512382 -1306
rect 511826 -1862 512062 -1626
rect 512146 -1862 512382 -1626
rect 512986 54038 513222 54274
rect 513306 54038 513542 54274
rect 512986 34038 513222 34274
rect 513306 34038 513542 34274
rect 512986 14038 513222 14274
rect 513306 14038 513542 14274
rect 509266 -4422 509502 -4186
rect 509586 -4422 509822 -4186
rect 509266 -4742 509502 -4506
rect 509586 -4742 509822 -4506
rect 502986 -7302 503222 -7066
rect 503306 -7302 503542 -7066
rect 502986 -7622 503222 -7386
rect 503306 -7622 503542 -7386
rect 515546 56718 515782 56954
rect 515866 56718 516102 56954
rect 515546 36718 515782 36954
rect 515866 36718 516102 36954
rect 515546 16718 515782 16954
rect 515866 16718 516102 16954
rect 515546 -3462 515782 -3226
rect 515866 -3462 516102 -3226
rect 515546 -3782 515782 -3546
rect 515866 -3782 516102 -3546
rect 519266 40378 519502 40614
rect 519586 40378 519822 40614
rect 519266 20378 519502 20614
rect 519586 20378 519822 20614
rect 521826 43058 522062 43294
rect 522146 43058 522382 43294
rect 521826 23058 522062 23294
rect 522146 23058 522382 23294
rect 521826 3058 522062 3294
rect 522146 3058 522382 3294
rect 521826 -582 522062 -346
rect 522146 -582 522382 -346
rect 521826 -902 522062 -666
rect 522146 -902 522382 -666
rect 522986 44038 523222 44274
rect 523306 44038 523542 44274
rect 522986 24038 523222 24274
rect 523306 24038 523542 24274
rect 519266 -5382 519502 -5146
rect 519586 -5382 519822 -5146
rect 519266 -5702 519502 -5466
rect 519586 -5702 519822 -5466
rect 512986 -6342 513222 -6106
rect 513306 -6342 513542 -6106
rect 512986 -6662 513222 -6426
rect 513306 -6662 513542 -6426
rect 525546 46718 525782 46954
rect 525866 46718 526102 46954
rect 525546 26718 525782 26954
rect 525866 26718 526102 26954
rect 525546 6718 525782 6954
rect 525866 6718 526102 6954
rect 525546 -2502 525782 -2266
rect 525866 -2502 526102 -2266
rect 525546 -2822 525782 -2586
rect 525866 -2822 526102 -2586
rect 529266 50378 529502 50614
rect 529586 50378 529822 50614
rect 529266 30378 529502 30614
rect 529586 30378 529822 30614
rect 529266 10378 529502 10614
rect 529586 10378 529822 10614
rect 531826 53058 532062 53294
rect 532146 53058 532382 53294
rect 531826 33058 532062 33294
rect 532146 33058 532382 33294
rect 531826 13058 532062 13294
rect 532146 13058 532382 13294
rect 531826 -1542 532062 -1306
rect 532146 -1542 532382 -1306
rect 531826 -1862 532062 -1626
rect 532146 -1862 532382 -1626
rect 532986 54038 533222 54274
rect 533306 54038 533542 54274
rect 532986 34038 533222 34274
rect 533306 34038 533542 34274
rect 532986 14038 533222 14274
rect 533306 14038 533542 14274
rect 529266 -4422 529502 -4186
rect 529586 -4422 529822 -4186
rect 529266 -4742 529502 -4506
rect 529586 -4742 529822 -4506
rect 522986 -7302 523222 -7066
rect 523306 -7302 523542 -7066
rect 522986 -7622 523222 -7386
rect 523306 -7622 523542 -7386
rect 535546 56718 535782 56954
rect 535866 56718 536102 56954
rect 535546 36718 535782 36954
rect 535866 36718 536102 36954
rect 535546 16718 535782 16954
rect 535866 16718 536102 16954
rect 535546 -3462 535782 -3226
rect 535866 -3462 536102 -3226
rect 535546 -3782 535782 -3546
rect 535866 -3782 536102 -3546
rect 539266 40378 539502 40614
rect 539586 40378 539822 40614
rect 539266 20378 539502 20614
rect 539586 20378 539822 20614
rect 541826 43058 542062 43294
rect 542146 43058 542382 43294
rect 541826 23058 542062 23294
rect 542146 23058 542382 23294
rect 541826 3058 542062 3294
rect 542146 3058 542382 3294
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 542986 44038 543222 44274
rect 543306 44038 543542 44274
rect 542986 24038 543222 24274
rect 543306 24038 543542 24274
rect 539266 -5382 539502 -5146
rect 539586 -5382 539822 -5146
rect 539266 -5702 539502 -5466
rect 539586 -5702 539822 -5466
rect 532986 -6342 533222 -6106
rect 533306 -6342 533542 -6106
rect 532986 -6662 533222 -6426
rect 533306 -6662 533542 -6426
rect 545546 46718 545782 46954
rect 545866 46718 546102 46954
rect 545546 26718 545782 26954
rect 545866 26718 546102 26954
rect 545546 6718 545782 6954
rect 545866 6718 546102 6954
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 50378 549502 50614
rect 549586 50378 549822 50614
rect 549266 30378 549502 30614
rect 549586 30378 549822 30614
rect 549266 10378 549502 10614
rect 549586 10378 549822 10614
rect 551826 53058 552062 53294
rect 552146 53058 552382 53294
rect 551826 33058 552062 33294
rect 552146 33058 552382 33294
rect 551826 13058 552062 13294
rect 552146 13058 552382 13294
rect 551826 -1542 552062 -1306
rect 552146 -1542 552382 -1306
rect 551826 -1862 552062 -1626
rect 552146 -1862 552382 -1626
rect 552986 54038 553222 54274
rect 553306 54038 553542 54274
rect 552986 34038 553222 34274
rect 553306 34038 553542 34274
rect 552986 14038 553222 14274
rect 553306 14038 553542 14274
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 542986 -7302 543222 -7066
rect 543306 -7302 543542 -7066
rect 542986 -7622 543222 -7386
rect 543306 -7622 543542 -7386
rect 555546 56718 555782 56954
rect 555866 56718 556102 56954
rect 555546 36718 555782 36954
rect 555866 36718 556102 36954
rect 555546 16718 555782 16954
rect 555866 16718 556102 16954
rect 555546 -3462 555782 -3226
rect 555866 -3462 556102 -3226
rect 555546 -3782 555782 -3546
rect 555866 -3782 556102 -3546
rect 559266 40378 559502 40614
rect 559586 40378 559822 40614
rect 559266 20378 559502 20614
rect 559586 20378 559822 20614
rect 561826 704602 562062 704838
rect 562146 704602 562382 704838
rect 561826 704282 562062 704518
rect 562146 704282 562382 704518
rect 561826 683058 562062 683294
rect 562146 683058 562382 683294
rect 561826 663058 562062 663294
rect 562146 663058 562382 663294
rect 561826 643058 562062 643294
rect 562146 643058 562382 643294
rect 561826 623058 562062 623294
rect 562146 623058 562382 623294
rect 561826 603058 562062 603294
rect 562146 603058 562382 603294
rect 561826 583058 562062 583294
rect 562146 583058 562382 583294
rect 561826 563058 562062 563294
rect 562146 563058 562382 563294
rect 561826 543058 562062 543294
rect 562146 543058 562382 543294
rect 561826 523058 562062 523294
rect 562146 523058 562382 523294
rect 561826 503058 562062 503294
rect 562146 503058 562382 503294
rect 561826 483058 562062 483294
rect 562146 483058 562382 483294
rect 561826 463058 562062 463294
rect 562146 463058 562382 463294
rect 561826 443058 562062 443294
rect 562146 443058 562382 443294
rect 561826 423058 562062 423294
rect 562146 423058 562382 423294
rect 561826 403058 562062 403294
rect 562146 403058 562382 403294
rect 561826 383058 562062 383294
rect 562146 383058 562382 383294
rect 561826 363058 562062 363294
rect 562146 363058 562382 363294
rect 561826 343058 562062 343294
rect 562146 343058 562382 343294
rect 561826 323058 562062 323294
rect 562146 323058 562382 323294
rect 561826 303058 562062 303294
rect 562146 303058 562382 303294
rect 561826 283058 562062 283294
rect 562146 283058 562382 283294
rect 561826 263058 562062 263294
rect 562146 263058 562382 263294
rect 561826 243058 562062 243294
rect 562146 243058 562382 243294
rect 561826 223058 562062 223294
rect 562146 223058 562382 223294
rect 561826 203058 562062 203294
rect 562146 203058 562382 203294
rect 561826 183058 562062 183294
rect 562146 183058 562382 183294
rect 561826 163058 562062 163294
rect 562146 163058 562382 163294
rect 561826 143058 562062 143294
rect 562146 143058 562382 143294
rect 561826 123058 562062 123294
rect 562146 123058 562382 123294
rect 561826 103058 562062 103294
rect 562146 103058 562382 103294
rect 561826 83058 562062 83294
rect 562146 83058 562382 83294
rect 561826 63058 562062 63294
rect 562146 63058 562382 63294
rect 561826 43058 562062 43294
rect 562146 43058 562382 43294
rect 561826 23058 562062 23294
rect 562146 23058 562382 23294
rect 561826 3058 562062 3294
rect 562146 3058 562382 3294
rect 561826 -582 562062 -346
rect 562146 -582 562382 -346
rect 561826 -902 562062 -666
rect 562146 -902 562382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 572986 710362 573222 710598
rect 573306 710362 573542 710598
rect 572986 710042 573222 710278
rect 573306 710042 573542 710278
rect 569266 708442 569502 708678
rect 569586 708442 569822 708678
rect 569266 708122 569502 708358
rect 569586 708122 569822 708358
rect 562986 684038 563222 684274
rect 563306 684038 563542 684274
rect 562986 664038 563222 664274
rect 563306 664038 563542 664274
rect 562986 644038 563222 644274
rect 563306 644038 563542 644274
rect 562986 624038 563222 624274
rect 563306 624038 563542 624274
rect 562986 604038 563222 604274
rect 563306 604038 563542 604274
rect 562986 584038 563222 584274
rect 563306 584038 563542 584274
rect 562986 564038 563222 564274
rect 563306 564038 563542 564274
rect 562986 544038 563222 544274
rect 563306 544038 563542 544274
rect 562986 524038 563222 524274
rect 563306 524038 563542 524274
rect 562986 504038 563222 504274
rect 563306 504038 563542 504274
rect 562986 484038 563222 484274
rect 563306 484038 563542 484274
rect 562986 464038 563222 464274
rect 563306 464038 563542 464274
rect 562986 444038 563222 444274
rect 563306 444038 563542 444274
rect 562986 424038 563222 424274
rect 563306 424038 563542 424274
rect 562986 404038 563222 404274
rect 563306 404038 563542 404274
rect 562986 384038 563222 384274
rect 563306 384038 563542 384274
rect 562986 364038 563222 364274
rect 563306 364038 563542 364274
rect 562986 344038 563222 344274
rect 563306 344038 563542 344274
rect 562986 324038 563222 324274
rect 563306 324038 563542 324274
rect 562986 304038 563222 304274
rect 563306 304038 563542 304274
rect 562986 284038 563222 284274
rect 563306 284038 563542 284274
rect 562986 264038 563222 264274
rect 563306 264038 563542 264274
rect 562986 244038 563222 244274
rect 563306 244038 563542 244274
rect 562986 224038 563222 224274
rect 563306 224038 563542 224274
rect 562986 204038 563222 204274
rect 563306 204038 563542 204274
rect 562986 184038 563222 184274
rect 563306 184038 563542 184274
rect 562986 164038 563222 164274
rect 563306 164038 563542 164274
rect 562986 144038 563222 144274
rect 563306 144038 563542 144274
rect 562986 124038 563222 124274
rect 563306 124038 563542 124274
rect 562986 104038 563222 104274
rect 563306 104038 563542 104274
rect 562986 84038 563222 84274
rect 563306 84038 563542 84274
rect 562986 64038 563222 64274
rect 563306 64038 563542 64274
rect 562986 44038 563222 44274
rect 563306 44038 563542 44274
rect 562986 24038 563222 24274
rect 563306 24038 563542 24274
rect 559266 -5382 559502 -5146
rect 559586 -5382 559822 -5146
rect 559266 -5702 559502 -5466
rect 559586 -5702 559822 -5466
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 565546 706522 565782 706758
rect 565866 706522 566102 706758
rect 565546 706202 565782 706438
rect 565866 706202 566102 706438
rect 565546 686718 565782 686954
rect 565866 686718 566102 686954
rect 565546 666718 565782 666954
rect 565866 666718 566102 666954
rect 565546 646718 565782 646954
rect 565866 646718 566102 646954
rect 565546 626718 565782 626954
rect 565866 626718 566102 626954
rect 565546 606718 565782 606954
rect 565866 606718 566102 606954
rect 565546 586718 565782 586954
rect 565866 586718 566102 586954
rect 565546 566718 565782 566954
rect 565866 566718 566102 566954
rect 565546 546718 565782 546954
rect 565866 546718 566102 546954
rect 565546 526718 565782 526954
rect 565866 526718 566102 526954
rect 565546 506718 565782 506954
rect 565866 506718 566102 506954
rect 565546 486718 565782 486954
rect 565866 486718 566102 486954
rect 565546 466718 565782 466954
rect 565866 466718 566102 466954
rect 565546 446718 565782 446954
rect 565866 446718 566102 446954
rect 565546 426718 565782 426954
rect 565866 426718 566102 426954
rect 565546 406718 565782 406954
rect 565866 406718 566102 406954
rect 565546 386718 565782 386954
rect 565866 386718 566102 386954
rect 565546 366718 565782 366954
rect 565866 366718 566102 366954
rect 565546 346718 565782 346954
rect 565866 346718 566102 346954
rect 565546 326718 565782 326954
rect 565866 326718 566102 326954
rect 565546 306718 565782 306954
rect 565866 306718 566102 306954
rect 565546 286718 565782 286954
rect 565866 286718 566102 286954
rect 565546 266718 565782 266954
rect 565866 266718 566102 266954
rect 565546 246718 565782 246954
rect 565866 246718 566102 246954
rect 565546 226718 565782 226954
rect 565866 226718 566102 226954
rect 565546 206718 565782 206954
rect 565866 206718 566102 206954
rect 565546 186718 565782 186954
rect 565866 186718 566102 186954
rect 565546 166718 565782 166954
rect 565866 166718 566102 166954
rect 565546 146718 565782 146954
rect 565866 146718 566102 146954
rect 565546 126718 565782 126954
rect 565866 126718 566102 126954
rect 565546 106718 565782 106954
rect 565866 106718 566102 106954
rect 565546 86718 565782 86954
rect 565866 86718 566102 86954
rect 565546 66718 565782 66954
rect 565866 66718 566102 66954
rect 565546 46718 565782 46954
rect 565866 46718 566102 46954
rect 565546 26718 565782 26954
rect 565866 26718 566102 26954
rect 565546 6718 565782 6954
rect 565866 6718 566102 6954
rect 565546 -2502 565782 -2266
rect 565866 -2502 566102 -2266
rect 565546 -2822 565782 -2586
rect 565866 -2822 566102 -2586
rect 569266 690378 569502 690614
rect 569586 690378 569822 690614
rect 569266 670378 569502 670614
rect 569586 670378 569822 670614
rect 569266 650378 569502 650614
rect 569586 650378 569822 650614
rect 569266 630378 569502 630614
rect 569586 630378 569822 630614
rect 569266 610378 569502 610614
rect 569586 610378 569822 610614
rect 569266 590378 569502 590614
rect 569586 590378 569822 590614
rect 569266 570378 569502 570614
rect 569586 570378 569822 570614
rect 569266 550378 569502 550614
rect 569586 550378 569822 550614
rect 569266 530378 569502 530614
rect 569586 530378 569822 530614
rect 569266 510378 569502 510614
rect 569586 510378 569822 510614
rect 569266 490378 569502 490614
rect 569586 490378 569822 490614
rect 569266 470378 569502 470614
rect 569586 470378 569822 470614
rect 569266 450378 569502 450614
rect 569586 450378 569822 450614
rect 569266 430378 569502 430614
rect 569586 430378 569822 430614
rect 569266 410378 569502 410614
rect 569586 410378 569822 410614
rect 569266 390378 569502 390614
rect 569586 390378 569822 390614
rect 569266 370378 569502 370614
rect 569586 370378 569822 370614
rect 569266 350378 569502 350614
rect 569586 350378 569822 350614
rect 569266 330378 569502 330614
rect 569586 330378 569822 330614
rect 569266 310378 569502 310614
rect 569586 310378 569822 310614
rect 569266 290378 569502 290614
rect 569586 290378 569822 290614
rect 569266 270378 569502 270614
rect 569586 270378 569822 270614
rect 569266 250378 569502 250614
rect 569586 250378 569822 250614
rect 569266 230378 569502 230614
rect 569586 230378 569822 230614
rect 569266 210378 569502 210614
rect 569586 210378 569822 210614
rect 569266 190378 569502 190614
rect 569586 190378 569822 190614
rect 569266 170378 569502 170614
rect 569586 170378 569822 170614
rect 569266 150378 569502 150614
rect 569586 150378 569822 150614
rect 569266 130378 569502 130614
rect 569586 130378 569822 130614
rect 569266 110378 569502 110614
rect 569586 110378 569822 110614
rect 569266 90378 569502 90614
rect 569586 90378 569822 90614
rect 569266 70378 569502 70614
rect 569586 70378 569822 70614
rect 569266 50378 569502 50614
rect 569586 50378 569822 50614
rect 569266 30378 569502 30614
rect 569586 30378 569822 30614
rect 569266 10378 569502 10614
rect 569586 10378 569822 10614
rect 571826 705562 572062 705798
rect 572146 705562 572382 705798
rect 571826 705242 572062 705478
rect 572146 705242 572382 705478
rect 571826 693058 572062 693294
rect 572146 693058 572382 693294
rect 571826 673058 572062 673294
rect 572146 673058 572382 673294
rect 571826 653058 572062 653294
rect 572146 653058 572382 653294
rect 571826 633058 572062 633294
rect 572146 633058 572382 633294
rect 571826 613058 572062 613294
rect 572146 613058 572382 613294
rect 571826 593058 572062 593294
rect 572146 593058 572382 593294
rect 571826 573058 572062 573294
rect 572146 573058 572382 573294
rect 571826 553058 572062 553294
rect 572146 553058 572382 553294
rect 571826 533058 572062 533294
rect 572146 533058 572382 533294
rect 571826 513058 572062 513294
rect 572146 513058 572382 513294
rect 571826 493058 572062 493294
rect 572146 493058 572382 493294
rect 571826 473058 572062 473294
rect 572146 473058 572382 473294
rect 571826 453058 572062 453294
rect 572146 453058 572382 453294
rect 571826 433058 572062 433294
rect 572146 433058 572382 433294
rect 571826 413058 572062 413294
rect 572146 413058 572382 413294
rect 571826 393058 572062 393294
rect 572146 393058 572382 393294
rect 571826 373058 572062 373294
rect 572146 373058 572382 373294
rect 571826 353058 572062 353294
rect 572146 353058 572382 353294
rect 571826 333058 572062 333294
rect 572146 333058 572382 333294
rect 571826 313058 572062 313294
rect 572146 313058 572382 313294
rect 571826 293058 572062 293294
rect 572146 293058 572382 293294
rect 571826 273058 572062 273294
rect 572146 273058 572382 273294
rect 571826 253058 572062 253294
rect 572146 253058 572382 253294
rect 571826 233058 572062 233294
rect 572146 233058 572382 233294
rect 571826 213058 572062 213294
rect 572146 213058 572382 213294
rect 571826 193058 572062 193294
rect 572146 193058 572382 193294
rect 571826 173058 572062 173294
rect 572146 173058 572382 173294
rect 571826 153058 572062 153294
rect 572146 153058 572382 153294
rect 571826 133058 572062 133294
rect 572146 133058 572382 133294
rect 571826 113058 572062 113294
rect 572146 113058 572382 113294
rect 571826 93058 572062 93294
rect 572146 93058 572382 93294
rect 571826 73058 572062 73294
rect 572146 73058 572382 73294
rect 571826 53058 572062 53294
rect 572146 53058 572382 53294
rect 571826 33058 572062 33294
rect 572146 33058 572382 33294
rect 571826 13058 572062 13294
rect 572146 13058 572382 13294
rect 571826 -1542 572062 -1306
rect 572146 -1542 572382 -1306
rect 571826 -1862 572062 -1626
rect 572146 -1862 572382 -1626
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 579266 709402 579502 709638
rect 579586 709402 579822 709638
rect 579266 709082 579502 709318
rect 579586 709082 579822 709318
rect 572986 694038 573222 694274
rect 573306 694038 573542 694274
rect 572986 674038 573222 674274
rect 573306 674038 573542 674274
rect 572986 654038 573222 654274
rect 573306 654038 573542 654274
rect 572986 634038 573222 634274
rect 573306 634038 573542 634274
rect 572986 614038 573222 614274
rect 573306 614038 573542 614274
rect 572986 594038 573222 594274
rect 573306 594038 573542 594274
rect 572986 574038 573222 574274
rect 573306 574038 573542 574274
rect 572986 554038 573222 554274
rect 573306 554038 573542 554274
rect 572986 534038 573222 534274
rect 573306 534038 573542 534274
rect 572986 514038 573222 514274
rect 573306 514038 573542 514274
rect 572986 494038 573222 494274
rect 573306 494038 573542 494274
rect 572986 474038 573222 474274
rect 573306 474038 573542 474274
rect 572986 454038 573222 454274
rect 573306 454038 573542 454274
rect 572986 434038 573222 434274
rect 573306 434038 573542 434274
rect 572986 414038 573222 414274
rect 573306 414038 573542 414274
rect 572986 394038 573222 394274
rect 573306 394038 573542 394274
rect 572986 374038 573222 374274
rect 573306 374038 573542 374274
rect 572986 354038 573222 354274
rect 573306 354038 573542 354274
rect 572986 334038 573222 334274
rect 573306 334038 573542 334274
rect 572986 314038 573222 314274
rect 573306 314038 573542 314274
rect 572986 294038 573222 294274
rect 573306 294038 573542 294274
rect 572986 274038 573222 274274
rect 573306 274038 573542 274274
rect 572986 254038 573222 254274
rect 573306 254038 573542 254274
rect 572986 234038 573222 234274
rect 573306 234038 573542 234274
rect 572986 214038 573222 214274
rect 573306 214038 573542 214274
rect 572986 194038 573222 194274
rect 573306 194038 573542 194274
rect 572986 174038 573222 174274
rect 573306 174038 573542 174274
rect 572986 154038 573222 154274
rect 573306 154038 573542 154274
rect 572986 134038 573222 134274
rect 573306 134038 573542 134274
rect 572986 114038 573222 114274
rect 573306 114038 573542 114274
rect 572986 94038 573222 94274
rect 573306 94038 573542 94274
rect 572986 74038 573222 74274
rect 573306 74038 573542 74274
rect 572986 54038 573222 54274
rect 573306 54038 573542 54274
rect 572986 34038 573222 34274
rect 573306 34038 573542 34274
rect 572986 14038 573222 14274
rect 573306 14038 573542 14274
rect 569266 -4422 569502 -4186
rect 569586 -4422 569822 -4186
rect 569266 -4742 569502 -4506
rect 569586 -4742 569822 -4506
rect 562986 -7302 563222 -7066
rect 563306 -7302 563542 -7066
rect 562986 -7622 563222 -7386
rect 563306 -7622 563542 -7386
rect 575546 707482 575782 707718
rect 575866 707482 576102 707718
rect 575546 707162 575782 707398
rect 575866 707162 576102 707398
rect 575546 696718 575782 696954
rect 575866 696718 576102 696954
rect 575546 676718 575782 676954
rect 575866 676718 576102 676954
rect 575546 656718 575782 656954
rect 575866 656718 576102 656954
rect 575546 636718 575782 636954
rect 575866 636718 576102 636954
rect 575546 616718 575782 616954
rect 575866 616718 576102 616954
rect 575546 596718 575782 596954
rect 575866 596718 576102 596954
rect 575546 576718 575782 576954
rect 575866 576718 576102 576954
rect 575546 556718 575782 556954
rect 575866 556718 576102 556954
rect 575546 536718 575782 536954
rect 575866 536718 576102 536954
rect 575546 516718 575782 516954
rect 575866 516718 576102 516954
rect 575546 496718 575782 496954
rect 575866 496718 576102 496954
rect 575546 476718 575782 476954
rect 575866 476718 576102 476954
rect 575546 456718 575782 456954
rect 575866 456718 576102 456954
rect 575546 436718 575782 436954
rect 575866 436718 576102 436954
rect 575546 416718 575782 416954
rect 575866 416718 576102 416954
rect 575546 396718 575782 396954
rect 575866 396718 576102 396954
rect 575546 376718 575782 376954
rect 575866 376718 576102 376954
rect 575546 356718 575782 356954
rect 575866 356718 576102 356954
rect 575546 336718 575782 336954
rect 575866 336718 576102 336954
rect 575546 316718 575782 316954
rect 575866 316718 576102 316954
rect 575546 296718 575782 296954
rect 575866 296718 576102 296954
rect 575546 276718 575782 276954
rect 575866 276718 576102 276954
rect 575546 256718 575782 256954
rect 575866 256718 576102 256954
rect 575546 236718 575782 236954
rect 575866 236718 576102 236954
rect 575546 216718 575782 216954
rect 575866 216718 576102 216954
rect 575546 196718 575782 196954
rect 575866 196718 576102 196954
rect 575546 176718 575782 176954
rect 575866 176718 576102 176954
rect 575546 156718 575782 156954
rect 575866 156718 576102 156954
rect 575546 136718 575782 136954
rect 575866 136718 576102 136954
rect 575546 116718 575782 116954
rect 575866 116718 576102 116954
rect 575546 96718 575782 96954
rect 575866 96718 576102 96954
rect 575546 76718 575782 76954
rect 575866 76718 576102 76954
rect 575546 56718 575782 56954
rect 575866 56718 576102 56954
rect 575546 36718 575782 36954
rect 575866 36718 576102 36954
rect 575546 16718 575782 16954
rect 575866 16718 576102 16954
rect 575546 -3462 575782 -3226
rect 575866 -3462 576102 -3226
rect 575546 -3782 575782 -3546
rect 575866 -3782 576102 -3546
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 579266 700378 579502 700614
rect 579586 700378 579822 700614
rect 579266 680378 579502 680614
rect 579586 680378 579822 680614
rect 579266 660378 579502 660614
rect 579586 660378 579822 660614
rect 579266 640378 579502 640614
rect 579586 640378 579822 640614
rect 579266 620378 579502 620614
rect 579586 620378 579822 620614
rect 579266 600378 579502 600614
rect 579586 600378 579822 600614
rect 579266 580378 579502 580614
rect 579586 580378 579822 580614
rect 579266 560378 579502 560614
rect 579586 560378 579822 560614
rect 579266 540378 579502 540614
rect 579586 540378 579822 540614
rect 579266 520378 579502 520614
rect 579586 520378 579822 520614
rect 579266 500378 579502 500614
rect 579586 500378 579822 500614
rect 579266 480378 579502 480614
rect 579586 480378 579822 480614
rect 579266 460378 579502 460614
rect 579586 460378 579822 460614
rect 579266 440378 579502 440614
rect 579586 440378 579822 440614
rect 579266 420378 579502 420614
rect 579586 420378 579822 420614
rect 579266 400378 579502 400614
rect 579586 400378 579822 400614
rect 579266 380378 579502 380614
rect 579586 380378 579822 380614
rect 579266 360378 579502 360614
rect 579586 360378 579822 360614
rect 579266 340378 579502 340614
rect 579586 340378 579822 340614
rect 579266 320378 579502 320614
rect 579586 320378 579822 320614
rect 579266 300378 579502 300614
rect 579586 300378 579822 300614
rect 579266 280378 579502 280614
rect 579586 280378 579822 280614
rect 579266 260378 579502 260614
rect 579586 260378 579822 260614
rect 579266 240378 579502 240614
rect 579586 240378 579822 240614
rect 579266 220378 579502 220614
rect 579586 220378 579822 220614
rect 579266 200378 579502 200614
rect 579586 200378 579822 200614
rect 579266 180378 579502 180614
rect 579586 180378 579822 180614
rect 579266 160378 579502 160614
rect 579586 160378 579822 160614
rect 579266 140378 579502 140614
rect 579586 140378 579822 140614
rect 579266 120378 579502 120614
rect 579586 120378 579822 120614
rect 579266 100378 579502 100614
rect 579586 100378 579822 100614
rect 579266 80378 579502 80614
rect 579586 80378 579822 80614
rect 579266 60378 579502 60614
rect 579586 60378 579822 60614
rect 579266 40378 579502 40614
rect 579586 40378 579822 40614
rect 579266 20378 579502 20614
rect 579586 20378 579822 20614
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581826 704602 582062 704838
rect 582146 704602 582382 704838
rect 581826 704282 582062 704518
rect 582146 704282 582382 704518
rect 581826 683058 582062 683294
rect 582146 683058 582382 683294
rect 581826 663058 582062 663294
rect 582146 663058 582382 663294
rect 581826 643058 582062 643294
rect 582146 643058 582382 643294
rect 581826 623058 582062 623294
rect 582146 623058 582382 623294
rect 581826 603058 582062 603294
rect 582146 603058 582382 603294
rect 581826 583058 582062 583294
rect 582146 583058 582382 583294
rect 581826 563058 582062 563294
rect 582146 563058 582382 563294
rect 581826 543058 582062 543294
rect 582146 543058 582382 543294
rect 581826 523058 582062 523294
rect 582146 523058 582382 523294
rect 581826 503058 582062 503294
rect 582146 503058 582382 503294
rect 581826 483058 582062 483294
rect 582146 483058 582382 483294
rect 581826 463058 582062 463294
rect 582146 463058 582382 463294
rect 581826 443058 582062 443294
rect 582146 443058 582382 443294
rect 581826 423058 582062 423294
rect 582146 423058 582382 423294
rect 581826 403058 582062 403294
rect 582146 403058 582382 403294
rect 581826 383058 582062 383294
rect 582146 383058 582382 383294
rect 581826 363058 582062 363294
rect 582146 363058 582382 363294
rect 581826 343058 582062 343294
rect 582146 343058 582382 343294
rect 581826 323058 582062 323294
rect 582146 323058 582382 323294
rect 581826 303058 582062 303294
rect 582146 303058 582382 303294
rect 581826 283058 582062 283294
rect 582146 283058 582382 283294
rect 581826 263058 582062 263294
rect 582146 263058 582382 263294
rect 581826 243058 582062 243294
rect 582146 243058 582382 243294
rect 581826 223058 582062 223294
rect 582146 223058 582382 223294
rect 581826 203058 582062 203294
rect 582146 203058 582382 203294
rect 581826 183058 582062 183294
rect 582146 183058 582382 183294
rect 581826 163058 582062 163294
rect 582146 163058 582382 163294
rect 581826 143058 582062 143294
rect 582146 143058 582382 143294
rect 581826 123058 582062 123294
rect 582146 123058 582382 123294
rect 581826 103058 582062 103294
rect 582146 103058 582382 103294
rect 581826 83058 582062 83294
rect 582146 83058 582382 83294
rect 581826 63058 582062 63294
rect 582146 63058 582382 63294
rect 581826 43058 582062 43294
rect 582146 43058 582382 43294
rect 581826 23058 582062 23294
rect 582146 23058 582382 23294
rect 581826 3058 582062 3294
rect 582146 3058 582382 3294
rect 581826 -582 582062 -346
rect 582146 -582 582382 -346
rect 581826 -902 582062 -666
rect 582146 -902 582382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 683058 585578 683294
rect 585662 683058 585898 683294
rect 585342 663058 585578 663294
rect 585662 663058 585898 663294
rect 585342 643058 585578 643294
rect 585662 643058 585898 643294
rect 585342 623058 585578 623294
rect 585662 623058 585898 623294
rect 585342 603058 585578 603294
rect 585662 603058 585898 603294
rect 585342 583058 585578 583294
rect 585662 583058 585898 583294
rect 585342 563058 585578 563294
rect 585662 563058 585898 563294
rect 585342 543058 585578 543294
rect 585662 543058 585898 543294
rect 585342 523058 585578 523294
rect 585662 523058 585898 523294
rect 585342 503058 585578 503294
rect 585662 503058 585898 503294
rect 585342 483058 585578 483294
rect 585662 483058 585898 483294
rect 585342 463058 585578 463294
rect 585662 463058 585898 463294
rect 585342 443058 585578 443294
rect 585662 443058 585898 443294
rect 585342 423058 585578 423294
rect 585662 423058 585898 423294
rect 585342 403058 585578 403294
rect 585662 403058 585898 403294
rect 585342 383058 585578 383294
rect 585662 383058 585898 383294
rect 585342 363058 585578 363294
rect 585662 363058 585898 363294
rect 585342 343058 585578 343294
rect 585662 343058 585898 343294
rect 585342 323058 585578 323294
rect 585662 323058 585898 323294
rect 585342 303058 585578 303294
rect 585662 303058 585898 303294
rect 585342 283058 585578 283294
rect 585662 283058 585898 283294
rect 585342 263058 585578 263294
rect 585662 263058 585898 263294
rect 585342 243058 585578 243294
rect 585662 243058 585898 243294
rect 585342 223058 585578 223294
rect 585662 223058 585898 223294
rect 585342 203058 585578 203294
rect 585662 203058 585898 203294
rect 585342 183058 585578 183294
rect 585662 183058 585898 183294
rect 585342 163058 585578 163294
rect 585662 163058 585898 163294
rect 585342 143058 585578 143294
rect 585662 143058 585898 143294
rect 585342 123058 585578 123294
rect 585662 123058 585898 123294
rect 585342 103058 585578 103294
rect 585662 103058 585898 103294
rect 585342 83058 585578 83294
rect 585662 83058 585898 83294
rect 585342 63058 585578 63294
rect 585662 63058 585898 63294
rect 585342 43058 585578 43294
rect 585662 43058 585898 43294
rect 585342 23058 585578 23294
rect 585662 23058 585898 23294
rect 585342 3058 585578 3294
rect 585662 3058 585898 3294
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 693058 586538 693294
rect 586622 693058 586858 693294
rect 586302 673058 586538 673294
rect 586622 673058 586858 673294
rect 586302 653058 586538 653294
rect 586622 653058 586858 653294
rect 586302 633058 586538 633294
rect 586622 633058 586858 633294
rect 586302 613058 586538 613294
rect 586622 613058 586858 613294
rect 586302 593058 586538 593294
rect 586622 593058 586858 593294
rect 586302 573058 586538 573294
rect 586622 573058 586858 573294
rect 586302 553058 586538 553294
rect 586622 553058 586858 553294
rect 586302 533058 586538 533294
rect 586622 533058 586858 533294
rect 586302 513058 586538 513294
rect 586622 513058 586858 513294
rect 586302 493058 586538 493294
rect 586622 493058 586858 493294
rect 586302 473058 586538 473294
rect 586622 473058 586858 473294
rect 586302 453058 586538 453294
rect 586622 453058 586858 453294
rect 586302 433058 586538 433294
rect 586622 433058 586858 433294
rect 586302 413058 586538 413294
rect 586622 413058 586858 413294
rect 586302 393058 586538 393294
rect 586622 393058 586858 393294
rect 586302 373058 586538 373294
rect 586622 373058 586858 373294
rect 586302 353058 586538 353294
rect 586622 353058 586858 353294
rect 586302 333058 586538 333294
rect 586622 333058 586858 333294
rect 586302 313058 586538 313294
rect 586622 313058 586858 313294
rect 586302 293058 586538 293294
rect 586622 293058 586858 293294
rect 586302 273058 586538 273294
rect 586622 273058 586858 273294
rect 586302 253058 586538 253294
rect 586622 253058 586858 253294
rect 586302 233058 586538 233294
rect 586622 233058 586858 233294
rect 586302 213058 586538 213294
rect 586622 213058 586858 213294
rect 586302 193058 586538 193294
rect 586622 193058 586858 193294
rect 586302 173058 586538 173294
rect 586622 173058 586858 173294
rect 586302 153058 586538 153294
rect 586622 153058 586858 153294
rect 586302 133058 586538 133294
rect 586622 133058 586858 133294
rect 586302 113058 586538 113294
rect 586622 113058 586858 113294
rect 586302 93058 586538 93294
rect 586622 93058 586858 93294
rect 586302 73058 586538 73294
rect 586622 73058 586858 73294
rect 586302 53058 586538 53294
rect 586622 53058 586858 53294
rect 586302 33058 586538 33294
rect 586622 33058 586858 33294
rect 586302 13058 586538 13294
rect 586622 13058 586858 13294
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 686718 587498 686954
rect 587582 686718 587818 686954
rect 587262 666718 587498 666954
rect 587582 666718 587818 666954
rect 587262 646718 587498 646954
rect 587582 646718 587818 646954
rect 587262 626718 587498 626954
rect 587582 626718 587818 626954
rect 587262 606718 587498 606954
rect 587582 606718 587818 606954
rect 587262 586718 587498 586954
rect 587582 586718 587818 586954
rect 587262 566718 587498 566954
rect 587582 566718 587818 566954
rect 587262 546718 587498 546954
rect 587582 546718 587818 546954
rect 587262 526718 587498 526954
rect 587582 526718 587818 526954
rect 587262 506718 587498 506954
rect 587582 506718 587818 506954
rect 587262 486718 587498 486954
rect 587582 486718 587818 486954
rect 587262 466718 587498 466954
rect 587582 466718 587818 466954
rect 587262 446718 587498 446954
rect 587582 446718 587818 446954
rect 587262 426718 587498 426954
rect 587582 426718 587818 426954
rect 587262 406718 587498 406954
rect 587582 406718 587818 406954
rect 587262 386718 587498 386954
rect 587582 386718 587818 386954
rect 587262 366718 587498 366954
rect 587582 366718 587818 366954
rect 587262 346718 587498 346954
rect 587582 346718 587818 346954
rect 587262 326718 587498 326954
rect 587582 326718 587818 326954
rect 587262 306718 587498 306954
rect 587582 306718 587818 306954
rect 587262 286718 587498 286954
rect 587582 286718 587818 286954
rect 587262 266718 587498 266954
rect 587582 266718 587818 266954
rect 587262 246718 587498 246954
rect 587582 246718 587818 246954
rect 587262 226718 587498 226954
rect 587582 226718 587818 226954
rect 587262 206718 587498 206954
rect 587582 206718 587818 206954
rect 587262 186718 587498 186954
rect 587582 186718 587818 186954
rect 587262 166718 587498 166954
rect 587582 166718 587818 166954
rect 587262 146718 587498 146954
rect 587582 146718 587818 146954
rect 587262 126718 587498 126954
rect 587582 126718 587818 126954
rect 587262 106718 587498 106954
rect 587582 106718 587818 106954
rect 587262 86718 587498 86954
rect 587582 86718 587818 86954
rect 587262 66718 587498 66954
rect 587582 66718 587818 66954
rect 587262 46718 587498 46954
rect 587582 46718 587818 46954
rect 587262 26718 587498 26954
rect 587582 26718 587818 26954
rect 587262 6718 587498 6954
rect 587582 6718 587818 6954
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 696718 588458 696954
rect 588542 696718 588778 696954
rect 588222 676718 588458 676954
rect 588542 676718 588778 676954
rect 588222 656718 588458 656954
rect 588542 656718 588778 656954
rect 588222 636718 588458 636954
rect 588542 636718 588778 636954
rect 588222 616718 588458 616954
rect 588542 616718 588778 616954
rect 588222 596718 588458 596954
rect 588542 596718 588778 596954
rect 588222 576718 588458 576954
rect 588542 576718 588778 576954
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 536718 588458 536954
rect 588542 536718 588778 536954
rect 588222 516718 588458 516954
rect 588542 516718 588778 516954
rect 588222 496718 588458 496954
rect 588542 496718 588778 496954
rect 588222 476718 588458 476954
rect 588542 476718 588778 476954
rect 588222 456718 588458 456954
rect 588542 456718 588778 456954
rect 588222 436718 588458 436954
rect 588542 436718 588778 436954
rect 588222 416718 588458 416954
rect 588542 416718 588778 416954
rect 588222 396718 588458 396954
rect 588542 396718 588778 396954
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 356718 588458 356954
rect 588542 356718 588778 356954
rect 588222 336718 588458 336954
rect 588542 336718 588778 336954
rect 588222 316718 588458 316954
rect 588542 316718 588778 316954
rect 588222 296718 588458 296954
rect 588542 296718 588778 296954
rect 588222 276718 588458 276954
rect 588542 276718 588778 276954
rect 588222 256718 588458 256954
rect 588542 256718 588778 256954
rect 588222 236718 588458 236954
rect 588542 236718 588778 236954
rect 588222 216718 588458 216954
rect 588542 216718 588778 216954
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 176718 588458 176954
rect 588542 176718 588778 176954
rect 588222 156718 588458 156954
rect 588542 156718 588778 156954
rect 588222 136718 588458 136954
rect 588542 136718 588778 136954
rect 588222 116718 588458 116954
rect 588542 116718 588778 116954
rect 588222 96718 588458 96954
rect 588542 96718 588778 96954
rect 588222 76718 588458 76954
rect 588542 76718 588778 76954
rect 588222 56718 588458 56954
rect 588542 56718 588778 56954
rect 588222 36718 588458 36954
rect 588542 36718 588778 36954
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 690378 589418 690614
rect 589502 690378 589738 690614
rect 589182 670378 589418 670614
rect 589502 670378 589738 670614
rect 589182 650378 589418 650614
rect 589502 650378 589738 650614
rect 589182 630378 589418 630614
rect 589502 630378 589738 630614
rect 589182 610378 589418 610614
rect 589502 610378 589738 610614
rect 589182 590378 589418 590614
rect 589502 590378 589738 590614
rect 589182 570378 589418 570614
rect 589502 570378 589738 570614
rect 589182 550378 589418 550614
rect 589502 550378 589738 550614
rect 589182 530378 589418 530614
rect 589502 530378 589738 530614
rect 589182 510378 589418 510614
rect 589502 510378 589738 510614
rect 589182 490378 589418 490614
rect 589502 490378 589738 490614
rect 589182 470378 589418 470614
rect 589502 470378 589738 470614
rect 589182 450378 589418 450614
rect 589502 450378 589738 450614
rect 589182 430378 589418 430614
rect 589502 430378 589738 430614
rect 589182 410378 589418 410614
rect 589502 410378 589738 410614
rect 589182 390378 589418 390614
rect 589502 390378 589738 390614
rect 589182 370378 589418 370614
rect 589502 370378 589738 370614
rect 589182 350378 589418 350614
rect 589502 350378 589738 350614
rect 589182 330378 589418 330614
rect 589502 330378 589738 330614
rect 589182 310378 589418 310614
rect 589502 310378 589738 310614
rect 589182 290378 589418 290614
rect 589502 290378 589738 290614
rect 589182 270378 589418 270614
rect 589502 270378 589738 270614
rect 589182 250378 589418 250614
rect 589502 250378 589738 250614
rect 589182 230378 589418 230614
rect 589502 230378 589738 230614
rect 589182 210378 589418 210614
rect 589502 210378 589738 210614
rect 589182 190378 589418 190614
rect 589502 190378 589738 190614
rect 589182 170378 589418 170614
rect 589502 170378 589738 170614
rect 589182 150378 589418 150614
rect 589502 150378 589738 150614
rect 589182 130378 589418 130614
rect 589502 130378 589738 130614
rect 589182 110378 589418 110614
rect 589502 110378 589738 110614
rect 589182 90378 589418 90614
rect 589502 90378 589738 90614
rect 589182 70378 589418 70614
rect 589502 70378 589738 70614
rect 589182 50378 589418 50614
rect 589502 50378 589738 50614
rect 589182 30378 589418 30614
rect 589502 30378 589738 30614
rect 589182 10378 589418 10614
rect 589502 10378 589738 10614
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 700378 590378 700614
rect 590462 700378 590698 700614
rect 590142 680378 590378 680614
rect 590462 680378 590698 680614
rect 590142 660378 590378 660614
rect 590462 660378 590698 660614
rect 590142 640378 590378 640614
rect 590462 640378 590698 640614
rect 590142 620378 590378 620614
rect 590462 620378 590698 620614
rect 590142 600378 590378 600614
rect 590462 600378 590698 600614
rect 590142 580378 590378 580614
rect 590462 580378 590698 580614
rect 590142 560378 590378 560614
rect 590462 560378 590698 560614
rect 590142 540378 590378 540614
rect 590462 540378 590698 540614
rect 590142 520378 590378 520614
rect 590462 520378 590698 520614
rect 590142 500378 590378 500614
rect 590462 500378 590698 500614
rect 590142 480378 590378 480614
rect 590462 480378 590698 480614
rect 590142 460378 590378 460614
rect 590462 460378 590698 460614
rect 590142 440378 590378 440614
rect 590462 440378 590698 440614
rect 590142 420378 590378 420614
rect 590462 420378 590698 420614
rect 590142 400378 590378 400614
rect 590462 400378 590698 400614
rect 590142 380378 590378 380614
rect 590462 380378 590698 380614
rect 590142 360378 590378 360614
rect 590462 360378 590698 360614
rect 590142 340378 590378 340614
rect 590462 340378 590698 340614
rect 590142 320378 590378 320614
rect 590462 320378 590698 320614
rect 590142 300378 590378 300614
rect 590462 300378 590698 300614
rect 590142 280378 590378 280614
rect 590462 280378 590698 280614
rect 590142 260378 590378 260614
rect 590462 260378 590698 260614
rect 590142 240378 590378 240614
rect 590462 240378 590698 240614
rect 590142 220378 590378 220614
rect 590462 220378 590698 220614
rect 590142 200378 590378 200614
rect 590462 200378 590698 200614
rect 590142 180378 590378 180614
rect 590462 180378 590698 180614
rect 590142 160378 590378 160614
rect 590462 160378 590698 160614
rect 590142 140378 590378 140614
rect 590462 140378 590698 140614
rect 590142 120378 590378 120614
rect 590462 120378 590698 120614
rect 590142 100378 590378 100614
rect 590462 100378 590698 100614
rect 590142 80378 590378 80614
rect 590462 80378 590698 80614
rect 590142 60378 590378 60614
rect 590462 60378 590698 60614
rect 590142 40378 590378 40614
rect 590462 40378 590698 40614
rect 590142 20378 590378 20614
rect 590462 20378 590698 20614
rect 579266 -5382 579502 -5146
rect 579586 -5382 579822 -5146
rect 579266 -5702 579502 -5466
rect 579586 -5702 579822 -5466
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 694038 591338 694274
rect 591422 694038 591658 694274
rect 591102 674038 591338 674274
rect 591422 674038 591658 674274
rect 591102 654038 591338 654274
rect 591422 654038 591658 654274
rect 591102 634038 591338 634274
rect 591422 634038 591658 634274
rect 591102 614038 591338 614274
rect 591422 614038 591658 614274
rect 591102 594038 591338 594274
rect 591422 594038 591658 594274
rect 591102 574038 591338 574274
rect 591422 574038 591658 574274
rect 591102 554038 591338 554274
rect 591422 554038 591658 554274
rect 591102 534038 591338 534274
rect 591422 534038 591658 534274
rect 591102 514038 591338 514274
rect 591422 514038 591658 514274
rect 591102 494038 591338 494274
rect 591422 494038 591658 494274
rect 591102 474038 591338 474274
rect 591422 474038 591658 474274
rect 591102 454038 591338 454274
rect 591422 454038 591658 454274
rect 591102 434038 591338 434274
rect 591422 434038 591658 434274
rect 591102 414038 591338 414274
rect 591422 414038 591658 414274
rect 591102 394038 591338 394274
rect 591422 394038 591658 394274
rect 591102 374038 591338 374274
rect 591422 374038 591658 374274
rect 591102 354038 591338 354274
rect 591422 354038 591658 354274
rect 591102 334038 591338 334274
rect 591422 334038 591658 334274
rect 591102 314038 591338 314274
rect 591422 314038 591658 314274
rect 591102 294038 591338 294274
rect 591422 294038 591658 294274
rect 591102 274038 591338 274274
rect 591422 274038 591658 274274
rect 591102 254038 591338 254274
rect 591422 254038 591658 254274
rect 591102 234038 591338 234274
rect 591422 234038 591658 234274
rect 591102 214038 591338 214274
rect 591422 214038 591658 214274
rect 591102 194038 591338 194274
rect 591422 194038 591658 194274
rect 591102 174038 591338 174274
rect 591422 174038 591658 174274
rect 591102 154038 591338 154274
rect 591422 154038 591658 154274
rect 591102 134038 591338 134274
rect 591422 134038 591658 134274
rect 591102 114038 591338 114274
rect 591422 114038 591658 114274
rect 591102 94038 591338 94274
rect 591422 94038 591658 94274
rect 591102 74038 591338 74274
rect 591422 74038 591658 74274
rect 591102 54038 591338 54274
rect 591422 54038 591658 54274
rect 591102 34038 591338 34274
rect 591422 34038 591658 34274
rect 591102 14038 591338 14274
rect 591422 14038 591658 14274
rect 572986 -6342 573222 -6106
rect 573306 -6342 573542 -6106
rect 572986 -6662 573222 -6426
rect 573306 -6662 573542 -6426
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 684038 592298 684274
rect 592382 684038 592618 684274
rect 592062 664038 592298 664274
rect 592382 664038 592618 664274
rect 592062 644038 592298 644274
rect 592382 644038 592618 644274
rect 592062 624038 592298 624274
rect 592382 624038 592618 624274
rect 592062 604038 592298 604274
rect 592382 604038 592618 604274
rect 592062 584038 592298 584274
rect 592382 584038 592618 584274
rect 592062 564038 592298 564274
rect 592382 564038 592618 564274
rect 592062 544038 592298 544274
rect 592382 544038 592618 544274
rect 592062 524038 592298 524274
rect 592382 524038 592618 524274
rect 592062 504038 592298 504274
rect 592382 504038 592618 504274
rect 592062 484038 592298 484274
rect 592382 484038 592618 484274
rect 592062 464038 592298 464274
rect 592382 464038 592618 464274
rect 592062 444038 592298 444274
rect 592382 444038 592618 444274
rect 592062 424038 592298 424274
rect 592382 424038 592618 424274
rect 592062 404038 592298 404274
rect 592382 404038 592618 404274
rect 592062 384038 592298 384274
rect 592382 384038 592618 384274
rect 592062 364038 592298 364274
rect 592382 364038 592618 364274
rect 592062 344038 592298 344274
rect 592382 344038 592618 344274
rect 592062 324038 592298 324274
rect 592382 324038 592618 324274
rect 592062 304038 592298 304274
rect 592382 304038 592618 304274
rect 592062 284038 592298 284274
rect 592382 284038 592618 284274
rect 592062 264038 592298 264274
rect 592382 264038 592618 264274
rect 592062 244038 592298 244274
rect 592382 244038 592618 244274
rect 592062 224038 592298 224274
rect 592382 224038 592618 224274
rect 592062 204038 592298 204274
rect 592382 204038 592618 204274
rect 592062 184038 592298 184274
rect 592382 184038 592618 184274
rect 592062 164038 592298 164274
rect 592382 164038 592618 164274
rect 592062 144038 592298 144274
rect 592382 144038 592618 144274
rect 592062 124038 592298 124274
rect 592382 124038 592618 124274
rect 592062 104038 592298 104274
rect 592382 104038 592618 104274
rect 592062 84038 592298 84274
rect 592382 84038 592618 84274
rect 592062 64038 592298 64274
rect 592382 64038 592618 64274
rect 592062 44038 592298 44274
rect 592382 44038 592618 44274
rect 592062 24038 592298 24274
rect 592382 24038 592618 24274
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 22986 711558
rect 23222 711322 23306 711558
rect 23542 711322 42986 711558
rect 43222 711322 43306 711558
rect 43542 711322 62986 711558
rect 63222 711322 63306 711558
rect 63542 711322 82986 711558
rect 83222 711322 83306 711558
rect 83542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 122986 711558
rect 123222 711322 123306 711558
rect 123542 711322 142986 711558
rect 143222 711322 143306 711558
rect 143542 711322 162986 711558
rect 163222 711322 163306 711558
rect 163542 711322 182986 711558
rect 183222 711322 183306 711558
rect 183542 711322 202986 711558
rect 203222 711322 203306 711558
rect 203542 711322 222986 711558
rect 223222 711322 223306 711558
rect 223542 711322 242986 711558
rect 243222 711322 243306 711558
rect 243542 711322 262986 711558
rect 263222 711322 263306 711558
rect 263542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 302986 711558
rect 303222 711322 303306 711558
rect 303542 711322 322986 711558
rect 323222 711322 323306 711558
rect 323542 711322 342986 711558
rect 343222 711322 343306 711558
rect 343542 711322 362986 711558
rect 363222 711322 363306 711558
rect 363542 711322 382986 711558
rect 383222 711322 383306 711558
rect 383542 711322 402986 711558
rect 403222 711322 403306 711558
rect 403542 711322 422986 711558
rect 423222 711322 423306 711558
rect 423542 711322 442986 711558
rect 443222 711322 443306 711558
rect 443542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 482986 711558
rect 483222 711322 483306 711558
rect 483542 711322 502986 711558
rect 503222 711322 503306 711558
rect 503542 711322 522986 711558
rect 523222 711322 523306 711558
rect 523542 711322 542986 711558
rect 543222 711322 543306 711558
rect 543542 711322 562986 711558
rect 563222 711322 563306 711558
rect 563542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 22986 711238
rect 23222 711002 23306 711238
rect 23542 711002 42986 711238
rect 43222 711002 43306 711238
rect 43542 711002 62986 711238
rect 63222 711002 63306 711238
rect 63542 711002 82986 711238
rect 83222 711002 83306 711238
rect 83542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 122986 711238
rect 123222 711002 123306 711238
rect 123542 711002 142986 711238
rect 143222 711002 143306 711238
rect 143542 711002 162986 711238
rect 163222 711002 163306 711238
rect 163542 711002 182986 711238
rect 183222 711002 183306 711238
rect 183542 711002 202986 711238
rect 203222 711002 203306 711238
rect 203542 711002 222986 711238
rect 223222 711002 223306 711238
rect 223542 711002 242986 711238
rect 243222 711002 243306 711238
rect 243542 711002 262986 711238
rect 263222 711002 263306 711238
rect 263542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 302986 711238
rect 303222 711002 303306 711238
rect 303542 711002 322986 711238
rect 323222 711002 323306 711238
rect 323542 711002 342986 711238
rect 343222 711002 343306 711238
rect 343542 711002 362986 711238
rect 363222 711002 363306 711238
rect 363542 711002 382986 711238
rect 383222 711002 383306 711238
rect 383542 711002 402986 711238
rect 403222 711002 403306 711238
rect 403542 711002 422986 711238
rect 423222 711002 423306 711238
rect 423542 711002 442986 711238
rect 443222 711002 443306 711238
rect 443542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 482986 711238
rect 483222 711002 483306 711238
rect 483542 711002 502986 711238
rect 503222 711002 503306 711238
rect 503542 711002 522986 711238
rect 523222 711002 523306 711238
rect 523542 711002 542986 711238
rect 543222 711002 543306 711238
rect 543542 711002 562986 711238
rect 563222 711002 563306 711238
rect 563542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 32986 710598
rect 33222 710362 33306 710598
rect 33542 710362 52986 710598
rect 53222 710362 53306 710598
rect 53542 710362 72986 710598
rect 73222 710362 73306 710598
rect 73542 710362 92986 710598
rect 93222 710362 93306 710598
rect 93542 710362 112986 710598
rect 113222 710362 113306 710598
rect 113542 710362 132986 710598
rect 133222 710362 133306 710598
rect 133542 710362 152986 710598
rect 153222 710362 153306 710598
rect 153542 710362 172986 710598
rect 173222 710362 173306 710598
rect 173542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 212986 710598
rect 213222 710362 213306 710598
rect 213542 710362 232986 710598
rect 233222 710362 233306 710598
rect 233542 710362 252986 710598
rect 253222 710362 253306 710598
rect 253542 710362 272986 710598
rect 273222 710362 273306 710598
rect 273542 710362 292986 710598
rect 293222 710362 293306 710598
rect 293542 710362 312986 710598
rect 313222 710362 313306 710598
rect 313542 710362 332986 710598
rect 333222 710362 333306 710598
rect 333542 710362 352986 710598
rect 353222 710362 353306 710598
rect 353542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 392986 710598
rect 393222 710362 393306 710598
rect 393542 710362 412986 710598
rect 413222 710362 413306 710598
rect 413542 710362 432986 710598
rect 433222 710362 433306 710598
rect 433542 710362 452986 710598
rect 453222 710362 453306 710598
rect 453542 710362 472986 710598
rect 473222 710362 473306 710598
rect 473542 710362 492986 710598
rect 493222 710362 493306 710598
rect 493542 710362 512986 710598
rect 513222 710362 513306 710598
rect 513542 710362 532986 710598
rect 533222 710362 533306 710598
rect 533542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 572986 710598
rect 573222 710362 573306 710598
rect 573542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 32986 710278
rect 33222 710042 33306 710278
rect 33542 710042 52986 710278
rect 53222 710042 53306 710278
rect 53542 710042 72986 710278
rect 73222 710042 73306 710278
rect 73542 710042 92986 710278
rect 93222 710042 93306 710278
rect 93542 710042 112986 710278
rect 113222 710042 113306 710278
rect 113542 710042 132986 710278
rect 133222 710042 133306 710278
rect 133542 710042 152986 710278
rect 153222 710042 153306 710278
rect 153542 710042 172986 710278
rect 173222 710042 173306 710278
rect 173542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 212986 710278
rect 213222 710042 213306 710278
rect 213542 710042 232986 710278
rect 233222 710042 233306 710278
rect 233542 710042 252986 710278
rect 253222 710042 253306 710278
rect 253542 710042 272986 710278
rect 273222 710042 273306 710278
rect 273542 710042 292986 710278
rect 293222 710042 293306 710278
rect 293542 710042 312986 710278
rect 313222 710042 313306 710278
rect 313542 710042 332986 710278
rect 333222 710042 333306 710278
rect 333542 710042 352986 710278
rect 353222 710042 353306 710278
rect 353542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 392986 710278
rect 393222 710042 393306 710278
rect 393542 710042 412986 710278
rect 413222 710042 413306 710278
rect 413542 710042 432986 710278
rect 433222 710042 433306 710278
rect 433542 710042 452986 710278
rect 453222 710042 453306 710278
rect 453542 710042 472986 710278
rect 473222 710042 473306 710278
rect 473542 710042 492986 710278
rect 493222 710042 493306 710278
rect 493542 710042 512986 710278
rect 513222 710042 513306 710278
rect 513542 710042 532986 710278
rect 533222 710042 533306 710278
rect 533542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 572986 710278
rect 573222 710042 573306 710278
rect 573542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 19266 709638
rect 19502 709402 19586 709638
rect 19822 709402 39266 709638
rect 39502 709402 39586 709638
rect 39822 709402 59266 709638
rect 59502 709402 59586 709638
rect 59822 709402 79266 709638
rect 79502 709402 79586 709638
rect 79822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 119266 709638
rect 119502 709402 119586 709638
rect 119822 709402 139266 709638
rect 139502 709402 139586 709638
rect 139822 709402 159266 709638
rect 159502 709402 159586 709638
rect 159822 709402 179266 709638
rect 179502 709402 179586 709638
rect 179822 709402 199266 709638
rect 199502 709402 199586 709638
rect 199822 709402 219266 709638
rect 219502 709402 219586 709638
rect 219822 709402 239266 709638
rect 239502 709402 239586 709638
rect 239822 709402 259266 709638
rect 259502 709402 259586 709638
rect 259822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 299266 709638
rect 299502 709402 299586 709638
rect 299822 709402 319266 709638
rect 319502 709402 319586 709638
rect 319822 709402 339266 709638
rect 339502 709402 339586 709638
rect 339822 709402 359266 709638
rect 359502 709402 359586 709638
rect 359822 709402 379266 709638
rect 379502 709402 379586 709638
rect 379822 709402 399266 709638
rect 399502 709402 399586 709638
rect 399822 709402 419266 709638
rect 419502 709402 419586 709638
rect 419822 709402 439266 709638
rect 439502 709402 439586 709638
rect 439822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 479266 709638
rect 479502 709402 479586 709638
rect 479822 709402 499266 709638
rect 499502 709402 499586 709638
rect 499822 709402 519266 709638
rect 519502 709402 519586 709638
rect 519822 709402 539266 709638
rect 539502 709402 539586 709638
rect 539822 709402 559266 709638
rect 559502 709402 559586 709638
rect 559822 709402 579266 709638
rect 579502 709402 579586 709638
rect 579822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 19266 709318
rect 19502 709082 19586 709318
rect 19822 709082 39266 709318
rect 39502 709082 39586 709318
rect 39822 709082 59266 709318
rect 59502 709082 59586 709318
rect 59822 709082 79266 709318
rect 79502 709082 79586 709318
rect 79822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 119266 709318
rect 119502 709082 119586 709318
rect 119822 709082 139266 709318
rect 139502 709082 139586 709318
rect 139822 709082 159266 709318
rect 159502 709082 159586 709318
rect 159822 709082 179266 709318
rect 179502 709082 179586 709318
rect 179822 709082 199266 709318
rect 199502 709082 199586 709318
rect 199822 709082 219266 709318
rect 219502 709082 219586 709318
rect 219822 709082 239266 709318
rect 239502 709082 239586 709318
rect 239822 709082 259266 709318
rect 259502 709082 259586 709318
rect 259822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 299266 709318
rect 299502 709082 299586 709318
rect 299822 709082 319266 709318
rect 319502 709082 319586 709318
rect 319822 709082 339266 709318
rect 339502 709082 339586 709318
rect 339822 709082 359266 709318
rect 359502 709082 359586 709318
rect 359822 709082 379266 709318
rect 379502 709082 379586 709318
rect 379822 709082 399266 709318
rect 399502 709082 399586 709318
rect 399822 709082 419266 709318
rect 419502 709082 419586 709318
rect 419822 709082 439266 709318
rect 439502 709082 439586 709318
rect 439822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 479266 709318
rect 479502 709082 479586 709318
rect 479822 709082 499266 709318
rect 499502 709082 499586 709318
rect 499822 709082 519266 709318
rect 519502 709082 519586 709318
rect 519822 709082 539266 709318
rect 539502 709082 539586 709318
rect 539822 709082 559266 709318
rect 559502 709082 559586 709318
rect 559822 709082 579266 709318
rect 579502 709082 579586 709318
rect 579822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 29266 708678
rect 29502 708442 29586 708678
rect 29822 708442 49266 708678
rect 49502 708442 49586 708678
rect 49822 708442 69266 708678
rect 69502 708442 69586 708678
rect 69822 708442 89266 708678
rect 89502 708442 89586 708678
rect 89822 708442 109266 708678
rect 109502 708442 109586 708678
rect 109822 708442 129266 708678
rect 129502 708442 129586 708678
rect 129822 708442 149266 708678
rect 149502 708442 149586 708678
rect 149822 708442 169266 708678
rect 169502 708442 169586 708678
rect 169822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 209266 708678
rect 209502 708442 209586 708678
rect 209822 708442 229266 708678
rect 229502 708442 229586 708678
rect 229822 708442 249266 708678
rect 249502 708442 249586 708678
rect 249822 708442 269266 708678
rect 269502 708442 269586 708678
rect 269822 708442 289266 708678
rect 289502 708442 289586 708678
rect 289822 708442 309266 708678
rect 309502 708442 309586 708678
rect 309822 708442 329266 708678
rect 329502 708442 329586 708678
rect 329822 708442 349266 708678
rect 349502 708442 349586 708678
rect 349822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 389266 708678
rect 389502 708442 389586 708678
rect 389822 708442 409266 708678
rect 409502 708442 409586 708678
rect 409822 708442 429266 708678
rect 429502 708442 429586 708678
rect 429822 708442 449266 708678
rect 449502 708442 449586 708678
rect 449822 708442 469266 708678
rect 469502 708442 469586 708678
rect 469822 708442 489266 708678
rect 489502 708442 489586 708678
rect 489822 708442 509266 708678
rect 509502 708442 509586 708678
rect 509822 708442 529266 708678
rect 529502 708442 529586 708678
rect 529822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 569266 708678
rect 569502 708442 569586 708678
rect 569822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 29266 708358
rect 29502 708122 29586 708358
rect 29822 708122 49266 708358
rect 49502 708122 49586 708358
rect 49822 708122 69266 708358
rect 69502 708122 69586 708358
rect 69822 708122 89266 708358
rect 89502 708122 89586 708358
rect 89822 708122 109266 708358
rect 109502 708122 109586 708358
rect 109822 708122 129266 708358
rect 129502 708122 129586 708358
rect 129822 708122 149266 708358
rect 149502 708122 149586 708358
rect 149822 708122 169266 708358
rect 169502 708122 169586 708358
rect 169822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 209266 708358
rect 209502 708122 209586 708358
rect 209822 708122 229266 708358
rect 229502 708122 229586 708358
rect 229822 708122 249266 708358
rect 249502 708122 249586 708358
rect 249822 708122 269266 708358
rect 269502 708122 269586 708358
rect 269822 708122 289266 708358
rect 289502 708122 289586 708358
rect 289822 708122 309266 708358
rect 309502 708122 309586 708358
rect 309822 708122 329266 708358
rect 329502 708122 329586 708358
rect 329822 708122 349266 708358
rect 349502 708122 349586 708358
rect 349822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 389266 708358
rect 389502 708122 389586 708358
rect 389822 708122 409266 708358
rect 409502 708122 409586 708358
rect 409822 708122 429266 708358
rect 429502 708122 429586 708358
rect 429822 708122 449266 708358
rect 449502 708122 449586 708358
rect 449822 708122 469266 708358
rect 469502 708122 469586 708358
rect 469822 708122 489266 708358
rect 489502 708122 489586 708358
rect 489822 708122 509266 708358
rect 509502 708122 509586 708358
rect 509822 708122 529266 708358
rect 529502 708122 529586 708358
rect 529822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 569266 708358
rect 569502 708122 569586 708358
rect 569822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15546 707718
rect 15782 707482 15866 707718
rect 16102 707482 35546 707718
rect 35782 707482 35866 707718
rect 36102 707482 55546 707718
rect 55782 707482 55866 707718
rect 56102 707482 75546 707718
rect 75782 707482 75866 707718
rect 76102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 115546 707718
rect 115782 707482 115866 707718
rect 116102 707482 135546 707718
rect 135782 707482 135866 707718
rect 136102 707482 155546 707718
rect 155782 707482 155866 707718
rect 156102 707482 175546 707718
rect 175782 707482 175866 707718
rect 176102 707482 195546 707718
rect 195782 707482 195866 707718
rect 196102 707482 215546 707718
rect 215782 707482 215866 707718
rect 216102 707482 235546 707718
rect 235782 707482 235866 707718
rect 236102 707482 255546 707718
rect 255782 707482 255866 707718
rect 256102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 295546 707718
rect 295782 707482 295866 707718
rect 296102 707482 315546 707718
rect 315782 707482 315866 707718
rect 316102 707482 335546 707718
rect 335782 707482 335866 707718
rect 336102 707482 355546 707718
rect 355782 707482 355866 707718
rect 356102 707482 375546 707718
rect 375782 707482 375866 707718
rect 376102 707482 395546 707718
rect 395782 707482 395866 707718
rect 396102 707482 415546 707718
rect 415782 707482 415866 707718
rect 416102 707482 435546 707718
rect 435782 707482 435866 707718
rect 436102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 475546 707718
rect 475782 707482 475866 707718
rect 476102 707482 495546 707718
rect 495782 707482 495866 707718
rect 496102 707482 515546 707718
rect 515782 707482 515866 707718
rect 516102 707482 535546 707718
rect 535782 707482 535866 707718
rect 536102 707482 555546 707718
rect 555782 707482 555866 707718
rect 556102 707482 575546 707718
rect 575782 707482 575866 707718
rect 576102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15546 707398
rect 15782 707162 15866 707398
rect 16102 707162 35546 707398
rect 35782 707162 35866 707398
rect 36102 707162 55546 707398
rect 55782 707162 55866 707398
rect 56102 707162 75546 707398
rect 75782 707162 75866 707398
rect 76102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 115546 707398
rect 115782 707162 115866 707398
rect 116102 707162 135546 707398
rect 135782 707162 135866 707398
rect 136102 707162 155546 707398
rect 155782 707162 155866 707398
rect 156102 707162 175546 707398
rect 175782 707162 175866 707398
rect 176102 707162 195546 707398
rect 195782 707162 195866 707398
rect 196102 707162 215546 707398
rect 215782 707162 215866 707398
rect 216102 707162 235546 707398
rect 235782 707162 235866 707398
rect 236102 707162 255546 707398
rect 255782 707162 255866 707398
rect 256102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 295546 707398
rect 295782 707162 295866 707398
rect 296102 707162 315546 707398
rect 315782 707162 315866 707398
rect 316102 707162 335546 707398
rect 335782 707162 335866 707398
rect 336102 707162 355546 707398
rect 355782 707162 355866 707398
rect 356102 707162 375546 707398
rect 375782 707162 375866 707398
rect 376102 707162 395546 707398
rect 395782 707162 395866 707398
rect 396102 707162 415546 707398
rect 415782 707162 415866 707398
rect 416102 707162 435546 707398
rect 435782 707162 435866 707398
rect 436102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 475546 707398
rect 475782 707162 475866 707398
rect 476102 707162 495546 707398
rect 495782 707162 495866 707398
rect 496102 707162 515546 707398
rect 515782 707162 515866 707398
rect 516102 707162 535546 707398
rect 535782 707162 535866 707398
rect 536102 707162 555546 707398
rect 555782 707162 555866 707398
rect 556102 707162 575546 707398
rect 575782 707162 575866 707398
rect 576102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 25546 706758
rect 25782 706522 25866 706758
rect 26102 706522 45546 706758
rect 45782 706522 45866 706758
rect 46102 706522 65546 706758
rect 65782 706522 65866 706758
rect 66102 706522 85546 706758
rect 85782 706522 85866 706758
rect 86102 706522 105546 706758
rect 105782 706522 105866 706758
rect 106102 706522 125546 706758
rect 125782 706522 125866 706758
rect 126102 706522 145546 706758
rect 145782 706522 145866 706758
rect 146102 706522 165546 706758
rect 165782 706522 165866 706758
rect 166102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 205546 706758
rect 205782 706522 205866 706758
rect 206102 706522 225546 706758
rect 225782 706522 225866 706758
rect 226102 706522 245546 706758
rect 245782 706522 245866 706758
rect 246102 706522 265546 706758
rect 265782 706522 265866 706758
rect 266102 706522 285546 706758
rect 285782 706522 285866 706758
rect 286102 706522 305546 706758
rect 305782 706522 305866 706758
rect 306102 706522 325546 706758
rect 325782 706522 325866 706758
rect 326102 706522 345546 706758
rect 345782 706522 345866 706758
rect 346102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 385546 706758
rect 385782 706522 385866 706758
rect 386102 706522 405546 706758
rect 405782 706522 405866 706758
rect 406102 706522 425546 706758
rect 425782 706522 425866 706758
rect 426102 706522 445546 706758
rect 445782 706522 445866 706758
rect 446102 706522 465546 706758
rect 465782 706522 465866 706758
rect 466102 706522 485546 706758
rect 485782 706522 485866 706758
rect 486102 706522 505546 706758
rect 505782 706522 505866 706758
rect 506102 706522 525546 706758
rect 525782 706522 525866 706758
rect 526102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 565546 706758
rect 565782 706522 565866 706758
rect 566102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 25546 706438
rect 25782 706202 25866 706438
rect 26102 706202 45546 706438
rect 45782 706202 45866 706438
rect 46102 706202 65546 706438
rect 65782 706202 65866 706438
rect 66102 706202 85546 706438
rect 85782 706202 85866 706438
rect 86102 706202 105546 706438
rect 105782 706202 105866 706438
rect 106102 706202 125546 706438
rect 125782 706202 125866 706438
rect 126102 706202 145546 706438
rect 145782 706202 145866 706438
rect 146102 706202 165546 706438
rect 165782 706202 165866 706438
rect 166102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 205546 706438
rect 205782 706202 205866 706438
rect 206102 706202 225546 706438
rect 225782 706202 225866 706438
rect 226102 706202 245546 706438
rect 245782 706202 245866 706438
rect 246102 706202 265546 706438
rect 265782 706202 265866 706438
rect 266102 706202 285546 706438
rect 285782 706202 285866 706438
rect 286102 706202 305546 706438
rect 305782 706202 305866 706438
rect 306102 706202 325546 706438
rect 325782 706202 325866 706438
rect 326102 706202 345546 706438
rect 345782 706202 345866 706438
rect 346102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 385546 706438
rect 385782 706202 385866 706438
rect 386102 706202 405546 706438
rect 405782 706202 405866 706438
rect 406102 706202 425546 706438
rect 425782 706202 425866 706438
rect 426102 706202 445546 706438
rect 445782 706202 445866 706438
rect 446102 706202 465546 706438
rect 465782 706202 465866 706438
rect 466102 706202 485546 706438
rect 485782 706202 485866 706438
rect 486102 706202 505546 706438
rect 505782 706202 505866 706438
rect 506102 706202 525546 706438
rect 525782 706202 525866 706438
rect 526102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 565546 706438
rect 565782 706202 565866 706438
rect 566102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 11826 705798
rect 12062 705562 12146 705798
rect 12382 705562 31826 705798
rect 32062 705562 32146 705798
rect 32382 705562 51826 705798
rect 52062 705562 52146 705798
rect 52382 705562 71826 705798
rect 72062 705562 72146 705798
rect 72382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 111826 705798
rect 112062 705562 112146 705798
rect 112382 705562 131826 705798
rect 132062 705562 132146 705798
rect 132382 705562 151826 705798
rect 152062 705562 152146 705798
rect 152382 705562 171826 705798
rect 172062 705562 172146 705798
rect 172382 705562 191826 705798
rect 192062 705562 192146 705798
rect 192382 705562 211826 705798
rect 212062 705562 212146 705798
rect 212382 705562 231826 705798
rect 232062 705562 232146 705798
rect 232382 705562 251826 705798
rect 252062 705562 252146 705798
rect 252382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 291826 705798
rect 292062 705562 292146 705798
rect 292382 705562 311826 705798
rect 312062 705562 312146 705798
rect 312382 705562 331826 705798
rect 332062 705562 332146 705798
rect 332382 705562 351826 705798
rect 352062 705562 352146 705798
rect 352382 705562 371826 705798
rect 372062 705562 372146 705798
rect 372382 705562 391826 705798
rect 392062 705562 392146 705798
rect 392382 705562 411826 705798
rect 412062 705562 412146 705798
rect 412382 705562 431826 705798
rect 432062 705562 432146 705798
rect 432382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 471826 705798
rect 472062 705562 472146 705798
rect 472382 705562 491826 705798
rect 492062 705562 492146 705798
rect 492382 705562 511826 705798
rect 512062 705562 512146 705798
rect 512382 705562 531826 705798
rect 532062 705562 532146 705798
rect 532382 705562 551826 705798
rect 552062 705562 552146 705798
rect 552382 705562 571826 705798
rect 572062 705562 572146 705798
rect 572382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 11826 705478
rect 12062 705242 12146 705478
rect 12382 705242 31826 705478
rect 32062 705242 32146 705478
rect 32382 705242 51826 705478
rect 52062 705242 52146 705478
rect 52382 705242 71826 705478
rect 72062 705242 72146 705478
rect 72382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 111826 705478
rect 112062 705242 112146 705478
rect 112382 705242 131826 705478
rect 132062 705242 132146 705478
rect 132382 705242 151826 705478
rect 152062 705242 152146 705478
rect 152382 705242 171826 705478
rect 172062 705242 172146 705478
rect 172382 705242 191826 705478
rect 192062 705242 192146 705478
rect 192382 705242 211826 705478
rect 212062 705242 212146 705478
rect 212382 705242 231826 705478
rect 232062 705242 232146 705478
rect 232382 705242 251826 705478
rect 252062 705242 252146 705478
rect 252382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 291826 705478
rect 292062 705242 292146 705478
rect 292382 705242 311826 705478
rect 312062 705242 312146 705478
rect 312382 705242 331826 705478
rect 332062 705242 332146 705478
rect 332382 705242 351826 705478
rect 352062 705242 352146 705478
rect 352382 705242 371826 705478
rect 372062 705242 372146 705478
rect 372382 705242 391826 705478
rect 392062 705242 392146 705478
rect 392382 705242 411826 705478
rect 412062 705242 412146 705478
rect 412382 705242 431826 705478
rect 432062 705242 432146 705478
rect 432382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 471826 705478
rect 472062 705242 472146 705478
rect 472382 705242 491826 705478
rect 492062 705242 492146 705478
rect 492382 705242 511826 705478
rect 512062 705242 512146 705478
rect 512382 705242 531826 705478
rect 532062 705242 532146 705478
rect 532382 705242 551826 705478
rect 552062 705242 552146 705478
rect 552382 705242 571826 705478
rect 572062 705242 572146 705478
rect 572382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 21826 704838
rect 22062 704602 22146 704838
rect 22382 704602 41826 704838
rect 42062 704602 42146 704838
rect 42382 704602 61826 704838
rect 62062 704602 62146 704838
rect 62382 704602 81826 704838
rect 82062 704602 82146 704838
rect 82382 704602 101826 704838
rect 102062 704602 102146 704838
rect 102382 704602 121826 704838
rect 122062 704602 122146 704838
rect 122382 704602 141826 704838
rect 142062 704602 142146 704838
rect 142382 704602 161826 704838
rect 162062 704602 162146 704838
rect 162382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 201826 704838
rect 202062 704602 202146 704838
rect 202382 704602 221826 704838
rect 222062 704602 222146 704838
rect 222382 704602 241826 704838
rect 242062 704602 242146 704838
rect 242382 704602 261826 704838
rect 262062 704602 262146 704838
rect 262382 704602 281826 704838
rect 282062 704602 282146 704838
rect 282382 704602 301826 704838
rect 302062 704602 302146 704838
rect 302382 704602 321826 704838
rect 322062 704602 322146 704838
rect 322382 704602 341826 704838
rect 342062 704602 342146 704838
rect 342382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 381826 704838
rect 382062 704602 382146 704838
rect 382382 704602 401826 704838
rect 402062 704602 402146 704838
rect 402382 704602 421826 704838
rect 422062 704602 422146 704838
rect 422382 704602 441826 704838
rect 442062 704602 442146 704838
rect 442382 704602 461826 704838
rect 462062 704602 462146 704838
rect 462382 704602 481826 704838
rect 482062 704602 482146 704838
rect 482382 704602 501826 704838
rect 502062 704602 502146 704838
rect 502382 704602 521826 704838
rect 522062 704602 522146 704838
rect 522382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 561826 704838
rect 562062 704602 562146 704838
rect 562382 704602 581826 704838
rect 582062 704602 582146 704838
rect 582382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 21826 704518
rect 22062 704282 22146 704518
rect 22382 704282 41826 704518
rect 42062 704282 42146 704518
rect 42382 704282 61826 704518
rect 62062 704282 62146 704518
rect 62382 704282 81826 704518
rect 82062 704282 82146 704518
rect 82382 704282 101826 704518
rect 102062 704282 102146 704518
rect 102382 704282 121826 704518
rect 122062 704282 122146 704518
rect 122382 704282 141826 704518
rect 142062 704282 142146 704518
rect 142382 704282 161826 704518
rect 162062 704282 162146 704518
rect 162382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 201826 704518
rect 202062 704282 202146 704518
rect 202382 704282 221826 704518
rect 222062 704282 222146 704518
rect 222382 704282 241826 704518
rect 242062 704282 242146 704518
rect 242382 704282 261826 704518
rect 262062 704282 262146 704518
rect 262382 704282 281826 704518
rect 282062 704282 282146 704518
rect 282382 704282 301826 704518
rect 302062 704282 302146 704518
rect 302382 704282 321826 704518
rect 322062 704282 322146 704518
rect 322382 704282 341826 704518
rect 342062 704282 342146 704518
rect 342382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 381826 704518
rect 382062 704282 382146 704518
rect 382382 704282 401826 704518
rect 402062 704282 402146 704518
rect 402382 704282 421826 704518
rect 422062 704282 422146 704518
rect 422382 704282 441826 704518
rect 442062 704282 442146 704518
rect 442382 704282 461826 704518
rect 462062 704282 462146 704518
rect 462382 704282 481826 704518
rect 482062 704282 482146 704518
rect 482382 704282 501826 704518
rect 502062 704282 502146 704518
rect 502382 704282 521826 704518
rect 522062 704282 522146 704518
rect 522382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 561826 704518
rect 562062 704282 562146 704518
rect 562382 704282 581826 704518
rect 582062 704282 582146 704518
rect 582382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -6806 700614 590730 700776
rect -6806 700378 -6774 700614
rect -6538 700378 -6454 700614
rect -6218 700378 19266 700614
rect 19502 700378 19586 700614
rect 19822 700378 39266 700614
rect 39502 700378 39586 700614
rect 39822 700378 59266 700614
rect 59502 700378 59586 700614
rect 59822 700378 79266 700614
rect 79502 700378 79586 700614
rect 79822 700378 99266 700614
rect 99502 700378 99586 700614
rect 99822 700378 119266 700614
rect 119502 700378 119586 700614
rect 119822 700378 139266 700614
rect 139502 700378 139586 700614
rect 139822 700378 159266 700614
rect 159502 700378 159586 700614
rect 159822 700378 179266 700614
rect 179502 700378 179586 700614
rect 179822 700378 199266 700614
rect 199502 700378 199586 700614
rect 199822 700378 219266 700614
rect 219502 700378 219586 700614
rect 219822 700378 239266 700614
rect 239502 700378 239586 700614
rect 239822 700378 259266 700614
rect 259502 700378 259586 700614
rect 259822 700378 279266 700614
rect 279502 700378 279586 700614
rect 279822 700378 299266 700614
rect 299502 700378 299586 700614
rect 299822 700378 319266 700614
rect 319502 700378 319586 700614
rect 319822 700378 339266 700614
rect 339502 700378 339586 700614
rect 339822 700378 359266 700614
rect 359502 700378 359586 700614
rect 359822 700378 379266 700614
rect 379502 700378 379586 700614
rect 379822 700378 399266 700614
rect 399502 700378 399586 700614
rect 399822 700378 419266 700614
rect 419502 700378 419586 700614
rect 419822 700378 439266 700614
rect 439502 700378 439586 700614
rect 439822 700378 459266 700614
rect 459502 700378 459586 700614
rect 459822 700378 479266 700614
rect 479502 700378 479586 700614
rect 479822 700378 499266 700614
rect 499502 700378 499586 700614
rect 499822 700378 519266 700614
rect 519502 700378 519586 700614
rect 519822 700378 539266 700614
rect 539502 700378 539586 700614
rect 539822 700378 559266 700614
rect 559502 700378 559586 700614
rect 559822 700378 579266 700614
rect 579502 700378 579586 700614
rect 579822 700378 590142 700614
rect 590378 700378 590462 700614
rect 590698 700378 590730 700614
rect -6806 700216 590730 700378
rect -4886 696954 588810 697116
rect -4886 696718 -4854 696954
rect -4618 696718 -4534 696954
rect -4298 696718 15546 696954
rect 15782 696718 15866 696954
rect 16102 696718 35546 696954
rect 35782 696718 35866 696954
rect 36102 696718 55546 696954
rect 55782 696718 55866 696954
rect 56102 696718 75546 696954
rect 75782 696718 75866 696954
rect 76102 696718 95546 696954
rect 95782 696718 95866 696954
rect 96102 696718 115546 696954
rect 115782 696718 115866 696954
rect 116102 696718 135546 696954
rect 135782 696718 135866 696954
rect 136102 696718 155546 696954
rect 155782 696718 155866 696954
rect 156102 696718 175546 696954
rect 175782 696718 175866 696954
rect 176102 696718 195546 696954
rect 195782 696718 195866 696954
rect 196102 696718 215546 696954
rect 215782 696718 215866 696954
rect 216102 696718 235546 696954
rect 235782 696718 235866 696954
rect 236102 696718 255546 696954
rect 255782 696718 255866 696954
rect 256102 696718 275546 696954
rect 275782 696718 275866 696954
rect 276102 696718 295546 696954
rect 295782 696718 295866 696954
rect 296102 696718 315546 696954
rect 315782 696718 315866 696954
rect 316102 696718 335546 696954
rect 335782 696718 335866 696954
rect 336102 696718 355546 696954
rect 355782 696718 355866 696954
rect 356102 696718 375546 696954
rect 375782 696718 375866 696954
rect 376102 696718 395546 696954
rect 395782 696718 395866 696954
rect 396102 696718 415546 696954
rect 415782 696718 415866 696954
rect 416102 696718 435546 696954
rect 435782 696718 435866 696954
rect 436102 696718 455546 696954
rect 455782 696718 455866 696954
rect 456102 696718 475546 696954
rect 475782 696718 475866 696954
rect 476102 696718 495546 696954
rect 495782 696718 495866 696954
rect 496102 696718 515546 696954
rect 515782 696718 515866 696954
rect 516102 696718 535546 696954
rect 535782 696718 535866 696954
rect 536102 696718 555546 696954
rect 555782 696718 555866 696954
rect 556102 696718 575546 696954
rect 575782 696718 575866 696954
rect 576102 696718 588222 696954
rect 588458 696718 588542 696954
rect 588778 696718 588810 696954
rect -4886 696556 588810 696718
rect -8726 694274 592650 694436
rect -8726 694038 -7734 694274
rect -7498 694038 -7414 694274
rect -7178 694038 12986 694274
rect 13222 694038 13306 694274
rect 13542 694038 32986 694274
rect 33222 694038 33306 694274
rect 33542 694038 52986 694274
rect 53222 694038 53306 694274
rect 53542 694038 72986 694274
rect 73222 694038 73306 694274
rect 73542 694038 92986 694274
rect 93222 694038 93306 694274
rect 93542 694038 112986 694274
rect 113222 694038 113306 694274
rect 113542 694038 132986 694274
rect 133222 694038 133306 694274
rect 133542 694038 152986 694274
rect 153222 694038 153306 694274
rect 153542 694038 172986 694274
rect 173222 694038 173306 694274
rect 173542 694038 192986 694274
rect 193222 694038 193306 694274
rect 193542 694038 212986 694274
rect 213222 694038 213306 694274
rect 213542 694038 232986 694274
rect 233222 694038 233306 694274
rect 233542 694038 252986 694274
rect 253222 694038 253306 694274
rect 253542 694038 272986 694274
rect 273222 694038 273306 694274
rect 273542 694038 292986 694274
rect 293222 694038 293306 694274
rect 293542 694038 312986 694274
rect 313222 694038 313306 694274
rect 313542 694038 332986 694274
rect 333222 694038 333306 694274
rect 333542 694038 352986 694274
rect 353222 694038 353306 694274
rect 353542 694038 372986 694274
rect 373222 694038 373306 694274
rect 373542 694038 392986 694274
rect 393222 694038 393306 694274
rect 393542 694038 412986 694274
rect 413222 694038 413306 694274
rect 413542 694038 432986 694274
rect 433222 694038 433306 694274
rect 433542 694038 452986 694274
rect 453222 694038 453306 694274
rect 453542 694038 472986 694274
rect 473222 694038 473306 694274
rect 473542 694038 492986 694274
rect 493222 694038 493306 694274
rect 493542 694038 512986 694274
rect 513222 694038 513306 694274
rect 513542 694038 532986 694274
rect 533222 694038 533306 694274
rect 533542 694038 552986 694274
rect 553222 694038 553306 694274
rect 553542 694038 572986 694274
rect 573222 694038 573306 694274
rect 573542 694038 591102 694274
rect 591338 694038 591422 694274
rect 591658 694038 592650 694274
rect -8726 693876 592650 694038
rect -2966 693294 586890 693456
rect -2966 693058 -2934 693294
rect -2698 693058 -2614 693294
rect -2378 693058 11826 693294
rect 12062 693058 12146 693294
rect 12382 693058 31826 693294
rect 32062 693058 32146 693294
rect 32382 693058 51826 693294
rect 52062 693058 52146 693294
rect 52382 693058 71826 693294
rect 72062 693058 72146 693294
rect 72382 693058 91826 693294
rect 92062 693058 92146 693294
rect 92382 693058 111826 693294
rect 112062 693058 112146 693294
rect 112382 693058 131826 693294
rect 132062 693058 132146 693294
rect 132382 693058 151826 693294
rect 152062 693058 152146 693294
rect 152382 693058 171826 693294
rect 172062 693058 172146 693294
rect 172382 693058 191826 693294
rect 192062 693058 192146 693294
rect 192382 693058 211826 693294
rect 212062 693058 212146 693294
rect 212382 693058 231826 693294
rect 232062 693058 232146 693294
rect 232382 693058 251826 693294
rect 252062 693058 252146 693294
rect 252382 693058 271826 693294
rect 272062 693058 272146 693294
rect 272382 693058 291826 693294
rect 292062 693058 292146 693294
rect 292382 693058 311826 693294
rect 312062 693058 312146 693294
rect 312382 693058 331826 693294
rect 332062 693058 332146 693294
rect 332382 693058 351826 693294
rect 352062 693058 352146 693294
rect 352382 693058 371826 693294
rect 372062 693058 372146 693294
rect 372382 693058 391826 693294
rect 392062 693058 392146 693294
rect 392382 693058 411826 693294
rect 412062 693058 412146 693294
rect 412382 693058 431826 693294
rect 432062 693058 432146 693294
rect 432382 693058 451826 693294
rect 452062 693058 452146 693294
rect 452382 693058 471826 693294
rect 472062 693058 472146 693294
rect 472382 693058 491826 693294
rect 492062 693058 492146 693294
rect 492382 693058 511826 693294
rect 512062 693058 512146 693294
rect 512382 693058 531826 693294
rect 532062 693058 532146 693294
rect 532382 693058 551826 693294
rect 552062 693058 552146 693294
rect 552382 693058 571826 693294
rect 572062 693058 572146 693294
rect 572382 693058 586302 693294
rect 586538 693058 586622 693294
rect 586858 693058 586890 693294
rect -2966 692896 586890 693058
rect -6806 690614 590730 690776
rect -6806 690378 -5814 690614
rect -5578 690378 -5494 690614
rect -5258 690378 9266 690614
rect 9502 690378 9586 690614
rect 9822 690378 29266 690614
rect 29502 690378 29586 690614
rect 29822 690378 49266 690614
rect 49502 690378 49586 690614
rect 49822 690378 69266 690614
rect 69502 690378 69586 690614
rect 69822 690378 89266 690614
rect 89502 690378 89586 690614
rect 89822 690378 109266 690614
rect 109502 690378 109586 690614
rect 109822 690378 129266 690614
rect 129502 690378 129586 690614
rect 129822 690378 149266 690614
rect 149502 690378 149586 690614
rect 149822 690378 169266 690614
rect 169502 690378 169586 690614
rect 169822 690378 189266 690614
rect 189502 690378 189586 690614
rect 189822 690378 209266 690614
rect 209502 690378 209586 690614
rect 209822 690378 229266 690614
rect 229502 690378 229586 690614
rect 229822 690378 249266 690614
rect 249502 690378 249586 690614
rect 249822 690378 269266 690614
rect 269502 690378 269586 690614
rect 269822 690378 289266 690614
rect 289502 690378 289586 690614
rect 289822 690378 309266 690614
rect 309502 690378 309586 690614
rect 309822 690378 329266 690614
rect 329502 690378 329586 690614
rect 329822 690378 349266 690614
rect 349502 690378 349586 690614
rect 349822 690378 369266 690614
rect 369502 690378 369586 690614
rect 369822 690378 389266 690614
rect 389502 690378 389586 690614
rect 389822 690378 409266 690614
rect 409502 690378 409586 690614
rect 409822 690378 429266 690614
rect 429502 690378 429586 690614
rect 429822 690378 449266 690614
rect 449502 690378 449586 690614
rect 449822 690378 469266 690614
rect 469502 690378 469586 690614
rect 469822 690378 489266 690614
rect 489502 690378 489586 690614
rect 489822 690378 509266 690614
rect 509502 690378 509586 690614
rect 509822 690378 529266 690614
rect 529502 690378 529586 690614
rect 529822 690378 549266 690614
rect 549502 690378 549586 690614
rect 549822 690378 569266 690614
rect 569502 690378 569586 690614
rect 569822 690378 589182 690614
rect 589418 690378 589502 690614
rect 589738 690378 590730 690614
rect -6806 690216 590730 690378
rect -4886 686954 588810 687116
rect -4886 686718 -3894 686954
rect -3658 686718 -3574 686954
rect -3338 686718 5546 686954
rect 5782 686718 5866 686954
rect 6102 686718 25546 686954
rect 25782 686718 25866 686954
rect 26102 686718 45546 686954
rect 45782 686718 45866 686954
rect 46102 686718 65546 686954
rect 65782 686718 65866 686954
rect 66102 686718 85546 686954
rect 85782 686718 85866 686954
rect 86102 686718 105546 686954
rect 105782 686718 105866 686954
rect 106102 686718 125546 686954
rect 125782 686718 125866 686954
rect 126102 686718 145546 686954
rect 145782 686718 145866 686954
rect 146102 686718 165546 686954
rect 165782 686718 165866 686954
rect 166102 686718 185546 686954
rect 185782 686718 185866 686954
rect 186102 686718 205546 686954
rect 205782 686718 205866 686954
rect 206102 686718 225546 686954
rect 225782 686718 225866 686954
rect 226102 686718 245546 686954
rect 245782 686718 245866 686954
rect 246102 686718 265546 686954
rect 265782 686718 265866 686954
rect 266102 686718 285546 686954
rect 285782 686718 285866 686954
rect 286102 686718 305546 686954
rect 305782 686718 305866 686954
rect 306102 686718 325546 686954
rect 325782 686718 325866 686954
rect 326102 686718 345546 686954
rect 345782 686718 345866 686954
rect 346102 686718 365546 686954
rect 365782 686718 365866 686954
rect 366102 686718 385546 686954
rect 385782 686718 385866 686954
rect 386102 686718 405546 686954
rect 405782 686718 405866 686954
rect 406102 686718 425546 686954
rect 425782 686718 425866 686954
rect 426102 686718 445546 686954
rect 445782 686718 445866 686954
rect 446102 686718 465546 686954
rect 465782 686718 465866 686954
rect 466102 686718 485546 686954
rect 485782 686718 485866 686954
rect 486102 686718 505546 686954
rect 505782 686718 505866 686954
rect 506102 686718 525546 686954
rect 525782 686718 525866 686954
rect 526102 686718 545546 686954
rect 545782 686718 545866 686954
rect 546102 686718 565546 686954
rect 565782 686718 565866 686954
rect 566102 686718 587262 686954
rect 587498 686718 587582 686954
rect 587818 686718 588810 686954
rect -4886 686556 588810 686718
rect -8726 684274 592650 684436
rect -8726 684038 -8694 684274
rect -8458 684038 -8374 684274
rect -8138 684038 22986 684274
rect 23222 684038 23306 684274
rect 23542 684038 42986 684274
rect 43222 684038 43306 684274
rect 43542 684038 62986 684274
rect 63222 684038 63306 684274
rect 63542 684038 82986 684274
rect 83222 684038 83306 684274
rect 83542 684038 102986 684274
rect 103222 684038 103306 684274
rect 103542 684038 122986 684274
rect 123222 684038 123306 684274
rect 123542 684038 142986 684274
rect 143222 684038 143306 684274
rect 143542 684038 162986 684274
rect 163222 684038 163306 684274
rect 163542 684038 182986 684274
rect 183222 684038 183306 684274
rect 183542 684038 202986 684274
rect 203222 684038 203306 684274
rect 203542 684038 222986 684274
rect 223222 684038 223306 684274
rect 223542 684038 242986 684274
rect 243222 684038 243306 684274
rect 243542 684038 262986 684274
rect 263222 684038 263306 684274
rect 263542 684038 282986 684274
rect 283222 684038 283306 684274
rect 283542 684038 302986 684274
rect 303222 684038 303306 684274
rect 303542 684038 322986 684274
rect 323222 684038 323306 684274
rect 323542 684038 342986 684274
rect 343222 684038 343306 684274
rect 343542 684038 362986 684274
rect 363222 684038 363306 684274
rect 363542 684038 382986 684274
rect 383222 684038 383306 684274
rect 383542 684038 402986 684274
rect 403222 684038 403306 684274
rect 403542 684038 422986 684274
rect 423222 684038 423306 684274
rect 423542 684038 442986 684274
rect 443222 684038 443306 684274
rect 443542 684038 462986 684274
rect 463222 684038 463306 684274
rect 463542 684038 482986 684274
rect 483222 684038 483306 684274
rect 483542 684038 502986 684274
rect 503222 684038 503306 684274
rect 503542 684038 522986 684274
rect 523222 684038 523306 684274
rect 523542 684038 542986 684274
rect 543222 684038 543306 684274
rect 543542 684038 562986 684274
rect 563222 684038 563306 684274
rect 563542 684038 592062 684274
rect 592298 684038 592382 684274
rect 592618 684038 592650 684274
rect -8726 683876 592650 684038
rect -2966 683294 586890 683456
rect -2966 683058 -1974 683294
rect -1738 683058 -1654 683294
rect -1418 683058 1826 683294
rect 2062 683058 2146 683294
rect 2382 683058 21826 683294
rect 22062 683058 22146 683294
rect 22382 683058 41826 683294
rect 42062 683058 42146 683294
rect 42382 683058 61826 683294
rect 62062 683058 62146 683294
rect 62382 683058 81826 683294
rect 82062 683058 82146 683294
rect 82382 683058 101826 683294
rect 102062 683058 102146 683294
rect 102382 683058 121826 683294
rect 122062 683058 122146 683294
rect 122382 683058 141826 683294
rect 142062 683058 142146 683294
rect 142382 683058 161826 683294
rect 162062 683058 162146 683294
rect 162382 683058 181826 683294
rect 182062 683058 182146 683294
rect 182382 683058 201826 683294
rect 202062 683058 202146 683294
rect 202382 683058 221826 683294
rect 222062 683058 222146 683294
rect 222382 683058 241826 683294
rect 242062 683058 242146 683294
rect 242382 683058 261826 683294
rect 262062 683058 262146 683294
rect 262382 683058 281826 683294
rect 282062 683058 282146 683294
rect 282382 683058 301826 683294
rect 302062 683058 302146 683294
rect 302382 683058 321826 683294
rect 322062 683058 322146 683294
rect 322382 683058 341826 683294
rect 342062 683058 342146 683294
rect 342382 683058 361826 683294
rect 362062 683058 362146 683294
rect 362382 683058 381826 683294
rect 382062 683058 382146 683294
rect 382382 683058 401826 683294
rect 402062 683058 402146 683294
rect 402382 683058 421826 683294
rect 422062 683058 422146 683294
rect 422382 683058 441826 683294
rect 442062 683058 442146 683294
rect 442382 683058 461826 683294
rect 462062 683058 462146 683294
rect 462382 683058 481826 683294
rect 482062 683058 482146 683294
rect 482382 683058 501826 683294
rect 502062 683058 502146 683294
rect 502382 683058 521826 683294
rect 522062 683058 522146 683294
rect 522382 683058 541826 683294
rect 542062 683058 542146 683294
rect 542382 683058 561826 683294
rect 562062 683058 562146 683294
rect 562382 683058 581826 683294
rect 582062 683058 582146 683294
rect 582382 683058 585342 683294
rect 585578 683058 585662 683294
rect 585898 683058 586890 683294
rect -2966 682896 586890 683058
rect -6806 680614 590730 680776
rect -6806 680378 -6774 680614
rect -6538 680378 -6454 680614
rect -6218 680378 19266 680614
rect 19502 680378 19586 680614
rect 19822 680378 39266 680614
rect 39502 680378 39586 680614
rect 39822 680378 59266 680614
rect 59502 680378 59586 680614
rect 59822 680378 79266 680614
rect 79502 680378 79586 680614
rect 79822 680378 99266 680614
rect 99502 680378 99586 680614
rect 99822 680378 119266 680614
rect 119502 680378 119586 680614
rect 119822 680378 139266 680614
rect 139502 680378 139586 680614
rect 139822 680378 159266 680614
rect 159502 680378 159586 680614
rect 159822 680378 179266 680614
rect 179502 680378 179586 680614
rect 179822 680378 199266 680614
rect 199502 680378 199586 680614
rect 199822 680378 219266 680614
rect 219502 680378 219586 680614
rect 219822 680378 239266 680614
rect 239502 680378 239586 680614
rect 239822 680378 259266 680614
rect 259502 680378 259586 680614
rect 259822 680378 279266 680614
rect 279502 680378 279586 680614
rect 279822 680378 299266 680614
rect 299502 680378 299586 680614
rect 299822 680378 319266 680614
rect 319502 680378 319586 680614
rect 319822 680378 339266 680614
rect 339502 680378 339586 680614
rect 339822 680378 359266 680614
rect 359502 680378 359586 680614
rect 359822 680378 379266 680614
rect 379502 680378 379586 680614
rect 379822 680378 399266 680614
rect 399502 680378 399586 680614
rect 399822 680378 419266 680614
rect 419502 680378 419586 680614
rect 419822 680378 439266 680614
rect 439502 680378 439586 680614
rect 439822 680378 459266 680614
rect 459502 680378 459586 680614
rect 459822 680378 479266 680614
rect 479502 680378 479586 680614
rect 479822 680378 499266 680614
rect 499502 680378 499586 680614
rect 499822 680378 519266 680614
rect 519502 680378 519586 680614
rect 519822 680378 539266 680614
rect 539502 680378 539586 680614
rect 539822 680378 559266 680614
rect 559502 680378 559586 680614
rect 559822 680378 579266 680614
rect 579502 680378 579586 680614
rect 579822 680378 590142 680614
rect 590378 680378 590462 680614
rect 590698 680378 590730 680614
rect -6806 680216 590730 680378
rect -4886 676954 588810 677116
rect -4886 676718 -4854 676954
rect -4618 676718 -4534 676954
rect -4298 676718 15546 676954
rect 15782 676718 15866 676954
rect 16102 676718 35546 676954
rect 35782 676718 35866 676954
rect 36102 676718 55546 676954
rect 55782 676718 55866 676954
rect 56102 676718 75546 676954
rect 75782 676718 75866 676954
rect 76102 676718 95546 676954
rect 95782 676718 95866 676954
rect 96102 676718 115546 676954
rect 115782 676718 115866 676954
rect 116102 676718 135546 676954
rect 135782 676718 135866 676954
rect 136102 676718 155546 676954
rect 155782 676718 155866 676954
rect 156102 676718 175546 676954
rect 175782 676718 175866 676954
rect 176102 676718 195546 676954
rect 195782 676718 195866 676954
rect 196102 676718 215546 676954
rect 215782 676718 215866 676954
rect 216102 676718 235546 676954
rect 235782 676718 235866 676954
rect 236102 676718 255546 676954
rect 255782 676718 255866 676954
rect 256102 676718 275546 676954
rect 275782 676718 275866 676954
rect 276102 676718 295546 676954
rect 295782 676718 295866 676954
rect 296102 676718 315546 676954
rect 315782 676718 315866 676954
rect 316102 676718 335546 676954
rect 335782 676718 335866 676954
rect 336102 676718 355546 676954
rect 355782 676718 355866 676954
rect 356102 676718 375546 676954
rect 375782 676718 375866 676954
rect 376102 676718 395546 676954
rect 395782 676718 395866 676954
rect 396102 676718 415546 676954
rect 415782 676718 415866 676954
rect 416102 676718 435546 676954
rect 435782 676718 435866 676954
rect 436102 676718 455546 676954
rect 455782 676718 455866 676954
rect 456102 676718 475546 676954
rect 475782 676718 475866 676954
rect 476102 676718 495546 676954
rect 495782 676718 495866 676954
rect 496102 676718 515546 676954
rect 515782 676718 515866 676954
rect 516102 676718 535546 676954
rect 535782 676718 535866 676954
rect 536102 676718 555546 676954
rect 555782 676718 555866 676954
rect 556102 676718 575546 676954
rect 575782 676718 575866 676954
rect 576102 676718 588222 676954
rect 588458 676718 588542 676954
rect 588778 676718 588810 676954
rect -4886 676556 588810 676718
rect -8726 674274 592650 674436
rect -8726 674038 -7734 674274
rect -7498 674038 -7414 674274
rect -7178 674038 12986 674274
rect 13222 674038 13306 674274
rect 13542 674038 172986 674274
rect 173222 674038 173306 674274
rect 173542 674038 192986 674274
rect 193222 674038 193306 674274
rect 193542 674038 212986 674274
rect 213222 674038 213306 674274
rect 213542 674038 232986 674274
rect 233222 674038 233306 674274
rect 233542 674038 252986 674274
rect 253222 674038 253306 674274
rect 253542 674038 272986 674274
rect 273222 674038 273306 674274
rect 273542 674038 292986 674274
rect 293222 674038 293306 674274
rect 293542 674038 312986 674274
rect 313222 674038 313306 674274
rect 313542 674038 332986 674274
rect 333222 674038 333306 674274
rect 333542 674038 352986 674274
rect 353222 674038 353306 674274
rect 353542 674038 372986 674274
rect 373222 674038 373306 674274
rect 373542 674038 392986 674274
rect 393222 674038 393306 674274
rect 393542 674038 412986 674274
rect 413222 674038 413306 674274
rect 413542 674038 432986 674274
rect 433222 674038 433306 674274
rect 433542 674038 452986 674274
rect 453222 674038 453306 674274
rect 453542 674038 472986 674274
rect 473222 674038 473306 674274
rect 473542 674038 492986 674274
rect 493222 674038 493306 674274
rect 493542 674038 512986 674274
rect 513222 674038 513306 674274
rect 513542 674038 532986 674274
rect 533222 674038 533306 674274
rect 533542 674038 552986 674274
rect 553222 674038 553306 674274
rect 553542 674038 572986 674274
rect 573222 674038 573306 674274
rect 573542 674038 591102 674274
rect 591338 674038 591422 674274
rect 591658 674038 592650 674274
rect -8726 673876 592650 674038
rect -2966 673294 586890 673456
rect -2966 673058 -2934 673294
rect -2698 673058 -2614 673294
rect -2378 673058 11826 673294
rect 12062 673058 12146 673294
rect 12382 673058 171826 673294
rect 172062 673058 172146 673294
rect 172382 673058 191826 673294
rect 192062 673058 192146 673294
rect 192382 673058 211826 673294
rect 212062 673058 212146 673294
rect 212382 673058 231826 673294
rect 232062 673058 232146 673294
rect 232382 673058 251826 673294
rect 252062 673058 252146 673294
rect 252382 673058 271826 673294
rect 272062 673058 272146 673294
rect 272382 673058 291826 673294
rect 292062 673058 292146 673294
rect 292382 673058 311826 673294
rect 312062 673058 312146 673294
rect 312382 673058 331826 673294
rect 332062 673058 332146 673294
rect 332382 673058 351826 673294
rect 352062 673058 352146 673294
rect 352382 673058 371826 673294
rect 372062 673058 372146 673294
rect 372382 673058 391826 673294
rect 392062 673058 392146 673294
rect 392382 673058 411826 673294
rect 412062 673058 412146 673294
rect 412382 673058 431826 673294
rect 432062 673058 432146 673294
rect 432382 673058 451826 673294
rect 452062 673058 452146 673294
rect 452382 673058 471826 673294
rect 472062 673058 472146 673294
rect 472382 673058 491826 673294
rect 492062 673058 492146 673294
rect 492382 673058 511826 673294
rect 512062 673058 512146 673294
rect 512382 673058 531826 673294
rect 532062 673058 532146 673294
rect 532382 673058 551826 673294
rect 552062 673058 552146 673294
rect 552382 673058 571826 673294
rect 572062 673058 572146 673294
rect 572382 673058 586302 673294
rect 586538 673058 586622 673294
rect 586858 673058 586890 673294
rect -2966 672896 586890 673058
rect -6806 670614 590730 670776
rect -6806 670378 -5814 670614
rect -5578 670378 -5494 670614
rect -5258 670378 9266 670614
rect 9502 670378 9586 670614
rect 9822 670378 169266 670614
rect 169502 670378 169586 670614
rect 169822 670378 189266 670614
rect 189502 670378 189586 670614
rect 189822 670378 209266 670614
rect 209502 670378 209586 670614
rect 209822 670378 229266 670614
rect 229502 670378 229586 670614
rect 229822 670378 249266 670614
rect 249502 670378 249586 670614
rect 249822 670378 269266 670614
rect 269502 670378 269586 670614
rect 269822 670378 289266 670614
rect 289502 670378 289586 670614
rect 289822 670378 309266 670614
rect 309502 670378 309586 670614
rect 309822 670378 329266 670614
rect 329502 670378 329586 670614
rect 329822 670378 349266 670614
rect 349502 670378 349586 670614
rect 349822 670378 369266 670614
rect 369502 670378 369586 670614
rect 369822 670378 389266 670614
rect 389502 670378 389586 670614
rect 389822 670378 409266 670614
rect 409502 670378 409586 670614
rect 409822 670378 429266 670614
rect 429502 670378 429586 670614
rect 429822 670378 449266 670614
rect 449502 670378 449586 670614
rect 449822 670378 469266 670614
rect 469502 670378 469586 670614
rect 469822 670378 489266 670614
rect 489502 670378 489586 670614
rect 489822 670378 509266 670614
rect 509502 670378 509586 670614
rect 509822 670378 529266 670614
rect 529502 670378 529586 670614
rect 529822 670378 549266 670614
rect 549502 670378 549586 670614
rect 549822 670378 569266 670614
rect 569502 670378 569586 670614
rect 569822 670378 589182 670614
rect 589418 670378 589502 670614
rect 589738 670378 590730 670614
rect -6806 670216 590730 670378
rect -4886 666954 588810 667116
rect -4886 666718 -3894 666954
rect -3658 666718 -3574 666954
rect -3338 666718 5546 666954
rect 5782 666718 5866 666954
rect 6102 666718 25546 666954
rect 25782 666718 25866 666954
rect 26102 666718 185546 666954
rect 185782 666718 185866 666954
rect 186102 666718 205546 666954
rect 205782 666718 205866 666954
rect 206102 666718 225546 666954
rect 225782 666718 225866 666954
rect 226102 666718 245546 666954
rect 245782 666718 245866 666954
rect 246102 666718 265546 666954
rect 265782 666718 265866 666954
rect 266102 666718 285546 666954
rect 285782 666718 285866 666954
rect 286102 666718 305546 666954
rect 305782 666718 305866 666954
rect 306102 666718 325546 666954
rect 325782 666718 325866 666954
rect 326102 666718 345546 666954
rect 345782 666718 345866 666954
rect 346102 666718 365546 666954
rect 365782 666718 365866 666954
rect 366102 666718 385546 666954
rect 385782 666718 385866 666954
rect 386102 666718 405546 666954
rect 405782 666718 405866 666954
rect 406102 666718 425546 666954
rect 425782 666718 425866 666954
rect 426102 666718 445546 666954
rect 445782 666718 445866 666954
rect 446102 666718 465546 666954
rect 465782 666718 465866 666954
rect 466102 666718 485546 666954
rect 485782 666718 485866 666954
rect 486102 666718 505546 666954
rect 505782 666718 505866 666954
rect 506102 666718 525546 666954
rect 525782 666718 525866 666954
rect 526102 666718 545546 666954
rect 545782 666718 545866 666954
rect 546102 666718 565546 666954
rect 565782 666718 565866 666954
rect 566102 666718 587262 666954
rect 587498 666718 587582 666954
rect 587818 666718 588810 666954
rect -4886 666556 588810 666718
rect -8726 664274 592650 664436
rect -8726 664038 -8694 664274
rect -8458 664038 -8374 664274
rect -8138 664038 22986 664274
rect 23222 664038 23306 664274
rect 23542 664038 182986 664274
rect 183222 664038 183306 664274
rect 183542 664038 202986 664274
rect 203222 664038 203306 664274
rect 203542 664038 222986 664274
rect 223222 664038 223306 664274
rect 223542 664038 242986 664274
rect 243222 664038 243306 664274
rect 243542 664038 262986 664274
rect 263222 664038 263306 664274
rect 263542 664038 282986 664274
rect 283222 664038 283306 664274
rect 283542 664038 302986 664274
rect 303222 664038 303306 664274
rect 303542 664038 322986 664274
rect 323222 664038 323306 664274
rect 323542 664038 342986 664274
rect 343222 664038 343306 664274
rect 343542 664038 362986 664274
rect 363222 664038 363306 664274
rect 363542 664038 382986 664274
rect 383222 664038 383306 664274
rect 383542 664038 402986 664274
rect 403222 664038 403306 664274
rect 403542 664038 422986 664274
rect 423222 664038 423306 664274
rect 423542 664038 442986 664274
rect 443222 664038 443306 664274
rect 443542 664038 462986 664274
rect 463222 664038 463306 664274
rect 463542 664038 482986 664274
rect 483222 664038 483306 664274
rect 483542 664038 502986 664274
rect 503222 664038 503306 664274
rect 503542 664038 522986 664274
rect 523222 664038 523306 664274
rect 523542 664038 542986 664274
rect 543222 664038 543306 664274
rect 543542 664038 562986 664274
rect 563222 664038 563306 664274
rect 563542 664038 592062 664274
rect 592298 664038 592382 664274
rect 592618 664038 592650 664274
rect -8726 663876 592650 664038
rect -2966 663294 586890 663456
rect -2966 663058 -1974 663294
rect -1738 663058 -1654 663294
rect -1418 663058 1826 663294
rect 2062 663058 2146 663294
rect 2382 663058 21826 663294
rect 22062 663058 22146 663294
rect 22382 663058 31008 663294
rect 31244 663058 165376 663294
rect 165612 663058 181826 663294
rect 182062 663058 182146 663294
rect 182382 663058 201826 663294
rect 202062 663058 202146 663294
rect 202382 663058 221826 663294
rect 222062 663058 222146 663294
rect 222382 663058 241826 663294
rect 242062 663058 242146 663294
rect 242382 663058 261826 663294
rect 262062 663058 262146 663294
rect 262382 663058 281826 663294
rect 282062 663058 282146 663294
rect 282382 663058 301826 663294
rect 302062 663058 302146 663294
rect 302382 663058 321826 663294
rect 322062 663058 322146 663294
rect 322382 663058 341826 663294
rect 342062 663058 342146 663294
rect 342382 663058 361826 663294
rect 362062 663058 362146 663294
rect 362382 663058 381826 663294
rect 382062 663058 382146 663294
rect 382382 663058 401826 663294
rect 402062 663058 402146 663294
rect 402382 663058 421826 663294
rect 422062 663058 422146 663294
rect 422382 663058 441826 663294
rect 442062 663058 442146 663294
rect 442382 663058 461826 663294
rect 462062 663058 462146 663294
rect 462382 663058 481826 663294
rect 482062 663058 482146 663294
rect 482382 663058 501826 663294
rect 502062 663058 502146 663294
rect 502382 663058 521826 663294
rect 522062 663058 522146 663294
rect 522382 663058 541826 663294
rect 542062 663058 542146 663294
rect 542382 663058 561826 663294
rect 562062 663058 562146 663294
rect 562382 663058 581826 663294
rect 582062 663058 582146 663294
rect 582382 663058 585342 663294
rect 585578 663058 585662 663294
rect 585898 663058 586890 663294
rect -2966 662896 586890 663058
rect -6806 660614 590730 660776
rect -6806 660378 -6774 660614
rect -6538 660378 -6454 660614
rect -6218 660378 19266 660614
rect 19502 660378 19586 660614
rect 19822 660378 179266 660614
rect 179502 660378 179586 660614
rect 179822 660378 199266 660614
rect 199502 660378 199586 660614
rect 199822 660378 219266 660614
rect 219502 660378 219586 660614
rect 219822 660378 239266 660614
rect 239502 660378 239586 660614
rect 239822 660378 259266 660614
rect 259502 660378 259586 660614
rect 259822 660378 279266 660614
rect 279502 660378 279586 660614
rect 279822 660378 299266 660614
rect 299502 660378 299586 660614
rect 299822 660378 319266 660614
rect 319502 660378 319586 660614
rect 319822 660378 339266 660614
rect 339502 660378 339586 660614
rect 339822 660378 359266 660614
rect 359502 660378 359586 660614
rect 359822 660378 379266 660614
rect 379502 660378 379586 660614
rect 379822 660378 399266 660614
rect 399502 660378 399586 660614
rect 399822 660378 419266 660614
rect 419502 660378 419586 660614
rect 419822 660378 439266 660614
rect 439502 660378 439586 660614
rect 439822 660378 459266 660614
rect 459502 660378 459586 660614
rect 459822 660378 479266 660614
rect 479502 660378 479586 660614
rect 479822 660378 499266 660614
rect 499502 660378 499586 660614
rect 499822 660378 519266 660614
rect 519502 660378 519586 660614
rect 519822 660378 539266 660614
rect 539502 660378 539586 660614
rect 539822 660378 559266 660614
rect 559502 660378 559586 660614
rect 559822 660378 579266 660614
rect 579502 660378 579586 660614
rect 579822 660378 590142 660614
rect 590378 660378 590462 660614
rect 590698 660378 590730 660614
rect -6806 660216 590730 660378
rect -4886 656954 588810 657116
rect -4886 656718 -4854 656954
rect -4618 656718 -4534 656954
rect -4298 656718 15546 656954
rect 15782 656718 15866 656954
rect 16102 656718 175546 656954
rect 175782 656718 175866 656954
rect 176102 656718 195546 656954
rect 195782 656718 195866 656954
rect 196102 656718 215546 656954
rect 215782 656718 215866 656954
rect 216102 656718 235546 656954
rect 235782 656718 235866 656954
rect 236102 656718 355546 656954
rect 355782 656718 355866 656954
rect 356102 656718 375546 656954
rect 375782 656718 375866 656954
rect 376102 656718 395546 656954
rect 395782 656718 395866 656954
rect 396102 656718 515546 656954
rect 515782 656718 515866 656954
rect 516102 656718 535546 656954
rect 535782 656718 535866 656954
rect 536102 656718 555546 656954
rect 555782 656718 555866 656954
rect 556102 656718 575546 656954
rect 575782 656718 575866 656954
rect 576102 656718 588222 656954
rect 588458 656718 588542 656954
rect 588778 656718 588810 656954
rect -4886 656556 588810 656718
rect -8726 654274 592650 654436
rect -8726 654038 -7734 654274
rect -7498 654038 -7414 654274
rect -7178 654038 12986 654274
rect 13222 654038 13306 654274
rect 13542 654038 172986 654274
rect 173222 654038 173306 654274
rect 173542 654038 192986 654274
rect 193222 654038 193306 654274
rect 193542 654038 212986 654274
rect 213222 654038 213306 654274
rect 213542 654038 232986 654274
rect 233222 654038 233306 654274
rect 233542 654038 352986 654274
rect 353222 654038 353306 654274
rect 353542 654038 372986 654274
rect 373222 654038 373306 654274
rect 373542 654038 392986 654274
rect 393222 654038 393306 654274
rect 393542 654038 512986 654274
rect 513222 654038 513306 654274
rect 513542 654038 532986 654274
rect 533222 654038 533306 654274
rect 533542 654038 552986 654274
rect 553222 654038 553306 654274
rect 553542 654038 572986 654274
rect 573222 654038 573306 654274
rect 573542 654038 591102 654274
rect 591338 654038 591422 654274
rect 591658 654038 592650 654274
rect -8726 653876 592650 654038
rect -2966 653294 586890 653456
rect -2966 653058 -2934 653294
rect -2698 653058 -2614 653294
rect -2378 653058 11826 653294
rect 12062 653058 12146 653294
rect 12382 653058 30328 653294
rect 30564 653058 166056 653294
rect 166292 653058 171826 653294
rect 172062 653058 172146 653294
rect 172382 653058 191826 653294
rect 192062 653058 192146 653294
rect 192382 653058 211826 653294
rect 212062 653058 212146 653294
rect 212382 653058 231826 653294
rect 232062 653058 232146 653294
rect 232382 653058 240328 653294
rect 240564 653058 335392 653294
rect 335628 653058 351826 653294
rect 352062 653058 352146 653294
rect 352382 653058 371826 653294
rect 372062 653058 372146 653294
rect 372382 653058 391826 653294
rect 392062 653058 392146 653294
rect 392382 653058 410328 653294
rect 410564 653058 505392 653294
rect 505628 653058 511826 653294
rect 512062 653058 512146 653294
rect 512382 653058 531826 653294
rect 532062 653058 532146 653294
rect 532382 653058 551826 653294
rect 552062 653058 552146 653294
rect 552382 653058 571826 653294
rect 572062 653058 572146 653294
rect 572382 653058 586302 653294
rect 586538 653058 586622 653294
rect 586858 653058 586890 653294
rect -2966 652896 586890 653058
rect -6806 650614 590730 650776
rect -6806 650378 -5814 650614
rect -5578 650378 -5494 650614
rect -5258 650378 9266 650614
rect 9502 650378 9586 650614
rect 9822 650378 169266 650614
rect 169502 650378 169586 650614
rect 169822 650378 189266 650614
rect 189502 650378 189586 650614
rect 189822 650378 209266 650614
rect 209502 650378 209586 650614
rect 209822 650378 229266 650614
rect 229502 650378 229586 650614
rect 229822 650378 349266 650614
rect 349502 650378 349586 650614
rect 349822 650378 369266 650614
rect 369502 650378 369586 650614
rect 369822 650378 389266 650614
rect 389502 650378 389586 650614
rect 389822 650378 509266 650614
rect 509502 650378 509586 650614
rect 509822 650378 529266 650614
rect 529502 650378 529586 650614
rect 529822 650378 549266 650614
rect 549502 650378 549586 650614
rect 549822 650378 569266 650614
rect 569502 650378 569586 650614
rect 569822 650378 589182 650614
rect 589418 650378 589502 650614
rect 589738 650378 590730 650614
rect -6806 650216 590730 650378
rect -4886 646954 588810 647116
rect -4886 646718 -3894 646954
rect -3658 646718 -3574 646954
rect -3338 646718 5546 646954
rect 5782 646718 5866 646954
rect 6102 646718 25546 646954
rect 25782 646718 25866 646954
rect 26102 646718 185546 646954
rect 185782 646718 185866 646954
rect 186102 646718 205546 646954
rect 205782 646718 205866 646954
rect 206102 646718 225546 646954
rect 225782 646718 225866 646954
rect 226102 646718 345546 646954
rect 345782 646718 345866 646954
rect 346102 646718 365546 646954
rect 365782 646718 365866 646954
rect 366102 646718 385546 646954
rect 385782 646718 385866 646954
rect 386102 646718 405546 646954
rect 405782 646718 405866 646954
rect 406102 646718 525546 646954
rect 525782 646718 525866 646954
rect 526102 646718 545546 646954
rect 545782 646718 545866 646954
rect 546102 646718 565546 646954
rect 565782 646718 565866 646954
rect 566102 646718 587262 646954
rect 587498 646718 587582 646954
rect 587818 646718 588810 646954
rect -4886 646556 588810 646718
rect -8726 644274 592650 644436
rect -8726 644038 -8694 644274
rect -8458 644038 -8374 644274
rect -8138 644038 22986 644274
rect 23222 644038 23306 644274
rect 23542 644038 182986 644274
rect 183222 644038 183306 644274
rect 183542 644038 202986 644274
rect 203222 644038 203306 644274
rect 203542 644038 222986 644274
rect 223222 644038 223306 644274
rect 223542 644038 342986 644274
rect 343222 644038 343306 644274
rect 343542 644038 362986 644274
rect 363222 644038 363306 644274
rect 363542 644038 382986 644274
rect 383222 644038 383306 644274
rect 383542 644038 402986 644274
rect 403222 644038 403306 644274
rect 403542 644038 522986 644274
rect 523222 644038 523306 644274
rect 523542 644038 542986 644274
rect 543222 644038 543306 644274
rect 543542 644038 562986 644274
rect 563222 644038 563306 644274
rect 563542 644038 592062 644274
rect 592298 644038 592382 644274
rect 592618 644038 592650 644274
rect -8726 643876 592650 644038
rect -2966 643294 586890 643456
rect -2966 643058 -1974 643294
rect -1738 643058 -1654 643294
rect -1418 643058 1826 643294
rect 2062 643058 2146 643294
rect 2382 643058 21826 643294
rect 22062 643058 22146 643294
rect 22382 643058 31008 643294
rect 31244 643058 165376 643294
rect 165612 643058 181826 643294
rect 182062 643058 182146 643294
rect 182382 643058 201826 643294
rect 202062 643058 202146 643294
rect 202382 643058 221826 643294
rect 222062 643058 222146 643294
rect 222382 643058 241008 643294
rect 241244 643058 334712 643294
rect 334948 643058 341826 643294
rect 342062 643058 342146 643294
rect 342382 643058 361826 643294
rect 362062 643058 362146 643294
rect 362382 643058 381826 643294
rect 382062 643058 382146 643294
rect 382382 643058 401826 643294
rect 402062 643058 402146 643294
rect 402382 643058 411008 643294
rect 411244 643058 504712 643294
rect 504948 643058 521826 643294
rect 522062 643058 522146 643294
rect 522382 643058 541826 643294
rect 542062 643058 542146 643294
rect 542382 643058 561826 643294
rect 562062 643058 562146 643294
rect 562382 643058 581826 643294
rect 582062 643058 582146 643294
rect 582382 643058 585342 643294
rect 585578 643058 585662 643294
rect 585898 643058 586890 643294
rect -2966 642896 586890 643058
rect -6806 640614 590730 640776
rect -6806 640378 -6774 640614
rect -6538 640378 -6454 640614
rect -6218 640378 19266 640614
rect 19502 640378 19586 640614
rect 19822 640378 179266 640614
rect 179502 640378 179586 640614
rect 179822 640378 199266 640614
rect 199502 640378 199586 640614
rect 199822 640378 219266 640614
rect 219502 640378 219586 640614
rect 219822 640378 339266 640614
rect 339502 640378 339586 640614
rect 339822 640378 359266 640614
rect 359502 640378 359586 640614
rect 359822 640378 379266 640614
rect 379502 640378 379586 640614
rect 379822 640378 399266 640614
rect 399502 640378 399586 640614
rect 399822 640378 519266 640614
rect 519502 640378 519586 640614
rect 519822 640378 539266 640614
rect 539502 640378 539586 640614
rect 539822 640378 559266 640614
rect 559502 640378 559586 640614
rect 559822 640378 579266 640614
rect 579502 640378 579586 640614
rect 579822 640378 590142 640614
rect 590378 640378 590462 640614
rect 590698 640378 590730 640614
rect -6806 640216 590730 640378
rect -4886 636954 588810 637116
rect -4886 636718 -4854 636954
rect -4618 636718 -4534 636954
rect -4298 636718 15546 636954
rect 15782 636718 15866 636954
rect 16102 636718 175546 636954
rect 175782 636718 175866 636954
rect 176102 636718 195546 636954
rect 195782 636718 195866 636954
rect 196102 636718 215546 636954
rect 215782 636718 215866 636954
rect 216102 636718 235546 636954
rect 235782 636718 235866 636954
rect 236102 636718 355546 636954
rect 355782 636718 355866 636954
rect 356102 636718 375546 636954
rect 375782 636718 375866 636954
rect 376102 636718 395546 636954
rect 395782 636718 395866 636954
rect 396102 636718 515546 636954
rect 515782 636718 515866 636954
rect 516102 636718 535546 636954
rect 535782 636718 535866 636954
rect 536102 636718 555546 636954
rect 555782 636718 555866 636954
rect 556102 636718 575546 636954
rect 575782 636718 575866 636954
rect 576102 636718 588222 636954
rect 588458 636718 588542 636954
rect 588778 636718 588810 636954
rect -4886 636556 588810 636718
rect -8726 634274 592650 634436
rect -8726 634038 -7734 634274
rect -7498 634038 -7414 634274
rect -7178 634038 12986 634274
rect 13222 634038 13306 634274
rect 13542 634038 172986 634274
rect 173222 634038 173306 634274
rect 173542 634038 192986 634274
rect 193222 634038 193306 634274
rect 193542 634038 212986 634274
rect 213222 634038 213306 634274
rect 213542 634038 232986 634274
rect 233222 634038 233306 634274
rect 233542 634038 352986 634274
rect 353222 634038 353306 634274
rect 353542 634038 372986 634274
rect 373222 634038 373306 634274
rect 373542 634038 392986 634274
rect 393222 634038 393306 634274
rect 393542 634038 512986 634274
rect 513222 634038 513306 634274
rect 513542 634038 532986 634274
rect 533222 634038 533306 634274
rect 533542 634038 552986 634274
rect 553222 634038 553306 634274
rect 553542 634038 572986 634274
rect 573222 634038 573306 634274
rect 573542 634038 591102 634274
rect 591338 634038 591422 634274
rect 591658 634038 592650 634274
rect -8726 633876 592650 634038
rect -2966 633294 586890 633456
rect -2966 633058 -2934 633294
rect -2698 633058 -2614 633294
rect -2378 633058 11826 633294
rect 12062 633058 12146 633294
rect 12382 633058 30328 633294
rect 30564 633058 166056 633294
rect 166292 633058 171826 633294
rect 172062 633058 172146 633294
rect 172382 633058 191826 633294
rect 192062 633058 192146 633294
rect 192382 633058 211826 633294
rect 212062 633058 212146 633294
rect 212382 633058 231826 633294
rect 232062 633058 232146 633294
rect 232382 633058 240328 633294
rect 240564 633058 335392 633294
rect 335628 633058 351826 633294
rect 352062 633058 352146 633294
rect 352382 633058 371826 633294
rect 372062 633058 372146 633294
rect 372382 633058 391826 633294
rect 392062 633058 392146 633294
rect 392382 633058 410328 633294
rect 410564 633058 505392 633294
rect 505628 633058 511826 633294
rect 512062 633058 512146 633294
rect 512382 633058 531826 633294
rect 532062 633058 532146 633294
rect 532382 633058 551826 633294
rect 552062 633058 552146 633294
rect 552382 633058 571826 633294
rect 572062 633058 572146 633294
rect 572382 633058 586302 633294
rect 586538 633058 586622 633294
rect 586858 633058 586890 633294
rect -2966 632896 586890 633058
rect -6806 630614 590730 630776
rect -6806 630378 -5814 630614
rect -5578 630378 -5494 630614
rect -5258 630378 9266 630614
rect 9502 630378 9586 630614
rect 9822 630378 169266 630614
rect 169502 630378 169586 630614
rect 169822 630378 189266 630614
rect 189502 630378 189586 630614
rect 189822 630378 209266 630614
rect 209502 630378 209586 630614
rect 209822 630378 229266 630614
rect 229502 630378 229586 630614
rect 229822 630378 349266 630614
rect 349502 630378 349586 630614
rect 349822 630378 369266 630614
rect 369502 630378 369586 630614
rect 369822 630378 389266 630614
rect 389502 630378 389586 630614
rect 389822 630378 509266 630614
rect 509502 630378 509586 630614
rect 509822 630378 529266 630614
rect 529502 630378 529586 630614
rect 529822 630378 549266 630614
rect 549502 630378 549586 630614
rect 549822 630378 569266 630614
rect 569502 630378 569586 630614
rect 569822 630378 589182 630614
rect 589418 630378 589502 630614
rect 589738 630378 590730 630614
rect -6806 630216 590730 630378
rect -4886 626954 588810 627116
rect -4886 626718 -3894 626954
rect -3658 626718 -3574 626954
rect -3338 626718 5546 626954
rect 5782 626718 5866 626954
rect 6102 626718 25546 626954
rect 25782 626718 25866 626954
rect 26102 626718 185546 626954
rect 185782 626718 185866 626954
rect 186102 626718 205546 626954
rect 205782 626718 205866 626954
rect 206102 626718 225546 626954
rect 225782 626718 225866 626954
rect 226102 626718 345546 626954
rect 345782 626718 345866 626954
rect 346102 626718 365546 626954
rect 365782 626718 365866 626954
rect 366102 626718 385546 626954
rect 385782 626718 385866 626954
rect 386102 626718 405546 626954
rect 405782 626718 405866 626954
rect 406102 626718 525546 626954
rect 525782 626718 525866 626954
rect 526102 626718 545546 626954
rect 545782 626718 545866 626954
rect 546102 626718 565546 626954
rect 565782 626718 565866 626954
rect 566102 626718 587262 626954
rect 587498 626718 587582 626954
rect 587818 626718 588810 626954
rect -4886 626556 588810 626718
rect -8726 624274 592650 624436
rect -8726 624038 -8694 624274
rect -8458 624038 -8374 624274
rect -8138 624038 22986 624274
rect 23222 624038 23306 624274
rect 23542 624038 182986 624274
rect 183222 624038 183306 624274
rect 183542 624038 202986 624274
rect 203222 624038 203306 624274
rect 203542 624038 222986 624274
rect 223222 624038 223306 624274
rect 223542 624038 342986 624274
rect 343222 624038 343306 624274
rect 343542 624038 362986 624274
rect 363222 624038 363306 624274
rect 363542 624038 382986 624274
rect 383222 624038 383306 624274
rect 383542 624038 402986 624274
rect 403222 624038 403306 624274
rect 403542 624038 522986 624274
rect 523222 624038 523306 624274
rect 523542 624038 542986 624274
rect 543222 624038 543306 624274
rect 543542 624038 562986 624274
rect 563222 624038 563306 624274
rect 563542 624038 592062 624274
rect 592298 624038 592382 624274
rect 592618 624038 592650 624274
rect -8726 623876 592650 624038
rect -2966 623294 586890 623456
rect -2966 623058 -1974 623294
rect -1738 623058 -1654 623294
rect -1418 623058 1826 623294
rect 2062 623058 2146 623294
rect 2382 623058 21826 623294
rect 22062 623058 22146 623294
rect 22382 623058 31008 623294
rect 31244 623058 165376 623294
rect 165612 623058 181826 623294
rect 182062 623058 182146 623294
rect 182382 623058 201826 623294
rect 202062 623058 202146 623294
rect 202382 623058 221826 623294
rect 222062 623058 222146 623294
rect 222382 623058 241008 623294
rect 241244 623058 334712 623294
rect 334948 623058 341826 623294
rect 342062 623058 342146 623294
rect 342382 623058 361826 623294
rect 362062 623058 362146 623294
rect 362382 623058 381826 623294
rect 382062 623058 382146 623294
rect 382382 623058 401826 623294
rect 402062 623058 402146 623294
rect 402382 623058 411008 623294
rect 411244 623058 504712 623294
rect 504948 623058 521826 623294
rect 522062 623058 522146 623294
rect 522382 623058 541826 623294
rect 542062 623058 542146 623294
rect 542382 623058 561826 623294
rect 562062 623058 562146 623294
rect 562382 623058 581826 623294
rect 582062 623058 582146 623294
rect 582382 623058 585342 623294
rect 585578 623058 585662 623294
rect 585898 623058 586890 623294
rect -2966 622896 586890 623058
rect -6806 620614 590730 620776
rect -6806 620378 -6774 620614
rect -6538 620378 -6454 620614
rect -6218 620378 19266 620614
rect 19502 620378 19586 620614
rect 19822 620378 179266 620614
rect 179502 620378 179586 620614
rect 179822 620378 199266 620614
rect 199502 620378 199586 620614
rect 199822 620378 219266 620614
rect 219502 620378 219586 620614
rect 219822 620378 339266 620614
rect 339502 620378 339586 620614
rect 339822 620378 359266 620614
rect 359502 620378 359586 620614
rect 359822 620378 379266 620614
rect 379502 620378 379586 620614
rect 379822 620378 399266 620614
rect 399502 620378 399586 620614
rect 399822 620378 519266 620614
rect 519502 620378 519586 620614
rect 519822 620378 539266 620614
rect 539502 620378 539586 620614
rect 539822 620378 559266 620614
rect 559502 620378 559586 620614
rect 559822 620378 579266 620614
rect 579502 620378 579586 620614
rect 579822 620378 590142 620614
rect 590378 620378 590462 620614
rect 590698 620378 590730 620614
rect -6806 620216 590730 620378
rect -4886 616954 588810 617116
rect -4886 616718 -4854 616954
rect -4618 616718 -4534 616954
rect -4298 616718 15546 616954
rect 15782 616718 15866 616954
rect 16102 616718 175546 616954
rect 175782 616718 175866 616954
rect 176102 616718 195546 616954
rect 195782 616718 195866 616954
rect 196102 616718 215546 616954
rect 215782 616718 215866 616954
rect 216102 616718 235546 616954
rect 235782 616718 235866 616954
rect 236102 616718 355546 616954
rect 355782 616718 355866 616954
rect 356102 616718 375546 616954
rect 375782 616718 375866 616954
rect 376102 616718 395546 616954
rect 395782 616718 395866 616954
rect 396102 616718 515546 616954
rect 515782 616718 515866 616954
rect 516102 616718 535546 616954
rect 535782 616718 535866 616954
rect 536102 616718 555546 616954
rect 555782 616718 555866 616954
rect 556102 616718 575546 616954
rect 575782 616718 575866 616954
rect 576102 616718 588222 616954
rect 588458 616718 588542 616954
rect 588778 616718 588810 616954
rect -4886 616556 588810 616718
rect -8726 614274 592650 614436
rect -8726 614038 -7734 614274
rect -7498 614038 -7414 614274
rect -7178 614038 12986 614274
rect 13222 614038 13306 614274
rect 13542 614038 172986 614274
rect 173222 614038 173306 614274
rect 173542 614038 192986 614274
rect 193222 614038 193306 614274
rect 193542 614038 212986 614274
rect 213222 614038 213306 614274
rect 213542 614038 232986 614274
rect 233222 614038 233306 614274
rect 233542 614038 352986 614274
rect 353222 614038 353306 614274
rect 353542 614038 372986 614274
rect 373222 614038 373306 614274
rect 373542 614038 392986 614274
rect 393222 614038 393306 614274
rect 393542 614038 512986 614274
rect 513222 614038 513306 614274
rect 513542 614038 532986 614274
rect 533222 614038 533306 614274
rect 533542 614038 552986 614274
rect 553222 614038 553306 614274
rect 553542 614038 572986 614274
rect 573222 614038 573306 614274
rect 573542 614038 591102 614274
rect 591338 614038 591422 614274
rect 591658 614038 592650 614274
rect -8726 613876 592650 614038
rect -2966 613294 586890 613456
rect -2966 613058 -2934 613294
rect -2698 613058 -2614 613294
rect -2378 613058 11826 613294
rect 12062 613058 12146 613294
rect 12382 613058 30328 613294
rect 30564 613058 166056 613294
rect 166292 613058 171826 613294
rect 172062 613058 172146 613294
rect 172382 613058 191826 613294
rect 192062 613058 192146 613294
rect 192382 613058 211826 613294
rect 212062 613058 212146 613294
rect 212382 613058 231826 613294
rect 232062 613058 232146 613294
rect 232382 613058 240328 613294
rect 240564 613058 335392 613294
rect 335628 613058 351826 613294
rect 352062 613058 352146 613294
rect 352382 613058 371826 613294
rect 372062 613058 372146 613294
rect 372382 613058 391826 613294
rect 392062 613058 392146 613294
rect 392382 613058 410328 613294
rect 410564 613058 505392 613294
rect 505628 613058 511826 613294
rect 512062 613058 512146 613294
rect 512382 613058 531826 613294
rect 532062 613058 532146 613294
rect 532382 613058 551826 613294
rect 552062 613058 552146 613294
rect 552382 613058 571826 613294
rect 572062 613058 572146 613294
rect 572382 613058 586302 613294
rect 586538 613058 586622 613294
rect 586858 613058 586890 613294
rect -2966 612896 586890 613058
rect -6806 610614 590730 610776
rect -6806 610378 -5814 610614
rect -5578 610378 -5494 610614
rect -5258 610378 9266 610614
rect 9502 610378 9586 610614
rect 9822 610378 169266 610614
rect 169502 610378 169586 610614
rect 169822 610378 189266 610614
rect 189502 610378 189586 610614
rect 189822 610378 209266 610614
rect 209502 610378 209586 610614
rect 209822 610378 229266 610614
rect 229502 610378 229586 610614
rect 229822 610378 349266 610614
rect 349502 610378 349586 610614
rect 349822 610378 369266 610614
rect 369502 610378 369586 610614
rect 369822 610378 389266 610614
rect 389502 610378 389586 610614
rect 389822 610378 509266 610614
rect 509502 610378 509586 610614
rect 509822 610378 529266 610614
rect 529502 610378 529586 610614
rect 529822 610378 549266 610614
rect 549502 610378 549586 610614
rect 549822 610378 569266 610614
rect 569502 610378 569586 610614
rect 569822 610378 589182 610614
rect 589418 610378 589502 610614
rect 589738 610378 590730 610614
rect -6806 610216 590730 610378
rect -4886 606954 588810 607116
rect -4886 606718 -3894 606954
rect -3658 606718 -3574 606954
rect -3338 606718 5546 606954
rect 5782 606718 5866 606954
rect 6102 606718 25546 606954
rect 25782 606718 25866 606954
rect 26102 606718 185546 606954
rect 185782 606718 185866 606954
rect 186102 606718 205546 606954
rect 205782 606718 205866 606954
rect 206102 606718 225546 606954
rect 225782 606718 225866 606954
rect 226102 606718 345546 606954
rect 345782 606718 345866 606954
rect 346102 606718 365546 606954
rect 365782 606718 365866 606954
rect 366102 606718 385546 606954
rect 385782 606718 385866 606954
rect 386102 606718 405546 606954
rect 405782 606718 405866 606954
rect 406102 606718 525546 606954
rect 525782 606718 525866 606954
rect 526102 606718 545546 606954
rect 545782 606718 545866 606954
rect 546102 606718 565546 606954
rect 565782 606718 565866 606954
rect 566102 606718 587262 606954
rect 587498 606718 587582 606954
rect 587818 606718 588810 606954
rect -4886 606556 588810 606718
rect -8726 604274 592650 604436
rect -8726 604038 -8694 604274
rect -8458 604038 -8374 604274
rect -8138 604038 22986 604274
rect 23222 604038 23306 604274
rect 23542 604038 182986 604274
rect 183222 604038 183306 604274
rect 183542 604038 202986 604274
rect 203222 604038 203306 604274
rect 203542 604038 222986 604274
rect 223222 604038 223306 604274
rect 223542 604038 342986 604274
rect 343222 604038 343306 604274
rect 343542 604038 362986 604274
rect 363222 604038 363306 604274
rect 363542 604038 382986 604274
rect 383222 604038 383306 604274
rect 383542 604038 402986 604274
rect 403222 604038 403306 604274
rect 403542 604038 522986 604274
rect 523222 604038 523306 604274
rect 523542 604038 542986 604274
rect 543222 604038 543306 604274
rect 543542 604038 562986 604274
rect 563222 604038 563306 604274
rect 563542 604038 592062 604274
rect 592298 604038 592382 604274
rect 592618 604038 592650 604274
rect -8726 603876 592650 604038
rect -2966 603294 586890 603456
rect -2966 603058 -1974 603294
rect -1738 603058 -1654 603294
rect -1418 603058 1826 603294
rect 2062 603058 2146 603294
rect 2382 603058 21826 603294
rect 22062 603058 22146 603294
rect 22382 603058 31008 603294
rect 31244 603058 165376 603294
rect 165612 603058 181826 603294
rect 182062 603058 182146 603294
rect 182382 603058 201826 603294
rect 202062 603058 202146 603294
rect 202382 603058 221826 603294
rect 222062 603058 222146 603294
rect 222382 603058 241008 603294
rect 241244 603058 334712 603294
rect 334948 603058 341826 603294
rect 342062 603058 342146 603294
rect 342382 603058 361826 603294
rect 362062 603058 362146 603294
rect 362382 603058 381826 603294
rect 382062 603058 382146 603294
rect 382382 603058 401826 603294
rect 402062 603058 402146 603294
rect 402382 603058 411008 603294
rect 411244 603058 504712 603294
rect 504948 603058 521826 603294
rect 522062 603058 522146 603294
rect 522382 603058 541826 603294
rect 542062 603058 542146 603294
rect 542382 603058 561826 603294
rect 562062 603058 562146 603294
rect 562382 603058 581826 603294
rect 582062 603058 582146 603294
rect 582382 603058 585342 603294
rect 585578 603058 585662 603294
rect 585898 603058 586890 603294
rect -2966 602896 586890 603058
rect -6806 600614 590730 600776
rect -6806 600378 -6774 600614
rect -6538 600378 -6454 600614
rect -6218 600378 19266 600614
rect 19502 600378 19586 600614
rect 19822 600378 179266 600614
rect 179502 600378 179586 600614
rect 179822 600378 199266 600614
rect 199502 600378 199586 600614
rect 199822 600378 219266 600614
rect 219502 600378 219586 600614
rect 219822 600378 339266 600614
rect 339502 600378 339586 600614
rect 339822 600378 359266 600614
rect 359502 600378 359586 600614
rect 359822 600378 379266 600614
rect 379502 600378 379586 600614
rect 379822 600378 399266 600614
rect 399502 600378 399586 600614
rect 399822 600378 519266 600614
rect 519502 600378 519586 600614
rect 519822 600378 539266 600614
rect 539502 600378 539586 600614
rect 539822 600378 559266 600614
rect 559502 600378 559586 600614
rect 559822 600378 579266 600614
rect 579502 600378 579586 600614
rect 579822 600378 590142 600614
rect 590378 600378 590462 600614
rect 590698 600378 590730 600614
rect -6806 600216 590730 600378
rect -4886 596954 588810 597116
rect -4886 596718 -4854 596954
rect -4618 596718 -4534 596954
rect -4298 596718 15546 596954
rect 15782 596718 15866 596954
rect 16102 596718 175546 596954
rect 175782 596718 175866 596954
rect 176102 596718 195546 596954
rect 195782 596718 195866 596954
rect 196102 596718 215546 596954
rect 215782 596718 215866 596954
rect 216102 596718 235546 596954
rect 235782 596718 235866 596954
rect 236102 596718 355546 596954
rect 355782 596718 355866 596954
rect 356102 596718 375546 596954
rect 375782 596718 375866 596954
rect 376102 596718 395546 596954
rect 395782 596718 395866 596954
rect 396102 596718 515546 596954
rect 515782 596718 515866 596954
rect 516102 596718 535546 596954
rect 535782 596718 535866 596954
rect 536102 596718 555546 596954
rect 555782 596718 555866 596954
rect 556102 596718 575546 596954
rect 575782 596718 575866 596954
rect 576102 596718 588222 596954
rect 588458 596718 588542 596954
rect 588778 596718 588810 596954
rect -4886 596556 588810 596718
rect -8726 594274 592650 594436
rect -8726 594038 -7734 594274
rect -7498 594038 -7414 594274
rect -7178 594038 12986 594274
rect 13222 594038 13306 594274
rect 13542 594038 172986 594274
rect 173222 594038 173306 594274
rect 173542 594038 192986 594274
rect 193222 594038 193306 594274
rect 193542 594038 212986 594274
rect 213222 594038 213306 594274
rect 213542 594038 232986 594274
rect 233222 594038 233306 594274
rect 233542 594038 352986 594274
rect 353222 594038 353306 594274
rect 353542 594038 372986 594274
rect 373222 594038 373306 594274
rect 373542 594038 392986 594274
rect 393222 594038 393306 594274
rect 393542 594038 512986 594274
rect 513222 594038 513306 594274
rect 513542 594038 532986 594274
rect 533222 594038 533306 594274
rect 533542 594038 552986 594274
rect 553222 594038 553306 594274
rect 553542 594038 572986 594274
rect 573222 594038 573306 594274
rect 573542 594038 591102 594274
rect 591338 594038 591422 594274
rect 591658 594038 592650 594274
rect -8726 593876 592650 594038
rect -2966 593294 586890 593456
rect -2966 593058 -2934 593294
rect -2698 593058 -2614 593294
rect -2378 593058 11826 593294
rect 12062 593058 12146 593294
rect 12382 593058 30328 593294
rect 30564 593058 166056 593294
rect 166292 593058 171826 593294
rect 172062 593058 172146 593294
rect 172382 593058 191826 593294
rect 192062 593058 192146 593294
rect 192382 593058 211826 593294
rect 212062 593058 212146 593294
rect 212382 593058 231826 593294
rect 232062 593058 232146 593294
rect 232382 593058 240328 593294
rect 240564 593058 335392 593294
rect 335628 593058 351826 593294
rect 352062 593058 352146 593294
rect 352382 593058 371826 593294
rect 372062 593058 372146 593294
rect 372382 593058 391826 593294
rect 392062 593058 392146 593294
rect 392382 593058 410328 593294
rect 410564 593058 505392 593294
rect 505628 593058 511826 593294
rect 512062 593058 512146 593294
rect 512382 593058 531826 593294
rect 532062 593058 532146 593294
rect 532382 593058 551826 593294
rect 552062 593058 552146 593294
rect 552382 593058 571826 593294
rect 572062 593058 572146 593294
rect 572382 593058 586302 593294
rect 586538 593058 586622 593294
rect 586858 593058 586890 593294
rect -2966 592896 586890 593058
rect -6806 590614 590730 590776
rect -6806 590378 -5814 590614
rect -5578 590378 -5494 590614
rect -5258 590378 9266 590614
rect 9502 590378 9586 590614
rect 9822 590378 169266 590614
rect 169502 590378 169586 590614
rect 169822 590378 189266 590614
rect 189502 590378 189586 590614
rect 189822 590378 209266 590614
rect 209502 590378 209586 590614
rect 209822 590378 229266 590614
rect 229502 590378 229586 590614
rect 229822 590378 349266 590614
rect 349502 590378 349586 590614
rect 349822 590378 369266 590614
rect 369502 590378 369586 590614
rect 369822 590378 389266 590614
rect 389502 590378 389586 590614
rect 389822 590378 509266 590614
rect 509502 590378 509586 590614
rect 509822 590378 529266 590614
rect 529502 590378 529586 590614
rect 529822 590378 549266 590614
rect 549502 590378 549586 590614
rect 549822 590378 569266 590614
rect 569502 590378 569586 590614
rect 569822 590378 589182 590614
rect 589418 590378 589502 590614
rect 589738 590378 590730 590614
rect -6806 590216 590730 590378
rect -4886 586954 588810 587116
rect -4886 586718 -3894 586954
rect -3658 586718 -3574 586954
rect -3338 586718 5546 586954
rect 5782 586718 5866 586954
rect 6102 586718 25546 586954
rect 25782 586718 25866 586954
rect 26102 586718 45546 586954
rect 45782 586718 45866 586954
rect 46102 586718 65546 586954
rect 65782 586718 65866 586954
rect 66102 586718 85546 586954
rect 85782 586718 85866 586954
rect 86102 586718 105546 586954
rect 105782 586718 105866 586954
rect 106102 586718 125546 586954
rect 125782 586718 125866 586954
rect 126102 586718 145546 586954
rect 145782 586718 145866 586954
rect 146102 586718 165546 586954
rect 165782 586718 165866 586954
rect 166102 586718 185546 586954
rect 185782 586718 185866 586954
rect 186102 586718 205546 586954
rect 205782 586718 205866 586954
rect 206102 586718 225546 586954
rect 225782 586718 225866 586954
rect 226102 586718 345546 586954
rect 345782 586718 345866 586954
rect 346102 586718 365546 586954
rect 365782 586718 365866 586954
rect 366102 586718 385546 586954
rect 385782 586718 385866 586954
rect 386102 586718 405546 586954
rect 405782 586718 405866 586954
rect 406102 586718 525546 586954
rect 525782 586718 525866 586954
rect 526102 586718 545546 586954
rect 545782 586718 545866 586954
rect 546102 586718 565546 586954
rect 565782 586718 565866 586954
rect 566102 586718 587262 586954
rect 587498 586718 587582 586954
rect 587818 586718 588810 586954
rect -4886 586556 588810 586718
rect -8726 584274 592650 584436
rect -8726 584038 -8694 584274
rect -8458 584038 -8374 584274
rect -8138 584038 22986 584274
rect 23222 584038 23306 584274
rect 23542 584038 42986 584274
rect 43222 584038 43306 584274
rect 43542 584038 62986 584274
rect 63222 584038 63306 584274
rect 63542 584038 82986 584274
rect 83222 584038 83306 584274
rect 83542 584038 102986 584274
rect 103222 584038 103306 584274
rect 103542 584038 122986 584274
rect 123222 584038 123306 584274
rect 123542 584038 142986 584274
rect 143222 584038 143306 584274
rect 143542 584038 162986 584274
rect 163222 584038 163306 584274
rect 163542 584038 182986 584274
rect 183222 584038 183306 584274
rect 183542 584038 202986 584274
rect 203222 584038 203306 584274
rect 203542 584038 222986 584274
rect 223222 584038 223306 584274
rect 223542 584038 342986 584274
rect 343222 584038 343306 584274
rect 343542 584038 362986 584274
rect 363222 584038 363306 584274
rect 363542 584038 382986 584274
rect 383222 584038 383306 584274
rect 383542 584038 402986 584274
rect 403222 584038 403306 584274
rect 403542 584038 522986 584274
rect 523222 584038 523306 584274
rect 523542 584038 542986 584274
rect 543222 584038 543306 584274
rect 543542 584038 562986 584274
rect 563222 584038 563306 584274
rect 563542 584038 592062 584274
rect 592298 584038 592382 584274
rect 592618 584038 592650 584274
rect -8726 583876 592650 584038
rect -2966 583294 586890 583456
rect -2966 583058 -1974 583294
rect -1738 583058 -1654 583294
rect -1418 583058 1826 583294
rect 2062 583058 2146 583294
rect 2382 583058 21826 583294
rect 22062 583058 22146 583294
rect 22382 583058 41826 583294
rect 42062 583058 42146 583294
rect 42382 583058 61826 583294
rect 62062 583058 62146 583294
rect 62382 583058 81826 583294
rect 82062 583058 82146 583294
rect 82382 583058 101826 583294
rect 102062 583058 102146 583294
rect 102382 583058 121826 583294
rect 122062 583058 122146 583294
rect 122382 583058 141826 583294
rect 142062 583058 142146 583294
rect 142382 583058 161826 583294
rect 162062 583058 162146 583294
rect 162382 583058 181826 583294
rect 182062 583058 182146 583294
rect 182382 583058 201826 583294
rect 202062 583058 202146 583294
rect 202382 583058 221826 583294
rect 222062 583058 222146 583294
rect 222382 583058 241008 583294
rect 241244 583058 334712 583294
rect 334948 583058 341826 583294
rect 342062 583058 342146 583294
rect 342382 583058 361826 583294
rect 362062 583058 362146 583294
rect 362382 583058 381826 583294
rect 382062 583058 382146 583294
rect 382382 583058 401826 583294
rect 402062 583058 402146 583294
rect 402382 583058 411008 583294
rect 411244 583058 504712 583294
rect 504948 583058 521826 583294
rect 522062 583058 522146 583294
rect 522382 583058 541826 583294
rect 542062 583058 542146 583294
rect 542382 583058 561826 583294
rect 562062 583058 562146 583294
rect 562382 583058 581826 583294
rect 582062 583058 582146 583294
rect 582382 583058 585342 583294
rect 585578 583058 585662 583294
rect 585898 583058 586890 583294
rect -2966 582896 586890 583058
rect -6806 580614 590730 580776
rect -6806 580378 -6774 580614
rect -6538 580378 -6454 580614
rect -6218 580378 19266 580614
rect 19502 580378 19586 580614
rect 19822 580378 39266 580614
rect 39502 580378 39586 580614
rect 39822 580378 59266 580614
rect 59502 580378 59586 580614
rect 59822 580378 79266 580614
rect 79502 580378 79586 580614
rect 79822 580378 99266 580614
rect 99502 580378 99586 580614
rect 99822 580378 119266 580614
rect 119502 580378 119586 580614
rect 119822 580378 139266 580614
rect 139502 580378 139586 580614
rect 139822 580378 159266 580614
rect 159502 580378 159586 580614
rect 159822 580378 179266 580614
rect 179502 580378 179586 580614
rect 179822 580378 199266 580614
rect 199502 580378 199586 580614
rect 199822 580378 219266 580614
rect 219502 580378 219586 580614
rect 219822 580378 339266 580614
rect 339502 580378 339586 580614
rect 339822 580378 359266 580614
rect 359502 580378 359586 580614
rect 359822 580378 379266 580614
rect 379502 580378 379586 580614
rect 379822 580378 399266 580614
rect 399502 580378 399586 580614
rect 399822 580378 519266 580614
rect 519502 580378 519586 580614
rect 519822 580378 539266 580614
rect 539502 580378 539586 580614
rect 539822 580378 559266 580614
rect 559502 580378 559586 580614
rect 559822 580378 579266 580614
rect 579502 580378 579586 580614
rect 579822 580378 590142 580614
rect 590378 580378 590462 580614
rect 590698 580378 590730 580614
rect -6806 580216 590730 580378
rect -4886 576954 588810 577116
rect -4886 576718 -4854 576954
rect -4618 576718 -4534 576954
rect -4298 576718 15546 576954
rect 15782 576718 15866 576954
rect 16102 576718 35546 576954
rect 35782 576718 35866 576954
rect 36102 576718 55546 576954
rect 55782 576718 55866 576954
rect 56102 576718 75546 576954
rect 75782 576718 75866 576954
rect 76102 576718 95546 576954
rect 95782 576718 95866 576954
rect 96102 576718 115546 576954
rect 115782 576718 115866 576954
rect 116102 576718 135546 576954
rect 135782 576718 135866 576954
rect 136102 576718 155546 576954
rect 155782 576718 155866 576954
rect 156102 576718 175546 576954
rect 175782 576718 175866 576954
rect 176102 576718 195546 576954
rect 195782 576718 195866 576954
rect 196102 576718 215546 576954
rect 215782 576718 215866 576954
rect 216102 576718 235546 576954
rect 235782 576718 235866 576954
rect 236102 576718 355546 576954
rect 355782 576718 355866 576954
rect 356102 576718 375546 576954
rect 375782 576718 375866 576954
rect 376102 576718 395546 576954
rect 395782 576718 395866 576954
rect 396102 576718 515546 576954
rect 515782 576718 515866 576954
rect 516102 576718 535546 576954
rect 535782 576718 535866 576954
rect 536102 576718 555546 576954
rect 555782 576718 555866 576954
rect 556102 576718 575546 576954
rect 575782 576718 575866 576954
rect 576102 576718 588222 576954
rect 588458 576718 588542 576954
rect 588778 576718 588810 576954
rect -4886 576556 588810 576718
rect -8726 574274 592650 574436
rect -8726 574038 -7734 574274
rect -7498 574038 -7414 574274
rect -7178 574038 12986 574274
rect 13222 574038 13306 574274
rect 13542 574038 32986 574274
rect 33222 574038 33306 574274
rect 33542 574038 52986 574274
rect 53222 574038 53306 574274
rect 53542 574038 72986 574274
rect 73222 574038 73306 574274
rect 73542 574038 92986 574274
rect 93222 574038 93306 574274
rect 93542 574038 112986 574274
rect 113222 574038 113306 574274
rect 113542 574038 132986 574274
rect 133222 574038 133306 574274
rect 133542 574038 152986 574274
rect 153222 574038 153306 574274
rect 153542 574038 172986 574274
rect 173222 574038 173306 574274
rect 173542 574038 192986 574274
rect 193222 574038 193306 574274
rect 193542 574038 212986 574274
rect 213222 574038 213306 574274
rect 213542 574038 232986 574274
rect 233222 574038 233306 574274
rect 233542 574038 252986 574274
rect 253222 574038 253306 574274
rect 253542 574038 272986 574274
rect 273222 574038 273306 574274
rect 273542 574038 292986 574274
rect 293222 574038 293306 574274
rect 293542 574038 312986 574274
rect 313222 574038 313306 574274
rect 313542 574038 332986 574274
rect 333222 574038 333306 574274
rect 333542 574038 352986 574274
rect 353222 574038 353306 574274
rect 353542 574038 372986 574274
rect 373222 574038 373306 574274
rect 373542 574038 392986 574274
rect 393222 574038 393306 574274
rect 393542 574038 412986 574274
rect 413222 574038 413306 574274
rect 413542 574038 432986 574274
rect 433222 574038 433306 574274
rect 433542 574038 452986 574274
rect 453222 574038 453306 574274
rect 453542 574038 472986 574274
rect 473222 574038 473306 574274
rect 473542 574038 492986 574274
rect 493222 574038 493306 574274
rect 493542 574038 512986 574274
rect 513222 574038 513306 574274
rect 513542 574038 532986 574274
rect 533222 574038 533306 574274
rect 533542 574038 552986 574274
rect 553222 574038 553306 574274
rect 553542 574038 572986 574274
rect 573222 574038 573306 574274
rect 573542 574038 591102 574274
rect 591338 574038 591422 574274
rect 591658 574038 592650 574274
rect -8726 573876 592650 574038
rect -2966 573294 586890 573456
rect -2966 573058 -2934 573294
rect -2698 573058 -2614 573294
rect -2378 573058 11826 573294
rect 12062 573058 12146 573294
rect 12382 573058 31826 573294
rect 32062 573058 32146 573294
rect 32382 573058 51826 573294
rect 52062 573058 52146 573294
rect 52382 573058 71826 573294
rect 72062 573058 72146 573294
rect 72382 573058 91826 573294
rect 92062 573058 92146 573294
rect 92382 573058 111826 573294
rect 112062 573058 112146 573294
rect 112382 573058 131826 573294
rect 132062 573058 132146 573294
rect 132382 573058 151826 573294
rect 152062 573058 152146 573294
rect 152382 573058 171826 573294
rect 172062 573058 172146 573294
rect 172382 573058 191826 573294
rect 192062 573058 192146 573294
rect 192382 573058 211826 573294
rect 212062 573058 212146 573294
rect 212382 573058 231826 573294
rect 232062 573058 232146 573294
rect 232382 573058 251826 573294
rect 252062 573058 252146 573294
rect 252382 573058 271826 573294
rect 272062 573058 272146 573294
rect 272382 573058 291826 573294
rect 292062 573058 292146 573294
rect 292382 573058 311826 573294
rect 312062 573058 312146 573294
rect 312382 573058 331826 573294
rect 332062 573058 332146 573294
rect 332382 573058 351826 573294
rect 352062 573058 352146 573294
rect 352382 573058 371826 573294
rect 372062 573058 372146 573294
rect 372382 573058 391826 573294
rect 392062 573058 392146 573294
rect 392382 573058 411826 573294
rect 412062 573058 412146 573294
rect 412382 573058 431826 573294
rect 432062 573058 432146 573294
rect 432382 573058 451826 573294
rect 452062 573058 452146 573294
rect 452382 573058 471826 573294
rect 472062 573058 472146 573294
rect 472382 573058 491826 573294
rect 492062 573058 492146 573294
rect 492382 573058 511826 573294
rect 512062 573058 512146 573294
rect 512382 573058 531826 573294
rect 532062 573058 532146 573294
rect 532382 573058 551826 573294
rect 552062 573058 552146 573294
rect 552382 573058 571826 573294
rect 572062 573058 572146 573294
rect 572382 573058 586302 573294
rect 586538 573058 586622 573294
rect 586858 573058 586890 573294
rect -2966 572896 586890 573058
rect -6806 570614 590730 570776
rect -6806 570378 -5814 570614
rect -5578 570378 -5494 570614
rect -5258 570378 9266 570614
rect 9502 570378 9586 570614
rect 9822 570378 29266 570614
rect 29502 570378 29586 570614
rect 29822 570378 49266 570614
rect 49502 570378 49586 570614
rect 49822 570378 69266 570614
rect 69502 570378 69586 570614
rect 69822 570378 89266 570614
rect 89502 570378 89586 570614
rect 89822 570378 109266 570614
rect 109502 570378 109586 570614
rect 109822 570378 129266 570614
rect 129502 570378 129586 570614
rect 129822 570378 149266 570614
rect 149502 570378 149586 570614
rect 149822 570378 169266 570614
rect 169502 570378 169586 570614
rect 169822 570378 189266 570614
rect 189502 570378 189586 570614
rect 189822 570378 209266 570614
rect 209502 570378 209586 570614
rect 209822 570378 229266 570614
rect 229502 570378 229586 570614
rect 229822 570378 249266 570614
rect 249502 570378 249586 570614
rect 249822 570378 269266 570614
rect 269502 570378 269586 570614
rect 269822 570378 289266 570614
rect 289502 570378 289586 570614
rect 289822 570378 309266 570614
rect 309502 570378 309586 570614
rect 309822 570378 329266 570614
rect 329502 570378 329586 570614
rect 329822 570378 349266 570614
rect 349502 570378 349586 570614
rect 349822 570378 369266 570614
rect 369502 570378 369586 570614
rect 369822 570378 389266 570614
rect 389502 570378 389586 570614
rect 389822 570378 409266 570614
rect 409502 570378 409586 570614
rect 409822 570378 429266 570614
rect 429502 570378 429586 570614
rect 429822 570378 449266 570614
rect 449502 570378 449586 570614
rect 449822 570378 469266 570614
rect 469502 570378 469586 570614
rect 469822 570378 489266 570614
rect 489502 570378 489586 570614
rect 489822 570378 509266 570614
rect 509502 570378 509586 570614
rect 509822 570378 529266 570614
rect 529502 570378 529586 570614
rect 529822 570378 549266 570614
rect 549502 570378 549586 570614
rect 549822 570378 569266 570614
rect 569502 570378 569586 570614
rect 569822 570378 589182 570614
rect 589418 570378 589502 570614
rect 589738 570378 590730 570614
rect -6806 570216 590730 570378
rect -4886 566954 588810 567116
rect -4886 566718 -3894 566954
rect -3658 566718 -3574 566954
rect -3338 566718 5546 566954
rect 5782 566718 5866 566954
rect 6102 566718 25546 566954
rect 25782 566718 25866 566954
rect 26102 566718 45546 566954
rect 45782 566718 45866 566954
rect 46102 566718 65546 566954
rect 65782 566718 65866 566954
rect 66102 566718 85546 566954
rect 85782 566718 85866 566954
rect 86102 566718 105546 566954
rect 105782 566718 105866 566954
rect 106102 566718 125546 566954
rect 125782 566718 125866 566954
rect 126102 566718 145546 566954
rect 145782 566718 145866 566954
rect 146102 566718 165546 566954
rect 165782 566718 165866 566954
rect 166102 566718 185546 566954
rect 185782 566718 185866 566954
rect 186102 566718 205546 566954
rect 205782 566718 205866 566954
rect 206102 566718 225546 566954
rect 225782 566718 225866 566954
rect 226102 566718 245546 566954
rect 245782 566718 245866 566954
rect 246102 566718 265546 566954
rect 265782 566718 265866 566954
rect 266102 566718 285546 566954
rect 285782 566718 285866 566954
rect 286102 566718 305546 566954
rect 305782 566718 305866 566954
rect 306102 566718 325546 566954
rect 325782 566718 325866 566954
rect 326102 566718 345546 566954
rect 345782 566718 345866 566954
rect 346102 566718 365546 566954
rect 365782 566718 365866 566954
rect 366102 566718 385546 566954
rect 385782 566718 385866 566954
rect 386102 566718 405546 566954
rect 405782 566718 405866 566954
rect 406102 566718 425546 566954
rect 425782 566718 425866 566954
rect 426102 566718 445546 566954
rect 445782 566718 445866 566954
rect 446102 566718 465546 566954
rect 465782 566718 465866 566954
rect 466102 566718 485546 566954
rect 485782 566718 485866 566954
rect 486102 566718 505546 566954
rect 505782 566718 505866 566954
rect 506102 566718 525546 566954
rect 525782 566718 525866 566954
rect 526102 566718 545546 566954
rect 545782 566718 545866 566954
rect 546102 566718 565546 566954
rect 565782 566718 565866 566954
rect 566102 566718 587262 566954
rect 587498 566718 587582 566954
rect 587818 566718 588810 566954
rect -4886 566556 588810 566718
rect -8726 564274 592650 564436
rect -8726 564038 -8694 564274
rect -8458 564038 -8374 564274
rect -8138 564038 22986 564274
rect 23222 564038 23306 564274
rect 23542 564038 42986 564274
rect 43222 564038 43306 564274
rect 43542 564038 62986 564274
rect 63222 564038 63306 564274
rect 63542 564038 82986 564274
rect 83222 564038 83306 564274
rect 83542 564038 102986 564274
rect 103222 564038 103306 564274
rect 103542 564038 122986 564274
rect 123222 564038 123306 564274
rect 123542 564038 142986 564274
rect 143222 564038 143306 564274
rect 143542 564038 162986 564274
rect 163222 564038 163306 564274
rect 163542 564038 182986 564274
rect 183222 564038 183306 564274
rect 183542 564038 202986 564274
rect 203222 564038 203306 564274
rect 203542 564038 222986 564274
rect 223222 564038 223306 564274
rect 223542 564038 242986 564274
rect 243222 564038 243306 564274
rect 243542 564038 262986 564274
rect 263222 564038 263306 564274
rect 263542 564038 282986 564274
rect 283222 564038 283306 564274
rect 283542 564038 302986 564274
rect 303222 564038 303306 564274
rect 303542 564038 322986 564274
rect 323222 564038 323306 564274
rect 323542 564038 342986 564274
rect 343222 564038 343306 564274
rect 343542 564038 362986 564274
rect 363222 564038 363306 564274
rect 363542 564038 382986 564274
rect 383222 564038 383306 564274
rect 383542 564038 402986 564274
rect 403222 564038 403306 564274
rect 403542 564038 422986 564274
rect 423222 564038 423306 564274
rect 423542 564038 442986 564274
rect 443222 564038 443306 564274
rect 443542 564038 462986 564274
rect 463222 564038 463306 564274
rect 463542 564038 482986 564274
rect 483222 564038 483306 564274
rect 483542 564038 502986 564274
rect 503222 564038 503306 564274
rect 503542 564038 522986 564274
rect 523222 564038 523306 564274
rect 523542 564038 542986 564274
rect 543222 564038 543306 564274
rect 543542 564038 562986 564274
rect 563222 564038 563306 564274
rect 563542 564038 592062 564274
rect 592298 564038 592382 564274
rect 592618 564038 592650 564274
rect -8726 563876 592650 564038
rect -2966 563294 586890 563456
rect -2966 563058 -1974 563294
rect -1738 563058 -1654 563294
rect -1418 563058 1826 563294
rect 2062 563058 2146 563294
rect 2382 563058 21826 563294
rect 22062 563058 22146 563294
rect 22382 563058 181826 563294
rect 182062 563058 182146 563294
rect 182382 563058 201826 563294
rect 202062 563058 202146 563294
rect 202382 563058 221826 563294
rect 222062 563058 222146 563294
rect 222382 563058 241826 563294
rect 242062 563058 242146 563294
rect 242382 563058 261826 563294
rect 262062 563058 262146 563294
rect 262382 563058 281826 563294
rect 282062 563058 282146 563294
rect 282382 563058 301826 563294
rect 302062 563058 302146 563294
rect 302382 563058 321826 563294
rect 322062 563058 322146 563294
rect 322382 563058 341826 563294
rect 342062 563058 342146 563294
rect 342382 563058 361826 563294
rect 362062 563058 362146 563294
rect 362382 563058 381826 563294
rect 382062 563058 382146 563294
rect 382382 563058 401826 563294
rect 402062 563058 402146 563294
rect 402382 563058 421826 563294
rect 422062 563058 422146 563294
rect 422382 563058 441826 563294
rect 442062 563058 442146 563294
rect 442382 563058 461826 563294
rect 462062 563058 462146 563294
rect 462382 563058 481826 563294
rect 482062 563058 482146 563294
rect 482382 563058 501826 563294
rect 502062 563058 502146 563294
rect 502382 563058 521826 563294
rect 522062 563058 522146 563294
rect 522382 563058 541826 563294
rect 542062 563058 542146 563294
rect 542382 563058 561826 563294
rect 562062 563058 562146 563294
rect 562382 563058 581826 563294
rect 582062 563058 582146 563294
rect 582382 563058 585342 563294
rect 585578 563058 585662 563294
rect 585898 563058 586890 563294
rect -2966 562896 586890 563058
rect -6806 560614 590730 560776
rect -6806 560378 -6774 560614
rect -6538 560378 -6454 560614
rect -6218 560378 19266 560614
rect 19502 560378 19586 560614
rect 19822 560378 179266 560614
rect 179502 560378 179586 560614
rect 179822 560378 199266 560614
rect 199502 560378 199586 560614
rect 199822 560378 219266 560614
rect 219502 560378 219586 560614
rect 219822 560378 239266 560614
rect 239502 560378 239586 560614
rect 239822 560378 259266 560614
rect 259502 560378 259586 560614
rect 259822 560378 279266 560614
rect 279502 560378 279586 560614
rect 279822 560378 299266 560614
rect 299502 560378 299586 560614
rect 299822 560378 319266 560614
rect 319502 560378 319586 560614
rect 319822 560378 339266 560614
rect 339502 560378 339586 560614
rect 339822 560378 359266 560614
rect 359502 560378 359586 560614
rect 359822 560378 379266 560614
rect 379502 560378 379586 560614
rect 379822 560378 399266 560614
rect 399502 560378 399586 560614
rect 399822 560378 419266 560614
rect 419502 560378 419586 560614
rect 419822 560378 439266 560614
rect 439502 560378 439586 560614
rect 439822 560378 459266 560614
rect 459502 560378 459586 560614
rect 459822 560378 479266 560614
rect 479502 560378 479586 560614
rect 479822 560378 499266 560614
rect 499502 560378 499586 560614
rect 499822 560378 519266 560614
rect 519502 560378 519586 560614
rect 519822 560378 539266 560614
rect 539502 560378 539586 560614
rect 539822 560378 559266 560614
rect 559502 560378 559586 560614
rect 559822 560378 579266 560614
rect 579502 560378 579586 560614
rect 579822 560378 590142 560614
rect 590378 560378 590462 560614
rect 590698 560378 590730 560614
rect -6806 560216 590730 560378
rect -4886 556954 588810 557116
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15546 556954
rect 15782 556718 15866 556954
rect 16102 556718 175546 556954
rect 175782 556718 175866 556954
rect 176102 556718 195546 556954
rect 195782 556718 195866 556954
rect 196102 556718 215546 556954
rect 215782 556718 215866 556954
rect 216102 556718 235546 556954
rect 235782 556718 235866 556954
rect 236102 556718 255546 556954
rect 255782 556718 255866 556954
rect 256102 556718 275546 556954
rect 275782 556718 275866 556954
rect 276102 556718 295546 556954
rect 295782 556718 295866 556954
rect 296102 556718 315546 556954
rect 315782 556718 315866 556954
rect 316102 556718 335546 556954
rect 335782 556718 335866 556954
rect 336102 556718 355546 556954
rect 355782 556718 355866 556954
rect 356102 556718 375546 556954
rect 375782 556718 375866 556954
rect 376102 556718 395546 556954
rect 395782 556718 395866 556954
rect 396102 556718 415546 556954
rect 415782 556718 415866 556954
rect 416102 556718 435546 556954
rect 435782 556718 435866 556954
rect 436102 556718 455546 556954
rect 455782 556718 455866 556954
rect 456102 556718 475546 556954
rect 475782 556718 475866 556954
rect 476102 556718 495546 556954
rect 495782 556718 495866 556954
rect 496102 556718 515546 556954
rect 515782 556718 515866 556954
rect 516102 556718 535546 556954
rect 535782 556718 535866 556954
rect 536102 556718 555546 556954
rect 555782 556718 555866 556954
rect 556102 556718 575546 556954
rect 575782 556718 575866 556954
rect 576102 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect -4886 556556 588810 556718
rect -8726 554274 592650 554436
rect -8726 554038 -7734 554274
rect -7498 554038 -7414 554274
rect -7178 554038 12986 554274
rect 13222 554038 13306 554274
rect 13542 554038 172986 554274
rect 173222 554038 173306 554274
rect 173542 554038 192986 554274
rect 193222 554038 193306 554274
rect 193542 554038 212986 554274
rect 213222 554038 213306 554274
rect 213542 554038 232986 554274
rect 233222 554038 233306 554274
rect 233542 554038 252986 554274
rect 253222 554038 253306 554274
rect 253542 554038 272986 554274
rect 273222 554038 273306 554274
rect 273542 554038 292986 554274
rect 293222 554038 293306 554274
rect 293542 554038 312986 554274
rect 313222 554038 313306 554274
rect 313542 554038 332986 554274
rect 333222 554038 333306 554274
rect 333542 554038 352986 554274
rect 353222 554038 353306 554274
rect 353542 554038 372986 554274
rect 373222 554038 373306 554274
rect 373542 554038 392986 554274
rect 393222 554038 393306 554274
rect 393542 554038 412986 554274
rect 413222 554038 413306 554274
rect 413542 554038 432986 554274
rect 433222 554038 433306 554274
rect 433542 554038 452986 554274
rect 453222 554038 453306 554274
rect 453542 554038 472986 554274
rect 473222 554038 473306 554274
rect 473542 554038 492986 554274
rect 493222 554038 493306 554274
rect 493542 554038 512986 554274
rect 513222 554038 513306 554274
rect 513542 554038 532986 554274
rect 533222 554038 533306 554274
rect 533542 554038 552986 554274
rect 553222 554038 553306 554274
rect 553542 554038 572986 554274
rect 573222 554038 573306 554274
rect 573542 554038 591102 554274
rect 591338 554038 591422 554274
rect 591658 554038 592650 554274
rect -8726 553876 592650 554038
rect -2966 553294 586890 553456
rect -2966 553058 -2934 553294
rect -2698 553058 -2614 553294
rect -2378 553058 11826 553294
rect 12062 553058 12146 553294
rect 12382 553058 30328 553294
rect 30564 553058 166056 553294
rect 166292 553058 171826 553294
rect 172062 553058 172146 553294
rect 172382 553058 191826 553294
rect 192062 553058 192146 553294
rect 192382 553058 211826 553294
rect 212062 553058 212146 553294
rect 212382 553058 231826 553294
rect 232062 553058 232146 553294
rect 232382 553058 251826 553294
rect 252062 553058 252146 553294
rect 252382 553058 271826 553294
rect 272062 553058 272146 553294
rect 272382 553058 291826 553294
rect 292062 553058 292146 553294
rect 292382 553058 311826 553294
rect 312062 553058 312146 553294
rect 312382 553058 331826 553294
rect 332062 553058 332146 553294
rect 332382 553058 351826 553294
rect 352062 553058 352146 553294
rect 352382 553058 371826 553294
rect 372062 553058 372146 553294
rect 372382 553058 391826 553294
rect 392062 553058 392146 553294
rect 392382 553058 411826 553294
rect 412062 553058 412146 553294
rect 412382 553058 431826 553294
rect 432062 553058 432146 553294
rect 432382 553058 451826 553294
rect 452062 553058 452146 553294
rect 452382 553058 471826 553294
rect 472062 553058 472146 553294
rect 472382 553058 491826 553294
rect 492062 553058 492146 553294
rect 492382 553058 511826 553294
rect 512062 553058 512146 553294
rect 512382 553058 531826 553294
rect 532062 553058 532146 553294
rect 532382 553058 551826 553294
rect 552062 553058 552146 553294
rect 552382 553058 571826 553294
rect 572062 553058 572146 553294
rect 572382 553058 586302 553294
rect 586538 553058 586622 553294
rect 586858 553058 586890 553294
rect -2966 552896 586890 553058
rect -6806 550614 590730 550776
rect -6806 550378 -5814 550614
rect -5578 550378 -5494 550614
rect -5258 550378 9266 550614
rect 9502 550378 9586 550614
rect 9822 550378 169266 550614
rect 169502 550378 169586 550614
rect 169822 550378 189266 550614
rect 189502 550378 189586 550614
rect 189822 550378 209266 550614
rect 209502 550378 209586 550614
rect 209822 550378 229266 550614
rect 229502 550378 229586 550614
rect 229822 550378 249266 550614
rect 249502 550378 249586 550614
rect 249822 550378 269266 550614
rect 269502 550378 269586 550614
rect 269822 550378 289266 550614
rect 289502 550378 289586 550614
rect 289822 550378 309266 550614
rect 309502 550378 309586 550614
rect 309822 550378 329266 550614
rect 329502 550378 329586 550614
rect 329822 550378 349266 550614
rect 349502 550378 349586 550614
rect 349822 550378 369266 550614
rect 369502 550378 369586 550614
rect 369822 550378 389266 550614
rect 389502 550378 389586 550614
rect 389822 550378 409266 550614
rect 409502 550378 409586 550614
rect 409822 550378 429266 550614
rect 429502 550378 429586 550614
rect 429822 550378 449266 550614
rect 449502 550378 449586 550614
rect 449822 550378 469266 550614
rect 469502 550378 469586 550614
rect 469822 550378 489266 550614
rect 489502 550378 489586 550614
rect 489822 550378 509266 550614
rect 509502 550378 509586 550614
rect 509822 550378 529266 550614
rect 529502 550378 529586 550614
rect 529822 550378 549266 550614
rect 549502 550378 549586 550614
rect 549822 550378 569266 550614
rect 569502 550378 569586 550614
rect 569822 550378 589182 550614
rect 589418 550378 589502 550614
rect 589738 550378 590730 550614
rect -6806 550216 590730 550378
rect -4886 546954 588810 547116
rect -4886 546718 -3894 546954
rect -3658 546718 -3574 546954
rect -3338 546718 5546 546954
rect 5782 546718 5866 546954
rect 6102 546718 25546 546954
rect 25782 546718 25866 546954
rect 26102 546718 185546 546954
rect 185782 546718 185866 546954
rect 186102 546718 205546 546954
rect 205782 546718 205866 546954
rect 206102 546718 225546 546954
rect 225782 546718 225866 546954
rect 226102 546718 245546 546954
rect 245782 546718 245866 546954
rect 246102 546718 265546 546954
rect 265782 546718 265866 546954
rect 266102 546718 285546 546954
rect 285782 546718 285866 546954
rect 286102 546718 305546 546954
rect 305782 546718 305866 546954
rect 306102 546718 325546 546954
rect 325782 546718 325866 546954
rect 326102 546718 345546 546954
rect 345782 546718 345866 546954
rect 346102 546718 365546 546954
rect 365782 546718 365866 546954
rect 366102 546718 385546 546954
rect 385782 546718 385866 546954
rect 386102 546718 405546 546954
rect 405782 546718 405866 546954
rect 406102 546718 425546 546954
rect 425782 546718 425866 546954
rect 426102 546718 445546 546954
rect 445782 546718 445866 546954
rect 446102 546718 465546 546954
rect 465782 546718 465866 546954
rect 466102 546718 485546 546954
rect 485782 546718 485866 546954
rect 486102 546718 505546 546954
rect 505782 546718 505866 546954
rect 506102 546718 525546 546954
rect 525782 546718 525866 546954
rect 526102 546718 545546 546954
rect 545782 546718 545866 546954
rect 546102 546718 565546 546954
rect 565782 546718 565866 546954
rect 566102 546718 587262 546954
rect 587498 546718 587582 546954
rect 587818 546718 588810 546954
rect -4886 546556 588810 546718
rect -8726 544274 592650 544436
rect -8726 544038 -8694 544274
rect -8458 544038 -8374 544274
rect -8138 544038 22986 544274
rect 23222 544038 23306 544274
rect 23542 544038 182986 544274
rect 183222 544038 183306 544274
rect 183542 544038 202986 544274
rect 203222 544038 203306 544274
rect 203542 544038 222986 544274
rect 223222 544038 223306 544274
rect 223542 544038 242986 544274
rect 243222 544038 243306 544274
rect 243542 544038 262986 544274
rect 263222 544038 263306 544274
rect 263542 544038 282986 544274
rect 283222 544038 283306 544274
rect 283542 544038 302986 544274
rect 303222 544038 303306 544274
rect 303542 544038 322986 544274
rect 323222 544038 323306 544274
rect 323542 544038 342986 544274
rect 343222 544038 343306 544274
rect 343542 544038 362986 544274
rect 363222 544038 363306 544274
rect 363542 544038 382986 544274
rect 383222 544038 383306 544274
rect 383542 544038 402986 544274
rect 403222 544038 403306 544274
rect 403542 544038 422986 544274
rect 423222 544038 423306 544274
rect 423542 544038 442986 544274
rect 443222 544038 443306 544274
rect 443542 544038 462986 544274
rect 463222 544038 463306 544274
rect 463542 544038 482986 544274
rect 483222 544038 483306 544274
rect 483542 544038 502986 544274
rect 503222 544038 503306 544274
rect 503542 544038 522986 544274
rect 523222 544038 523306 544274
rect 523542 544038 542986 544274
rect 543222 544038 543306 544274
rect 543542 544038 562986 544274
rect 563222 544038 563306 544274
rect 563542 544038 592062 544274
rect 592298 544038 592382 544274
rect 592618 544038 592650 544274
rect -8726 543876 592650 544038
rect -2966 543294 586890 543456
rect -2966 543058 -1974 543294
rect -1738 543058 -1654 543294
rect -1418 543058 1826 543294
rect 2062 543058 2146 543294
rect 2382 543058 21826 543294
rect 22062 543058 22146 543294
rect 22382 543058 31008 543294
rect 31244 543058 165376 543294
rect 165612 543058 181826 543294
rect 182062 543058 182146 543294
rect 182382 543058 201826 543294
rect 202062 543058 202146 543294
rect 202382 543058 221826 543294
rect 222062 543058 222146 543294
rect 222382 543058 241826 543294
rect 242062 543058 242146 543294
rect 242382 543058 261826 543294
rect 262062 543058 262146 543294
rect 262382 543058 281826 543294
rect 282062 543058 282146 543294
rect 282382 543058 301826 543294
rect 302062 543058 302146 543294
rect 302382 543058 321826 543294
rect 322062 543058 322146 543294
rect 322382 543058 341826 543294
rect 342062 543058 342146 543294
rect 342382 543058 361826 543294
rect 362062 543058 362146 543294
rect 362382 543058 381826 543294
rect 382062 543058 382146 543294
rect 382382 543058 401826 543294
rect 402062 543058 402146 543294
rect 402382 543058 421826 543294
rect 422062 543058 422146 543294
rect 422382 543058 441826 543294
rect 442062 543058 442146 543294
rect 442382 543058 461826 543294
rect 462062 543058 462146 543294
rect 462382 543058 481826 543294
rect 482062 543058 482146 543294
rect 482382 543058 501826 543294
rect 502062 543058 502146 543294
rect 502382 543058 521826 543294
rect 522062 543058 522146 543294
rect 522382 543058 541826 543294
rect 542062 543058 542146 543294
rect 542382 543058 561826 543294
rect 562062 543058 562146 543294
rect 562382 543058 581826 543294
rect 582062 543058 582146 543294
rect 582382 543058 585342 543294
rect 585578 543058 585662 543294
rect 585898 543058 586890 543294
rect -2966 542896 586890 543058
rect -6806 540614 590730 540776
rect -6806 540378 -6774 540614
rect -6538 540378 -6454 540614
rect -6218 540378 19266 540614
rect 19502 540378 19586 540614
rect 19822 540378 179266 540614
rect 179502 540378 179586 540614
rect 179822 540378 199266 540614
rect 199502 540378 199586 540614
rect 199822 540378 219266 540614
rect 219502 540378 219586 540614
rect 219822 540378 239266 540614
rect 239502 540378 239586 540614
rect 239822 540378 259266 540614
rect 259502 540378 259586 540614
rect 259822 540378 279266 540614
rect 279502 540378 279586 540614
rect 279822 540378 299266 540614
rect 299502 540378 299586 540614
rect 299822 540378 319266 540614
rect 319502 540378 319586 540614
rect 319822 540378 339266 540614
rect 339502 540378 339586 540614
rect 339822 540378 359266 540614
rect 359502 540378 359586 540614
rect 359822 540378 379266 540614
rect 379502 540378 379586 540614
rect 379822 540378 399266 540614
rect 399502 540378 399586 540614
rect 399822 540378 419266 540614
rect 419502 540378 419586 540614
rect 419822 540378 439266 540614
rect 439502 540378 439586 540614
rect 439822 540378 459266 540614
rect 459502 540378 459586 540614
rect 459822 540378 479266 540614
rect 479502 540378 479586 540614
rect 479822 540378 499266 540614
rect 499502 540378 499586 540614
rect 499822 540378 519266 540614
rect 519502 540378 519586 540614
rect 519822 540378 539266 540614
rect 539502 540378 539586 540614
rect 539822 540378 559266 540614
rect 559502 540378 559586 540614
rect 559822 540378 579266 540614
rect 579502 540378 579586 540614
rect 579822 540378 590142 540614
rect 590378 540378 590462 540614
rect 590698 540378 590730 540614
rect -6806 540216 590730 540378
rect -4886 536954 588810 537116
rect -4886 536718 -4854 536954
rect -4618 536718 -4534 536954
rect -4298 536718 15546 536954
rect 15782 536718 15866 536954
rect 16102 536718 175546 536954
rect 175782 536718 175866 536954
rect 176102 536718 195546 536954
rect 195782 536718 195866 536954
rect 196102 536718 355546 536954
rect 355782 536718 355866 536954
rect 356102 536718 375546 536954
rect 375782 536718 375866 536954
rect 376102 536718 395546 536954
rect 395782 536718 395866 536954
rect 396102 536718 555546 536954
rect 555782 536718 555866 536954
rect 556102 536718 575546 536954
rect 575782 536718 575866 536954
rect 576102 536718 588222 536954
rect 588458 536718 588542 536954
rect 588778 536718 588810 536954
rect -4886 536556 588810 536718
rect -8726 534274 592650 534436
rect -8726 534038 -7734 534274
rect -7498 534038 -7414 534274
rect -7178 534038 12986 534274
rect 13222 534038 13306 534274
rect 13542 534038 172986 534274
rect 173222 534038 173306 534274
rect 173542 534038 192986 534274
rect 193222 534038 193306 534274
rect 193542 534038 352986 534274
rect 353222 534038 353306 534274
rect 353542 534038 372986 534274
rect 373222 534038 373306 534274
rect 373542 534038 392986 534274
rect 393222 534038 393306 534274
rect 393542 534038 552986 534274
rect 553222 534038 553306 534274
rect 553542 534038 572986 534274
rect 573222 534038 573306 534274
rect 573542 534038 591102 534274
rect 591338 534038 591422 534274
rect 591658 534038 592650 534274
rect -8726 533876 592650 534038
rect -2966 533294 586890 533456
rect -2966 533058 -2934 533294
rect -2698 533058 -2614 533294
rect -2378 533058 11826 533294
rect 12062 533058 12146 533294
rect 12382 533058 30328 533294
rect 30564 533058 166056 533294
rect 166292 533058 171826 533294
rect 172062 533058 172146 533294
rect 172382 533058 191826 533294
rect 192062 533058 192146 533294
rect 192382 533058 200328 533294
rect 200564 533058 336056 533294
rect 336292 533058 351826 533294
rect 352062 533058 352146 533294
rect 352382 533058 371826 533294
rect 372062 533058 372146 533294
rect 372382 533058 391826 533294
rect 392062 533058 392146 533294
rect 392382 533058 410328 533294
rect 410564 533058 546056 533294
rect 546292 533058 551826 533294
rect 552062 533058 552146 533294
rect 552382 533058 571826 533294
rect 572062 533058 572146 533294
rect 572382 533058 586302 533294
rect 586538 533058 586622 533294
rect 586858 533058 586890 533294
rect -2966 532896 586890 533058
rect -6806 530614 590730 530776
rect -6806 530378 -5814 530614
rect -5578 530378 -5494 530614
rect -5258 530378 9266 530614
rect 9502 530378 9586 530614
rect 9822 530378 169266 530614
rect 169502 530378 169586 530614
rect 169822 530378 189266 530614
rect 189502 530378 189586 530614
rect 189822 530378 349266 530614
rect 349502 530378 349586 530614
rect 349822 530378 369266 530614
rect 369502 530378 369586 530614
rect 369822 530378 389266 530614
rect 389502 530378 389586 530614
rect 389822 530378 549266 530614
rect 549502 530378 549586 530614
rect 549822 530378 569266 530614
rect 569502 530378 569586 530614
rect 569822 530378 589182 530614
rect 589418 530378 589502 530614
rect 589738 530378 590730 530614
rect -6806 530216 590730 530378
rect -4886 526954 588810 527116
rect -4886 526718 -3894 526954
rect -3658 526718 -3574 526954
rect -3338 526718 5546 526954
rect 5782 526718 5866 526954
rect 6102 526718 25546 526954
rect 25782 526718 25866 526954
rect 26102 526718 185546 526954
rect 185782 526718 185866 526954
rect 186102 526718 345546 526954
rect 345782 526718 345866 526954
rect 346102 526718 365546 526954
rect 365782 526718 365866 526954
rect 366102 526718 385546 526954
rect 385782 526718 385866 526954
rect 386102 526718 405546 526954
rect 405782 526718 405866 526954
rect 406102 526718 565546 526954
rect 565782 526718 565866 526954
rect 566102 526718 587262 526954
rect 587498 526718 587582 526954
rect 587818 526718 588810 526954
rect -4886 526556 588810 526718
rect -8726 524274 592650 524436
rect -8726 524038 -8694 524274
rect -8458 524038 -8374 524274
rect -8138 524038 22986 524274
rect 23222 524038 23306 524274
rect 23542 524038 182986 524274
rect 183222 524038 183306 524274
rect 183542 524038 342986 524274
rect 343222 524038 343306 524274
rect 343542 524038 362986 524274
rect 363222 524038 363306 524274
rect 363542 524038 382986 524274
rect 383222 524038 383306 524274
rect 383542 524038 402986 524274
rect 403222 524038 403306 524274
rect 403542 524038 562986 524274
rect 563222 524038 563306 524274
rect 563542 524038 592062 524274
rect 592298 524038 592382 524274
rect 592618 524038 592650 524274
rect -8726 523876 592650 524038
rect -2966 523294 586890 523456
rect -2966 523058 -1974 523294
rect -1738 523058 -1654 523294
rect -1418 523058 1826 523294
rect 2062 523058 2146 523294
rect 2382 523058 21826 523294
rect 22062 523058 22146 523294
rect 22382 523058 31008 523294
rect 31244 523058 165376 523294
rect 165612 523058 181826 523294
rect 182062 523058 182146 523294
rect 182382 523058 201008 523294
rect 201244 523058 335376 523294
rect 335612 523058 341826 523294
rect 342062 523058 342146 523294
rect 342382 523058 361826 523294
rect 362062 523058 362146 523294
rect 362382 523058 381826 523294
rect 382062 523058 382146 523294
rect 382382 523058 401826 523294
rect 402062 523058 402146 523294
rect 402382 523058 411008 523294
rect 411244 523058 545376 523294
rect 545612 523058 561826 523294
rect 562062 523058 562146 523294
rect 562382 523058 581826 523294
rect 582062 523058 582146 523294
rect 582382 523058 585342 523294
rect 585578 523058 585662 523294
rect 585898 523058 586890 523294
rect -2966 522896 586890 523058
rect -6806 520614 590730 520776
rect -6806 520378 -6774 520614
rect -6538 520378 -6454 520614
rect -6218 520378 19266 520614
rect 19502 520378 19586 520614
rect 19822 520378 179266 520614
rect 179502 520378 179586 520614
rect 179822 520378 339266 520614
rect 339502 520378 339586 520614
rect 339822 520378 359266 520614
rect 359502 520378 359586 520614
rect 359822 520378 379266 520614
rect 379502 520378 379586 520614
rect 379822 520378 399266 520614
rect 399502 520378 399586 520614
rect 399822 520378 559266 520614
rect 559502 520378 559586 520614
rect 559822 520378 579266 520614
rect 579502 520378 579586 520614
rect 579822 520378 590142 520614
rect 590378 520378 590462 520614
rect 590698 520378 590730 520614
rect -6806 520216 590730 520378
rect -4886 516954 588810 517116
rect -4886 516718 -4854 516954
rect -4618 516718 -4534 516954
rect -4298 516718 15546 516954
rect 15782 516718 15866 516954
rect 16102 516718 175546 516954
rect 175782 516718 175866 516954
rect 176102 516718 195546 516954
rect 195782 516718 195866 516954
rect 196102 516718 355546 516954
rect 355782 516718 355866 516954
rect 356102 516718 375546 516954
rect 375782 516718 375866 516954
rect 376102 516718 395546 516954
rect 395782 516718 395866 516954
rect 396102 516718 555546 516954
rect 555782 516718 555866 516954
rect 556102 516718 575546 516954
rect 575782 516718 575866 516954
rect 576102 516718 588222 516954
rect 588458 516718 588542 516954
rect 588778 516718 588810 516954
rect -4886 516556 588810 516718
rect -8726 514274 592650 514436
rect -8726 514038 -7734 514274
rect -7498 514038 -7414 514274
rect -7178 514038 12986 514274
rect 13222 514038 13306 514274
rect 13542 514038 172986 514274
rect 173222 514038 173306 514274
rect 173542 514038 192986 514274
rect 193222 514038 193306 514274
rect 193542 514038 352986 514274
rect 353222 514038 353306 514274
rect 353542 514038 372986 514274
rect 373222 514038 373306 514274
rect 373542 514038 392986 514274
rect 393222 514038 393306 514274
rect 393542 514038 552986 514274
rect 553222 514038 553306 514274
rect 553542 514038 572986 514274
rect 573222 514038 573306 514274
rect 573542 514038 591102 514274
rect 591338 514038 591422 514274
rect 591658 514038 592650 514274
rect -8726 513876 592650 514038
rect -2966 513294 586890 513456
rect -2966 513058 -2934 513294
rect -2698 513058 -2614 513294
rect -2378 513058 11826 513294
rect 12062 513058 12146 513294
rect 12382 513058 30328 513294
rect 30564 513058 166056 513294
rect 166292 513058 171826 513294
rect 172062 513058 172146 513294
rect 172382 513058 191826 513294
rect 192062 513058 192146 513294
rect 192382 513058 200328 513294
rect 200564 513058 336056 513294
rect 336292 513058 351826 513294
rect 352062 513058 352146 513294
rect 352382 513058 371826 513294
rect 372062 513058 372146 513294
rect 372382 513058 391826 513294
rect 392062 513058 392146 513294
rect 392382 513058 410328 513294
rect 410564 513058 546056 513294
rect 546292 513058 551826 513294
rect 552062 513058 552146 513294
rect 552382 513058 571826 513294
rect 572062 513058 572146 513294
rect 572382 513058 586302 513294
rect 586538 513058 586622 513294
rect 586858 513058 586890 513294
rect -2966 512896 586890 513058
rect -6806 510614 590730 510776
rect -6806 510378 -5814 510614
rect -5578 510378 -5494 510614
rect -5258 510378 9266 510614
rect 9502 510378 9586 510614
rect 9822 510378 169266 510614
rect 169502 510378 169586 510614
rect 169822 510378 189266 510614
rect 189502 510378 189586 510614
rect 189822 510378 349266 510614
rect 349502 510378 349586 510614
rect 349822 510378 369266 510614
rect 369502 510378 369586 510614
rect 369822 510378 389266 510614
rect 389502 510378 389586 510614
rect 389822 510378 549266 510614
rect 549502 510378 549586 510614
rect 549822 510378 569266 510614
rect 569502 510378 569586 510614
rect 569822 510378 589182 510614
rect 589418 510378 589502 510614
rect 589738 510378 590730 510614
rect -6806 510216 590730 510378
rect -4886 506954 588810 507116
rect -4886 506718 -3894 506954
rect -3658 506718 -3574 506954
rect -3338 506718 5546 506954
rect 5782 506718 5866 506954
rect 6102 506718 25546 506954
rect 25782 506718 25866 506954
rect 26102 506718 185546 506954
rect 185782 506718 185866 506954
rect 186102 506718 345546 506954
rect 345782 506718 345866 506954
rect 346102 506718 365546 506954
rect 365782 506718 365866 506954
rect 366102 506718 385546 506954
rect 385782 506718 385866 506954
rect 386102 506718 405546 506954
rect 405782 506718 405866 506954
rect 406102 506718 565546 506954
rect 565782 506718 565866 506954
rect 566102 506718 587262 506954
rect 587498 506718 587582 506954
rect 587818 506718 588810 506954
rect -4886 506556 588810 506718
rect -8726 504274 592650 504436
rect -8726 504038 -8694 504274
rect -8458 504038 -8374 504274
rect -8138 504038 22986 504274
rect 23222 504038 23306 504274
rect 23542 504038 182986 504274
rect 183222 504038 183306 504274
rect 183542 504038 342986 504274
rect 343222 504038 343306 504274
rect 343542 504038 362986 504274
rect 363222 504038 363306 504274
rect 363542 504038 382986 504274
rect 383222 504038 383306 504274
rect 383542 504038 402986 504274
rect 403222 504038 403306 504274
rect 403542 504038 562986 504274
rect 563222 504038 563306 504274
rect 563542 504038 592062 504274
rect 592298 504038 592382 504274
rect 592618 504038 592650 504274
rect -8726 503876 592650 504038
rect -2966 503294 586890 503456
rect -2966 503058 -1974 503294
rect -1738 503058 -1654 503294
rect -1418 503058 1826 503294
rect 2062 503058 2146 503294
rect 2382 503058 21826 503294
rect 22062 503058 22146 503294
rect 22382 503058 31008 503294
rect 31244 503058 165376 503294
rect 165612 503058 181826 503294
rect 182062 503058 182146 503294
rect 182382 503058 201008 503294
rect 201244 503058 335376 503294
rect 335612 503058 341826 503294
rect 342062 503058 342146 503294
rect 342382 503058 361826 503294
rect 362062 503058 362146 503294
rect 362382 503058 381826 503294
rect 382062 503058 382146 503294
rect 382382 503058 401826 503294
rect 402062 503058 402146 503294
rect 402382 503058 411008 503294
rect 411244 503058 545376 503294
rect 545612 503058 561826 503294
rect 562062 503058 562146 503294
rect 562382 503058 581826 503294
rect 582062 503058 582146 503294
rect 582382 503058 585342 503294
rect 585578 503058 585662 503294
rect 585898 503058 586890 503294
rect -2966 502896 586890 503058
rect -6806 500614 590730 500776
rect -6806 500378 -6774 500614
rect -6538 500378 -6454 500614
rect -6218 500378 19266 500614
rect 19502 500378 19586 500614
rect 19822 500378 179266 500614
rect 179502 500378 179586 500614
rect 179822 500378 339266 500614
rect 339502 500378 339586 500614
rect 339822 500378 359266 500614
rect 359502 500378 359586 500614
rect 359822 500378 379266 500614
rect 379502 500378 379586 500614
rect 379822 500378 399266 500614
rect 399502 500378 399586 500614
rect 399822 500378 559266 500614
rect 559502 500378 559586 500614
rect 559822 500378 579266 500614
rect 579502 500378 579586 500614
rect 579822 500378 590142 500614
rect 590378 500378 590462 500614
rect 590698 500378 590730 500614
rect -6806 500216 590730 500378
rect -4886 496954 588810 497116
rect -4886 496718 -4854 496954
rect -4618 496718 -4534 496954
rect -4298 496718 15546 496954
rect 15782 496718 15866 496954
rect 16102 496718 175546 496954
rect 175782 496718 175866 496954
rect 176102 496718 195546 496954
rect 195782 496718 195866 496954
rect 196102 496718 355546 496954
rect 355782 496718 355866 496954
rect 356102 496718 375546 496954
rect 375782 496718 375866 496954
rect 376102 496718 395546 496954
rect 395782 496718 395866 496954
rect 396102 496718 555546 496954
rect 555782 496718 555866 496954
rect 556102 496718 575546 496954
rect 575782 496718 575866 496954
rect 576102 496718 588222 496954
rect 588458 496718 588542 496954
rect 588778 496718 588810 496954
rect -4886 496556 588810 496718
rect -8726 494274 592650 494436
rect -8726 494038 -7734 494274
rect -7498 494038 -7414 494274
rect -7178 494038 12986 494274
rect 13222 494038 13306 494274
rect 13542 494038 172986 494274
rect 173222 494038 173306 494274
rect 173542 494038 192986 494274
rect 193222 494038 193306 494274
rect 193542 494038 352986 494274
rect 353222 494038 353306 494274
rect 353542 494038 372986 494274
rect 373222 494038 373306 494274
rect 373542 494038 392986 494274
rect 393222 494038 393306 494274
rect 393542 494038 552986 494274
rect 553222 494038 553306 494274
rect 553542 494038 572986 494274
rect 573222 494038 573306 494274
rect 573542 494038 591102 494274
rect 591338 494038 591422 494274
rect 591658 494038 592650 494274
rect -8726 493876 592650 494038
rect -2966 493294 586890 493456
rect -2966 493058 -2934 493294
rect -2698 493058 -2614 493294
rect -2378 493058 11826 493294
rect 12062 493058 12146 493294
rect 12382 493058 30328 493294
rect 30564 493058 166056 493294
rect 166292 493058 171826 493294
rect 172062 493058 172146 493294
rect 172382 493058 191826 493294
rect 192062 493058 192146 493294
rect 192382 493058 200328 493294
rect 200564 493058 336056 493294
rect 336292 493058 351826 493294
rect 352062 493058 352146 493294
rect 352382 493058 371826 493294
rect 372062 493058 372146 493294
rect 372382 493058 391826 493294
rect 392062 493058 392146 493294
rect 392382 493058 410328 493294
rect 410564 493058 546056 493294
rect 546292 493058 551826 493294
rect 552062 493058 552146 493294
rect 552382 493058 571826 493294
rect 572062 493058 572146 493294
rect 572382 493058 586302 493294
rect 586538 493058 586622 493294
rect 586858 493058 586890 493294
rect -2966 492896 586890 493058
rect -6806 490614 590730 490776
rect -6806 490378 -5814 490614
rect -5578 490378 -5494 490614
rect -5258 490378 9266 490614
rect 9502 490378 9586 490614
rect 9822 490378 169266 490614
rect 169502 490378 169586 490614
rect 169822 490378 189266 490614
rect 189502 490378 189586 490614
rect 189822 490378 349266 490614
rect 349502 490378 349586 490614
rect 349822 490378 369266 490614
rect 369502 490378 369586 490614
rect 369822 490378 389266 490614
rect 389502 490378 389586 490614
rect 389822 490378 549266 490614
rect 549502 490378 549586 490614
rect 549822 490378 569266 490614
rect 569502 490378 569586 490614
rect 569822 490378 589182 490614
rect 589418 490378 589502 490614
rect 589738 490378 590730 490614
rect -6806 490216 590730 490378
rect -4886 486954 588810 487116
rect -4886 486718 -3894 486954
rect -3658 486718 -3574 486954
rect -3338 486718 5546 486954
rect 5782 486718 5866 486954
rect 6102 486718 25546 486954
rect 25782 486718 25866 486954
rect 26102 486718 185546 486954
rect 185782 486718 185866 486954
rect 186102 486718 345546 486954
rect 345782 486718 345866 486954
rect 346102 486718 365546 486954
rect 365782 486718 365866 486954
rect 366102 486718 385546 486954
rect 385782 486718 385866 486954
rect 386102 486718 405546 486954
rect 405782 486718 405866 486954
rect 406102 486718 565546 486954
rect 565782 486718 565866 486954
rect 566102 486718 587262 486954
rect 587498 486718 587582 486954
rect 587818 486718 588810 486954
rect -4886 486556 588810 486718
rect -8726 484274 592650 484436
rect -8726 484038 -8694 484274
rect -8458 484038 -8374 484274
rect -8138 484038 22986 484274
rect 23222 484038 23306 484274
rect 23542 484038 182986 484274
rect 183222 484038 183306 484274
rect 183542 484038 342986 484274
rect 343222 484038 343306 484274
rect 343542 484038 362986 484274
rect 363222 484038 363306 484274
rect 363542 484038 382986 484274
rect 383222 484038 383306 484274
rect 383542 484038 402986 484274
rect 403222 484038 403306 484274
rect 403542 484038 562986 484274
rect 563222 484038 563306 484274
rect 563542 484038 592062 484274
rect 592298 484038 592382 484274
rect 592618 484038 592650 484274
rect -8726 483876 592650 484038
rect -2966 483294 586890 483456
rect -2966 483058 -1974 483294
rect -1738 483058 -1654 483294
rect -1418 483058 1826 483294
rect 2062 483058 2146 483294
rect 2382 483058 21826 483294
rect 22062 483058 22146 483294
rect 22382 483058 31008 483294
rect 31244 483058 165376 483294
rect 165612 483058 181826 483294
rect 182062 483058 182146 483294
rect 182382 483058 201008 483294
rect 201244 483058 335376 483294
rect 335612 483058 341826 483294
rect 342062 483058 342146 483294
rect 342382 483058 361826 483294
rect 362062 483058 362146 483294
rect 362382 483058 381826 483294
rect 382062 483058 382146 483294
rect 382382 483058 401826 483294
rect 402062 483058 402146 483294
rect 402382 483058 411008 483294
rect 411244 483058 545376 483294
rect 545612 483058 561826 483294
rect 562062 483058 562146 483294
rect 562382 483058 581826 483294
rect 582062 483058 582146 483294
rect 582382 483058 585342 483294
rect 585578 483058 585662 483294
rect 585898 483058 586890 483294
rect -2966 482896 586890 483058
rect -6806 480614 590730 480776
rect -6806 480378 -6774 480614
rect -6538 480378 -6454 480614
rect -6218 480378 19266 480614
rect 19502 480378 19586 480614
rect 19822 480378 179266 480614
rect 179502 480378 179586 480614
rect 179822 480378 339266 480614
rect 339502 480378 339586 480614
rect 339822 480378 359266 480614
rect 359502 480378 359586 480614
rect 359822 480378 379266 480614
rect 379502 480378 379586 480614
rect 379822 480378 399266 480614
rect 399502 480378 399586 480614
rect 399822 480378 559266 480614
rect 559502 480378 559586 480614
rect 559822 480378 579266 480614
rect 579502 480378 579586 480614
rect 579822 480378 590142 480614
rect 590378 480378 590462 480614
rect 590698 480378 590730 480614
rect -6806 480216 590730 480378
rect -4886 476954 588810 477116
rect -4886 476718 -4854 476954
rect -4618 476718 -4534 476954
rect -4298 476718 15546 476954
rect 15782 476718 15866 476954
rect 16102 476718 175546 476954
rect 175782 476718 175866 476954
rect 176102 476718 195546 476954
rect 195782 476718 195866 476954
rect 196102 476718 355546 476954
rect 355782 476718 355866 476954
rect 356102 476718 375546 476954
rect 375782 476718 375866 476954
rect 376102 476718 395546 476954
rect 395782 476718 395866 476954
rect 396102 476718 555546 476954
rect 555782 476718 555866 476954
rect 556102 476718 575546 476954
rect 575782 476718 575866 476954
rect 576102 476718 588222 476954
rect 588458 476718 588542 476954
rect 588778 476718 588810 476954
rect -4886 476556 588810 476718
rect -8726 474274 592650 474436
rect -8726 474038 -7734 474274
rect -7498 474038 -7414 474274
rect -7178 474038 12986 474274
rect 13222 474038 13306 474274
rect 13542 474038 32986 474274
rect 33222 474038 33306 474274
rect 33542 474038 52986 474274
rect 53222 474038 53306 474274
rect 53542 474038 72986 474274
rect 73222 474038 73306 474274
rect 73542 474038 92986 474274
rect 93222 474038 93306 474274
rect 93542 474038 112986 474274
rect 113222 474038 113306 474274
rect 113542 474038 132986 474274
rect 133222 474038 133306 474274
rect 133542 474038 152986 474274
rect 153222 474038 153306 474274
rect 153542 474038 172986 474274
rect 173222 474038 173306 474274
rect 173542 474038 192986 474274
rect 193222 474038 193306 474274
rect 193542 474038 352986 474274
rect 353222 474038 353306 474274
rect 353542 474038 372986 474274
rect 373222 474038 373306 474274
rect 373542 474038 392986 474274
rect 393222 474038 393306 474274
rect 393542 474038 552986 474274
rect 553222 474038 553306 474274
rect 553542 474038 572986 474274
rect 573222 474038 573306 474274
rect 573542 474038 591102 474274
rect 591338 474038 591422 474274
rect 591658 474038 592650 474274
rect -8726 473876 592650 474038
rect -2966 473294 586890 473456
rect -2966 473058 -2934 473294
rect -2698 473058 -2614 473294
rect -2378 473058 11826 473294
rect 12062 473058 12146 473294
rect 12382 473058 31826 473294
rect 32062 473058 32146 473294
rect 32382 473058 51826 473294
rect 52062 473058 52146 473294
rect 52382 473058 71826 473294
rect 72062 473058 72146 473294
rect 72382 473058 91826 473294
rect 92062 473058 92146 473294
rect 92382 473058 111826 473294
rect 112062 473058 112146 473294
rect 112382 473058 131826 473294
rect 132062 473058 132146 473294
rect 132382 473058 151826 473294
rect 152062 473058 152146 473294
rect 152382 473058 171826 473294
rect 172062 473058 172146 473294
rect 172382 473058 191826 473294
rect 192062 473058 192146 473294
rect 192382 473058 200328 473294
rect 200564 473058 336056 473294
rect 336292 473058 351826 473294
rect 352062 473058 352146 473294
rect 352382 473058 371826 473294
rect 372062 473058 372146 473294
rect 372382 473058 391826 473294
rect 392062 473058 392146 473294
rect 392382 473058 410328 473294
rect 410564 473058 546056 473294
rect 546292 473058 551826 473294
rect 552062 473058 552146 473294
rect 552382 473058 571826 473294
rect 572062 473058 572146 473294
rect 572382 473058 586302 473294
rect 586538 473058 586622 473294
rect 586858 473058 586890 473294
rect -2966 472896 586890 473058
rect -6806 470614 590730 470776
rect -6806 470378 -5814 470614
rect -5578 470378 -5494 470614
rect -5258 470378 9266 470614
rect 9502 470378 9586 470614
rect 9822 470378 29266 470614
rect 29502 470378 29586 470614
rect 29822 470378 49266 470614
rect 49502 470378 49586 470614
rect 49822 470378 69266 470614
rect 69502 470378 69586 470614
rect 69822 470378 89266 470614
rect 89502 470378 89586 470614
rect 89822 470378 109266 470614
rect 109502 470378 109586 470614
rect 109822 470378 129266 470614
rect 129502 470378 129586 470614
rect 129822 470378 149266 470614
rect 149502 470378 149586 470614
rect 149822 470378 169266 470614
rect 169502 470378 169586 470614
rect 169822 470378 189266 470614
rect 189502 470378 189586 470614
rect 189822 470378 349266 470614
rect 349502 470378 349586 470614
rect 349822 470378 369266 470614
rect 369502 470378 369586 470614
rect 369822 470378 389266 470614
rect 389502 470378 389586 470614
rect 389822 470378 549266 470614
rect 549502 470378 549586 470614
rect 549822 470378 569266 470614
rect 569502 470378 569586 470614
rect 569822 470378 589182 470614
rect 589418 470378 589502 470614
rect 589738 470378 590730 470614
rect -6806 470216 590730 470378
rect -4886 466954 588810 467116
rect -4886 466718 -3894 466954
rect -3658 466718 -3574 466954
rect -3338 466718 5546 466954
rect 5782 466718 5866 466954
rect 6102 466718 25546 466954
rect 25782 466718 25866 466954
rect 26102 466718 45546 466954
rect 45782 466718 45866 466954
rect 46102 466718 65546 466954
rect 65782 466718 65866 466954
rect 66102 466718 85546 466954
rect 85782 466718 85866 466954
rect 86102 466718 105546 466954
rect 105782 466718 105866 466954
rect 106102 466718 125546 466954
rect 125782 466718 125866 466954
rect 126102 466718 145546 466954
rect 145782 466718 145866 466954
rect 146102 466718 165546 466954
rect 165782 466718 165866 466954
rect 166102 466718 185546 466954
rect 185782 466718 185866 466954
rect 186102 466718 345546 466954
rect 345782 466718 345866 466954
rect 346102 466718 365546 466954
rect 365782 466718 365866 466954
rect 366102 466718 385546 466954
rect 385782 466718 385866 466954
rect 386102 466718 405546 466954
rect 405782 466718 405866 466954
rect 406102 466718 565546 466954
rect 565782 466718 565866 466954
rect 566102 466718 587262 466954
rect 587498 466718 587582 466954
rect 587818 466718 588810 466954
rect -4886 466556 588810 466718
rect -8726 464274 592650 464436
rect -8726 464038 -8694 464274
rect -8458 464038 -8374 464274
rect -8138 464038 22986 464274
rect 23222 464038 23306 464274
rect 23542 464038 42986 464274
rect 43222 464038 43306 464274
rect 43542 464038 62986 464274
rect 63222 464038 63306 464274
rect 63542 464038 82986 464274
rect 83222 464038 83306 464274
rect 83542 464038 102986 464274
rect 103222 464038 103306 464274
rect 103542 464038 122986 464274
rect 123222 464038 123306 464274
rect 123542 464038 142986 464274
rect 143222 464038 143306 464274
rect 143542 464038 162986 464274
rect 163222 464038 163306 464274
rect 163542 464038 182986 464274
rect 183222 464038 183306 464274
rect 183542 464038 342986 464274
rect 343222 464038 343306 464274
rect 343542 464038 362986 464274
rect 363222 464038 363306 464274
rect 363542 464038 382986 464274
rect 383222 464038 383306 464274
rect 383542 464038 402986 464274
rect 403222 464038 403306 464274
rect 403542 464038 562986 464274
rect 563222 464038 563306 464274
rect 563542 464038 592062 464274
rect 592298 464038 592382 464274
rect 592618 464038 592650 464274
rect -8726 463876 592650 464038
rect -2966 463294 586890 463456
rect -2966 463058 -1974 463294
rect -1738 463058 -1654 463294
rect -1418 463058 1826 463294
rect 2062 463058 2146 463294
rect 2382 463058 21826 463294
rect 22062 463058 22146 463294
rect 22382 463058 41826 463294
rect 42062 463058 42146 463294
rect 42382 463058 61826 463294
rect 62062 463058 62146 463294
rect 62382 463058 81826 463294
rect 82062 463058 82146 463294
rect 82382 463058 101826 463294
rect 102062 463058 102146 463294
rect 102382 463058 121826 463294
rect 122062 463058 122146 463294
rect 122382 463058 141826 463294
rect 142062 463058 142146 463294
rect 142382 463058 161826 463294
rect 162062 463058 162146 463294
rect 162382 463058 181826 463294
rect 182062 463058 182146 463294
rect 182382 463058 201008 463294
rect 201244 463058 335376 463294
rect 335612 463058 341826 463294
rect 342062 463058 342146 463294
rect 342382 463058 361826 463294
rect 362062 463058 362146 463294
rect 362382 463058 381826 463294
rect 382062 463058 382146 463294
rect 382382 463058 401826 463294
rect 402062 463058 402146 463294
rect 402382 463058 411008 463294
rect 411244 463058 545376 463294
rect 545612 463058 561826 463294
rect 562062 463058 562146 463294
rect 562382 463058 581826 463294
rect 582062 463058 582146 463294
rect 582382 463058 585342 463294
rect 585578 463058 585662 463294
rect 585898 463058 586890 463294
rect -2966 462896 586890 463058
rect -6806 460614 590730 460776
rect -6806 460378 -6774 460614
rect -6538 460378 -6454 460614
rect -6218 460378 19266 460614
rect 19502 460378 19586 460614
rect 19822 460378 39266 460614
rect 39502 460378 39586 460614
rect 39822 460378 59266 460614
rect 59502 460378 59586 460614
rect 59822 460378 79266 460614
rect 79502 460378 79586 460614
rect 79822 460378 99266 460614
rect 99502 460378 99586 460614
rect 99822 460378 119266 460614
rect 119502 460378 119586 460614
rect 119822 460378 139266 460614
rect 139502 460378 139586 460614
rect 139822 460378 159266 460614
rect 159502 460378 159586 460614
rect 159822 460378 179266 460614
rect 179502 460378 179586 460614
rect 179822 460378 339266 460614
rect 339502 460378 339586 460614
rect 339822 460378 359266 460614
rect 359502 460378 359586 460614
rect 359822 460378 379266 460614
rect 379502 460378 379586 460614
rect 379822 460378 399266 460614
rect 399502 460378 399586 460614
rect 399822 460378 559266 460614
rect 559502 460378 559586 460614
rect 559822 460378 579266 460614
rect 579502 460378 579586 460614
rect 579822 460378 590142 460614
rect 590378 460378 590462 460614
rect 590698 460378 590730 460614
rect -6806 460216 590730 460378
rect -4886 456954 588810 457116
rect -4886 456718 -4854 456954
rect -4618 456718 -4534 456954
rect -4298 456718 15546 456954
rect 15782 456718 15866 456954
rect 16102 456718 35546 456954
rect 35782 456718 35866 456954
rect 36102 456718 55546 456954
rect 55782 456718 55866 456954
rect 56102 456718 75546 456954
rect 75782 456718 75866 456954
rect 76102 456718 95546 456954
rect 95782 456718 95866 456954
rect 96102 456718 115546 456954
rect 115782 456718 115866 456954
rect 116102 456718 135546 456954
rect 135782 456718 135866 456954
rect 136102 456718 155546 456954
rect 155782 456718 155866 456954
rect 156102 456718 175546 456954
rect 175782 456718 175866 456954
rect 176102 456718 195546 456954
rect 195782 456718 195866 456954
rect 196102 456718 355546 456954
rect 355782 456718 355866 456954
rect 356102 456718 375546 456954
rect 375782 456718 375866 456954
rect 376102 456718 395546 456954
rect 395782 456718 395866 456954
rect 396102 456718 555546 456954
rect 555782 456718 555866 456954
rect 556102 456718 575546 456954
rect 575782 456718 575866 456954
rect 576102 456718 588222 456954
rect 588458 456718 588542 456954
rect 588778 456718 588810 456954
rect -4886 456556 588810 456718
rect -8726 454274 592650 454436
rect -8726 454038 -7734 454274
rect -7498 454038 -7414 454274
rect -7178 454038 12986 454274
rect 13222 454038 13306 454274
rect 13542 454038 32986 454274
rect 33222 454038 33306 454274
rect 33542 454038 52986 454274
rect 53222 454038 53306 454274
rect 53542 454038 72986 454274
rect 73222 454038 73306 454274
rect 73542 454038 92986 454274
rect 93222 454038 93306 454274
rect 93542 454038 112986 454274
rect 113222 454038 113306 454274
rect 113542 454038 132986 454274
rect 133222 454038 133306 454274
rect 133542 454038 152986 454274
rect 153222 454038 153306 454274
rect 153542 454038 172986 454274
rect 173222 454038 173306 454274
rect 173542 454038 192986 454274
rect 193222 454038 193306 454274
rect 193542 454038 352986 454274
rect 353222 454038 353306 454274
rect 353542 454038 372986 454274
rect 373222 454038 373306 454274
rect 373542 454038 392986 454274
rect 393222 454038 393306 454274
rect 393542 454038 552986 454274
rect 553222 454038 553306 454274
rect 553542 454038 572986 454274
rect 573222 454038 573306 454274
rect 573542 454038 591102 454274
rect 591338 454038 591422 454274
rect 591658 454038 592650 454274
rect -8726 453876 592650 454038
rect -2966 453294 586890 453456
rect -2966 453058 -2934 453294
rect -2698 453058 -2614 453294
rect -2378 453058 11826 453294
rect 12062 453058 12146 453294
rect 12382 453058 31826 453294
rect 32062 453058 32146 453294
rect 32382 453058 51826 453294
rect 52062 453058 52146 453294
rect 52382 453058 71826 453294
rect 72062 453058 72146 453294
rect 72382 453058 91826 453294
rect 92062 453058 92146 453294
rect 92382 453058 111826 453294
rect 112062 453058 112146 453294
rect 112382 453058 131826 453294
rect 132062 453058 132146 453294
rect 132382 453058 151826 453294
rect 152062 453058 152146 453294
rect 152382 453058 171826 453294
rect 172062 453058 172146 453294
rect 172382 453058 191826 453294
rect 192062 453058 192146 453294
rect 192382 453058 351826 453294
rect 352062 453058 352146 453294
rect 352382 453058 371826 453294
rect 372062 453058 372146 453294
rect 372382 453058 391826 453294
rect 392062 453058 392146 453294
rect 392382 453058 551826 453294
rect 552062 453058 552146 453294
rect 552382 453058 571826 453294
rect 572062 453058 572146 453294
rect 572382 453058 586302 453294
rect 586538 453058 586622 453294
rect 586858 453058 586890 453294
rect -2966 452896 586890 453058
rect -6806 450614 590730 450776
rect -6806 450378 -5814 450614
rect -5578 450378 -5494 450614
rect -5258 450378 9266 450614
rect 9502 450378 9586 450614
rect 9822 450378 169266 450614
rect 169502 450378 169586 450614
rect 169822 450378 189266 450614
rect 189502 450378 189586 450614
rect 189822 450378 209266 450614
rect 209502 450378 209586 450614
rect 209822 450378 229266 450614
rect 229502 450378 229586 450614
rect 229822 450378 249266 450614
rect 249502 450378 249586 450614
rect 249822 450378 269266 450614
rect 269502 450378 269586 450614
rect 269822 450378 289266 450614
rect 289502 450378 289586 450614
rect 289822 450378 309266 450614
rect 309502 450378 309586 450614
rect 309822 450378 329266 450614
rect 329502 450378 329586 450614
rect 329822 450378 349266 450614
rect 349502 450378 349586 450614
rect 349822 450378 369266 450614
rect 369502 450378 369586 450614
rect 369822 450378 389266 450614
rect 389502 450378 389586 450614
rect 389822 450378 409266 450614
rect 409502 450378 409586 450614
rect 409822 450378 429266 450614
rect 429502 450378 429586 450614
rect 429822 450378 449266 450614
rect 449502 450378 449586 450614
rect 449822 450378 469266 450614
rect 469502 450378 469586 450614
rect 469822 450378 489266 450614
rect 489502 450378 489586 450614
rect 489822 450378 509266 450614
rect 509502 450378 509586 450614
rect 509822 450378 529266 450614
rect 529502 450378 529586 450614
rect 529822 450378 549266 450614
rect 549502 450378 549586 450614
rect 549822 450378 569266 450614
rect 569502 450378 569586 450614
rect 569822 450378 589182 450614
rect 589418 450378 589502 450614
rect 589738 450378 590730 450614
rect -6806 450216 590730 450378
rect -4886 446954 588810 447116
rect -4886 446718 -3894 446954
rect -3658 446718 -3574 446954
rect -3338 446718 5546 446954
rect 5782 446718 5866 446954
rect 6102 446718 25546 446954
rect 25782 446718 25866 446954
rect 26102 446718 185546 446954
rect 185782 446718 185866 446954
rect 186102 446718 205546 446954
rect 205782 446718 205866 446954
rect 206102 446718 225546 446954
rect 225782 446718 225866 446954
rect 226102 446718 245546 446954
rect 245782 446718 245866 446954
rect 246102 446718 265546 446954
rect 265782 446718 265866 446954
rect 266102 446718 285546 446954
rect 285782 446718 285866 446954
rect 286102 446718 305546 446954
rect 305782 446718 305866 446954
rect 306102 446718 325546 446954
rect 325782 446718 325866 446954
rect 326102 446718 345546 446954
rect 345782 446718 345866 446954
rect 346102 446718 365546 446954
rect 365782 446718 365866 446954
rect 366102 446718 385546 446954
rect 385782 446718 385866 446954
rect 386102 446718 405546 446954
rect 405782 446718 405866 446954
rect 406102 446718 425546 446954
rect 425782 446718 425866 446954
rect 426102 446718 445546 446954
rect 445782 446718 445866 446954
rect 446102 446718 465546 446954
rect 465782 446718 465866 446954
rect 466102 446718 485546 446954
rect 485782 446718 485866 446954
rect 486102 446718 505546 446954
rect 505782 446718 505866 446954
rect 506102 446718 525546 446954
rect 525782 446718 525866 446954
rect 526102 446718 545546 446954
rect 545782 446718 545866 446954
rect 546102 446718 565546 446954
rect 565782 446718 565866 446954
rect 566102 446718 587262 446954
rect 587498 446718 587582 446954
rect 587818 446718 588810 446954
rect -4886 446556 588810 446718
rect -8726 444274 592650 444436
rect -8726 444038 -8694 444274
rect -8458 444038 -8374 444274
rect -8138 444038 22986 444274
rect 23222 444038 23306 444274
rect 23542 444038 182986 444274
rect 183222 444038 183306 444274
rect 183542 444038 202986 444274
rect 203222 444038 203306 444274
rect 203542 444038 222986 444274
rect 223222 444038 223306 444274
rect 223542 444038 242986 444274
rect 243222 444038 243306 444274
rect 243542 444038 262986 444274
rect 263222 444038 263306 444274
rect 263542 444038 282986 444274
rect 283222 444038 283306 444274
rect 283542 444038 302986 444274
rect 303222 444038 303306 444274
rect 303542 444038 322986 444274
rect 323222 444038 323306 444274
rect 323542 444038 342986 444274
rect 343222 444038 343306 444274
rect 343542 444038 362986 444274
rect 363222 444038 363306 444274
rect 363542 444038 382986 444274
rect 383222 444038 383306 444274
rect 383542 444038 402986 444274
rect 403222 444038 403306 444274
rect 403542 444038 422986 444274
rect 423222 444038 423306 444274
rect 423542 444038 442986 444274
rect 443222 444038 443306 444274
rect 443542 444038 462986 444274
rect 463222 444038 463306 444274
rect 463542 444038 482986 444274
rect 483222 444038 483306 444274
rect 483542 444038 502986 444274
rect 503222 444038 503306 444274
rect 503542 444038 522986 444274
rect 523222 444038 523306 444274
rect 523542 444038 542986 444274
rect 543222 444038 543306 444274
rect 543542 444038 562986 444274
rect 563222 444038 563306 444274
rect 563542 444038 592062 444274
rect 592298 444038 592382 444274
rect 592618 444038 592650 444274
rect -8726 443876 592650 444038
rect -2966 443294 586890 443456
rect -2966 443058 -1974 443294
rect -1738 443058 -1654 443294
rect -1418 443058 1826 443294
rect 2062 443058 2146 443294
rect 2382 443058 21826 443294
rect 22062 443058 22146 443294
rect 22382 443058 31008 443294
rect 31244 443058 165376 443294
rect 165612 443058 181826 443294
rect 182062 443058 182146 443294
rect 182382 443058 201826 443294
rect 202062 443058 202146 443294
rect 202382 443058 221826 443294
rect 222062 443058 222146 443294
rect 222382 443058 241826 443294
rect 242062 443058 242146 443294
rect 242382 443058 261826 443294
rect 262062 443058 262146 443294
rect 262382 443058 281826 443294
rect 282062 443058 282146 443294
rect 282382 443058 301826 443294
rect 302062 443058 302146 443294
rect 302382 443058 321826 443294
rect 322062 443058 322146 443294
rect 322382 443058 341826 443294
rect 342062 443058 342146 443294
rect 342382 443058 361826 443294
rect 362062 443058 362146 443294
rect 362382 443058 381826 443294
rect 382062 443058 382146 443294
rect 382382 443058 401826 443294
rect 402062 443058 402146 443294
rect 402382 443058 421826 443294
rect 422062 443058 422146 443294
rect 422382 443058 441826 443294
rect 442062 443058 442146 443294
rect 442382 443058 461826 443294
rect 462062 443058 462146 443294
rect 462382 443058 481826 443294
rect 482062 443058 482146 443294
rect 482382 443058 501826 443294
rect 502062 443058 502146 443294
rect 502382 443058 521826 443294
rect 522062 443058 522146 443294
rect 522382 443058 541826 443294
rect 542062 443058 542146 443294
rect 542382 443058 561826 443294
rect 562062 443058 562146 443294
rect 562382 443058 581826 443294
rect 582062 443058 582146 443294
rect 582382 443058 585342 443294
rect 585578 443058 585662 443294
rect 585898 443058 586890 443294
rect -2966 442896 586890 443058
rect -6806 440614 590730 440776
rect -6806 440378 -6774 440614
rect -6538 440378 -6454 440614
rect -6218 440378 19266 440614
rect 19502 440378 19586 440614
rect 19822 440378 179266 440614
rect 179502 440378 179586 440614
rect 179822 440378 199266 440614
rect 199502 440378 199586 440614
rect 199822 440378 219266 440614
rect 219502 440378 219586 440614
rect 219822 440378 239266 440614
rect 239502 440378 239586 440614
rect 239822 440378 259266 440614
rect 259502 440378 259586 440614
rect 259822 440378 279266 440614
rect 279502 440378 279586 440614
rect 279822 440378 299266 440614
rect 299502 440378 299586 440614
rect 299822 440378 319266 440614
rect 319502 440378 319586 440614
rect 319822 440378 339266 440614
rect 339502 440378 339586 440614
rect 339822 440378 359266 440614
rect 359502 440378 359586 440614
rect 359822 440378 379266 440614
rect 379502 440378 379586 440614
rect 379822 440378 399266 440614
rect 399502 440378 399586 440614
rect 399822 440378 419266 440614
rect 419502 440378 419586 440614
rect 419822 440378 439266 440614
rect 439502 440378 439586 440614
rect 439822 440378 459266 440614
rect 459502 440378 459586 440614
rect 459822 440378 479266 440614
rect 479502 440378 479586 440614
rect 479822 440378 499266 440614
rect 499502 440378 499586 440614
rect 499822 440378 519266 440614
rect 519502 440378 519586 440614
rect 519822 440378 539266 440614
rect 539502 440378 539586 440614
rect 539822 440378 559266 440614
rect 559502 440378 559586 440614
rect 559822 440378 579266 440614
rect 579502 440378 579586 440614
rect 579822 440378 590142 440614
rect 590378 440378 590462 440614
rect 590698 440378 590730 440614
rect -6806 440216 590730 440378
rect -4886 436954 588810 437116
rect -4886 436718 -4854 436954
rect -4618 436718 -4534 436954
rect -4298 436718 15546 436954
rect 15782 436718 15866 436954
rect 16102 436718 175546 436954
rect 175782 436718 175866 436954
rect 176102 436718 195546 436954
rect 195782 436718 195866 436954
rect 196102 436718 215546 436954
rect 215782 436718 215866 436954
rect 216102 436718 235546 436954
rect 235782 436718 235866 436954
rect 236102 436718 255546 436954
rect 255782 436718 255866 436954
rect 256102 436718 275546 436954
rect 275782 436718 275866 436954
rect 276102 436718 295546 436954
rect 295782 436718 295866 436954
rect 296102 436718 315546 436954
rect 315782 436718 315866 436954
rect 316102 436718 335546 436954
rect 335782 436718 335866 436954
rect 336102 436718 355546 436954
rect 355782 436718 355866 436954
rect 356102 436718 375546 436954
rect 375782 436718 375866 436954
rect 376102 436718 395546 436954
rect 395782 436718 395866 436954
rect 396102 436718 415546 436954
rect 415782 436718 415866 436954
rect 416102 436718 435546 436954
rect 435782 436718 435866 436954
rect 436102 436718 455546 436954
rect 455782 436718 455866 436954
rect 456102 436718 475546 436954
rect 475782 436718 475866 436954
rect 476102 436718 495546 436954
rect 495782 436718 495866 436954
rect 496102 436718 515546 436954
rect 515782 436718 515866 436954
rect 516102 436718 535546 436954
rect 535782 436718 535866 436954
rect 536102 436718 555546 436954
rect 555782 436718 555866 436954
rect 556102 436718 575546 436954
rect 575782 436718 575866 436954
rect 576102 436718 588222 436954
rect 588458 436718 588542 436954
rect 588778 436718 588810 436954
rect -4886 436556 588810 436718
rect -8726 434274 592650 434436
rect -8726 434038 -7734 434274
rect -7498 434038 -7414 434274
rect -7178 434038 12986 434274
rect 13222 434038 13306 434274
rect 13542 434038 172986 434274
rect 173222 434038 173306 434274
rect 173542 434038 192986 434274
rect 193222 434038 193306 434274
rect 193542 434038 212986 434274
rect 213222 434038 213306 434274
rect 213542 434038 232986 434274
rect 233222 434038 233306 434274
rect 233542 434038 252986 434274
rect 253222 434038 253306 434274
rect 253542 434038 272986 434274
rect 273222 434038 273306 434274
rect 273542 434038 292986 434274
rect 293222 434038 293306 434274
rect 293542 434038 312986 434274
rect 313222 434038 313306 434274
rect 313542 434038 332986 434274
rect 333222 434038 333306 434274
rect 333542 434038 352986 434274
rect 353222 434038 353306 434274
rect 353542 434038 372986 434274
rect 373222 434038 373306 434274
rect 373542 434038 392986 434274
rect 393222 434038 393306 434274
rect 393542 434038 412986 434274
rect 413222 434038 413306 434274
rect 413542 434038 432986 434274
rect 433222 434038 433306 434274
rect 433542 434038 452986 434274
rect 453222 434038 453306 434274
rect 453542 434038 472986 434274
rect 473222 434038 473306 434274
rect 473542 434038 492986 434274
rect 493222 434038 493306 434274
rect 493542 434038 512986 434274
rect 513222 434038 513306 434274
rect 513542 434038 532986 434274
rect 533222 434038 533306 434274
rect 533542 434038 552986 434274
rect 553222 434038 553306 434274
rect 553542 434038 572986 434274
rect 573222 434038 573306 434274
rect 573542 434038 591102 434274
rect 591338 434038 591422 434274
rect 591658 434038 592650 434274
rect -8726 433876 592650 434038
rect -2966 433294 586890 433456
rect -2966 433058 -2934 433294
rect -2698 433058 -2614 433294
rect -2378 433058 11826 433294
rect 12062 433058 12146 433294
rect 12382 433058 30328 433294
rect 30564 433058 166056 433294
rect 166292 433058 171826 433294
rect 172062 433058 172146 433294
rect 172382 433058 191826 433294
rect 192062 433058 192146 433294
rect 192382 433058 211826 433294
rect 212062 433058 212146 433294
rect 212382 433058 231826 433294
rect 232062 433058 232146 433294
rect 232382 433058 251826 433294
rect 252062 433058 252146 433294
rect 252382 433058 271826 433294
rect 272062 433058 272146 433294
rect 272382 433058 291826 433294
rect 292062 433058 292146 433294
rect 292382 433058 311826 433294
rect 312062 433058 312146 433294
rect 312382 433058 331826 433294
rect 332062 433058 332146 433294
rect 332382 433058 351826 433294
rect 352062 433058 352146 433294
rect 352382 433058 371826 433294
rect 372062 433058 372146 433294
rect 372382 433058 391826 433294
rect 392062 433058 392146 433294
rect 392382 433058 411826 433294
rect 412062 433058 412146 433294
rect 412382 433058 431826 433294
rect 432062 433058 432146 433294
rect 432382 433058 451826 433294
rect 452062 433058 452146 433294
rect 452382 433058 471826 433294
rect 472062 433058 472146 433294
rect 472382 433058 491826 433294
rect 492062 433058 492146 433294
rect 492382 433058 511826 433294
rect 512062 433058 512146 433294
rect 512382 433058 531826 433294
rect 532062 433058 532146 433294
rect 532382 433058 551826 433294
rect 552062 433058 552146 433294
rect 552382 433058 571826 433294
rect 572062 433058 572146 433294
rect 572382 433058 586302 433294
rect 586538 433058 586622 433294
rect 586858 433058 586890 433294
rect -2966 432896 586890 433058
rect -6806 430614 590730 430776
rect -6806 430378 -5814 430614
rect -5578 430378 -5494 430614
rect -5258 430378 9266 430614
rect 9502 430378 9586 430614
rect 9822 430378 169266 430614
rect 169502 430378 169586 430614
rect 169822 430378 189266 430614
rect 189502 430378 189586 430614
rect 189822 430378 209266 430614
rect 209502 430378 209586 430614
rect 209822 430378 229266 430614
rect 229502 430378 229586 430614
rect 229822 430378 249266 430614
rect 249502 430378 249586 430614
rect 249822 430378 269266 430614
rect 269502 430378 269586 430614
rect 269822 430378 289266 430614
rect 289502 430378 289586 430614
rect 289822 430378 309266 430614
rect 309502 430378 309586 430614
rect 309822 430378 329266 430614
rect 329502 430378 329586 430614
rect 329822 430378 349266 430614
rect 349502 430378 349586 430614
rect 349822 430378 369266 430614
rect 369502 430378 369586 430614
rect 369822 430378 389266 430614
rect 389502 430378 389586 430614
rect 389822 430378 409266 430614
rect 409502 430378 409586 430614
rect 409822 430378 429266 430614
rect 429502 430378 429586 430614
rect 429822 430378 449266 430614
rect 449502 430378 449586 430614
rect 449822 430378 469266 430614
rect 469502 430378 469586 430614
rect 469822 430378 489266 430614
rect 489502 430378 489586 430614
rect 489822 430378 509266 430614
rect 509502 430378 509586 430614
rect 509822 430378 529266 430614
rect 529502 430378 529586 430614
rect 529822 430378 549266 430614
rect 549502 430378 549586 430614
rect 549822 430378 569266 430614
rect 569502 430378 569586 430614
rect 569822 430378 589182 430614
rect 589418 430378 589502 430614
rect 589738 430378 590730 430614
rect -6806 430216 590730 430378
rect -4886 426954 588810 427116
rect -4886 426718 -3894 426954
rect -3658 426718 -3574 426954
rect -3338 426718 5546 426954
rect 5782 426718 5866 426954
rect 6102 426718 25546 426954
rect 25782 426718 25866 426954
rect 26102 426718 185546 426954
rect 185782 426718 185866 426954
rect 186102 426718 205546 426954
rect 205782 426718 205866 426954
rect 206102 426718 225546 426954
rect 225782 426718 225866 426954
rect 226102 426718 245546 426954
rect 245782 426718 245866 426954
rect 246102 426718 265546 426954
rect 265782 426718 265866 426954
rect 266102 426718 285546 426954
rect 285782 426718 285866 426954
rect 286102 426718 305546 426954
rect 305782 426718 305866 426954
rect 306102 426718 325546 426954
rect 325782 426718 325866 426954
rect 326102 426718 345546 426954
rect 345782 426718 345866 426954
rect 346102 426718 365546 426954
rect 365782 426718 365866 426954
rect 366102 426718 385546 426954
rect 385782 426718 385866 426954
rect 386102 426718 405546 426954
rect 405782 426718 405866 426954
rect 406102 426718 425546 426954
rect 425782 426718 425866 426954
rect 426102 426718 445546 426954
rect 445782 426718 445866 426954
rect 446102 426718 465546 426954
rect 465782 426718 465866 426954
rect 466102 426718 485546 426954
rect 485782 426718 485866 426954
rect 486102 426718 505546 426954
rect 505782 426718 505866 426954
rect 506102 426718 525546 426954
rect 525782 426718 525866 426954
rect 526102 426718 545546 426954
rect 545782 426718 545866 426954
rect 546102 426718 565546 426954
rect 565782 426718 565866 426954
rect 566102 426718 587262 426954
rect 587498 426718 587582 426954
rect 587818 426718 588810 426954
rect -4886 426556 588810 426718
rect -8726 424274 592650 424436
rect -8726 424038 -8694 424274
rect -8458 424038 -8374 424274
rect -8138 424038 22986 424274
rect 23222 424038 23306 424274
rect 23542 424038 182986 424274
rect 183222 424038 183306 424274
rect 183542 424038 202986 424274
rect 203222 424038 203306 424274
rect 203542 424038 222986 424274
rect 223222 424038 223306 424274
rect 223542 424038 242986 424274
rect 243222 424038 243306 424274
rect 243542 424038 262986 424274
rect 263222 424038 263306 424274
rect 263542 424038 282986 424274
rect 283222 424038 283306 424274
rect 283542 424038 302986 424274
rect 303222 424038 303306 424274
rect 303542 424038 322986 424274
rect 323222 424038 323306 424274
rect 323542 424038 342986 424274
rect 343222 424038 343306 424274
rect 343542 424038 362986 424274
rect 363222 424038 363306 424274
rect 363542 424038 382986 424274
rect 383222 424038 383306 424274
rect 383542 424038 402986 424274
rect 403222 424038 403306 424274
rect 403542 424038 422986 424274
rect 423222 424038 423306 424274
rect 423542 424038 442986 424274
rect 443222 424038 443306 424274
rect 443542 424038 462986 424274
rect 463222 424038 463306 424274
rect 463542 424038 482986 424274
rect 483222 424038 483306 424274
rect 483542 424038 502986 424274
rect 503222 424038 503306 424274
rect 503542 424038 522986 424274
rect 523222 424038 523306 424274
rect 523542 424038 542986 424274
rect 543222 424038 543306 424274
rect 543542 424038 562986 424274
rect 563222 424038 563306 424274
rect 563542 424038 592062 424274
rect 592298 424038 592382 424274
rect 592618 424038 592650 424274
rect -8726 423876 592650 424038
rect -2966 423294 586890 423456
rect -2966 423058 -1974 423294
rect -1738 423058 -1654 423294
rect -1418 423058 1826 423294
rect 2062 423058 2146 423294
rect 2382 423058 21826 423294
rect 22062 423058 22146 423294
rect 22382 423058 31008 423294
rect 31244 423058 165376 423294
rect 165612 423058 181826 423294
rect 182062 423058 182146 423294
rect 182382 423058 201826 423294
rect 202062 423058 202146 423294
rect 202382 423058 221826 423294
rect 222062 423058 222146 423294
rect 222382 423058 241826 423294
rect 242062 423058 242146 423294
rect 242382 423058 261826 423294
rect 262062 423058 262146 423294
rect 262382 423058 281826 423294
rect 282062 423058 282146 423294
rect 282382 423058 301826 423294
rect 302062 423058 302146 423294
rect 302382 423058 321826 423294
rect 322062 423058 322146 423294
rect 322382 423058 341826 423294
rect 342062 423058 342146 423294
rect 342382 423058 361826 423294
rect 362062 423058 362146 423294
rect 362382 423058 381826 423294
rect 382062 423058 382146 423294
rect 382382 423058 401826 423294
rect 402062 423058 402146 423294
rect 402382 423058 421826 423294
rect 422062 423058 422146 423294
rect 422382 423058 441826 423294
rect 442062 423058 442146 423294
rect 442382 423058 461826 423294
rect 462062 423058 462146 423294
rect 462382 423058 481826 423294
rect 482062 423058 482146 423294
rect 482382 423058 501826 423294
rect 502062 423058 502146 423294
rect 502382 423058 521826 423294
rect 522062 423058 522146 423294
rect 522382 423058 541826 423294
rect 542062 423058 542146 423294
rect 542382 423058 561826 423294
rect 562062 423058 562146 423294
rect 562382 423058 581826 423294
rect 582062 423058 582146 423294
rect 582382 423058 585342 423294
rect 585578 423058 585662 423294
rect 585898 423058 586890 423294
rect -2966 422896 586890 423058
rect -6806 420614 590730 420776
rect -6806 420378 -6774 420614
rect -6538 420378 -6454 420614
rect -6218 420378 19266 420614
rect 19502 420378 19586 420614
rect 19822 420378 179266 420614
rect 179502 420378 179586 420614
rect 179822 420378 559266 420614
rect 559502 420378 559586 420614
rect 559822 420378 579266 420614
rect 579502 420378 579586 420614
rect 579822 420378 590142 420614
rect 590378 420378 590462 420614
rect 590698 420378 590730 420614
rect -6806 420216 590730 420378
rect -4886 416954 588810 417116
rect -4886 416718 -4854 416954
rect -4618 416718 -4534 416954
rect -4298 416718 15546 416954
rect 15782 416718 15866 416954
rect 16102 416718 175546 416954
rect 175782 416718 175866 416954
rect 176102 416718 195546 416954
rect 195782 416718 195866 416954
rect 196102 416718 575546 416954
rect 575782 416718 575866 416954
rect 576102 416718 588222 416954
rect 588458 416718 588542 416954
rect 588778 416718 588810 416954
rect -4886 416556 588810 416718
rect -8726 414274 592650 414436
rect -8726 414038 -7734 414274
rect -7498 414038 -7414 414274
rect -7178 414038 12986 414274
rect 13222 414038 13306 414274
rect 13542 414038 172986 414274
rect 173222 414038 173306 414274
rect 173542 414038 192986 414274
rect 193222 414038 193306 414274
rect 193542 414038 572986 414274
rect 573222 414038 573306 414274
rect 573542 414038 591102 414274
rect 591338 414038 591422 414274
rect 591658 414038 592650 414274
rect -8726 413876 592650 414038
rect -2966 413294 586890 413456
rect -2966 413058 -2934 413294
rect -2698 413058 -2614 413294
rect -2378 413058 11826 413294
rect 12062 413058 12146 413294
rect 12382 413058 30328 413294
rect 30564 413058 166056 413294
rect 166292 413058 171826 413294
rect 172062 413058 172146 413294
rect 172382 413058 191826 413294
rect 192062 413058 192146 413294
rect 192382 413058 219610 413294
rect 219846 413058 250330 413294
rect 250566 413058 281050 413294
rect 281286 413058 311770 413294
rect 312006 413058 342490 413294
rect 342726 413058 373210 413294
rect 373446 413058 403930 413294
rect 404166 413058 434650 413294
rect 434886 413058 465370 413294
rect 465606 413058 496090 413294
rect 496326 413058 526810 413294
rect 527046 413058 571826 413294
rect 572062 413058 572146 413294
rect 572382 413058 586302 413294
rect 586538 413058 586622 413294
rect 586858 413058 586890 413294
rect -2966 412896 586890 413058
rect -6806 410614 590730 410776
rect -6806 410378 -5814 410614
rect -5578 410378 -5494 410614
rect -5258 410378 9266 410614
rect 9502 410378 9586 410614
rect 9822 410378 169266 410614
rect 169502 410378 169586 410614
rect 169822 410378 189266 410614
rect 189502 410378 189586 410614
rect 189822 410378 569266 410614
rect 569502 410378 569586 410614
rect 569822 410378 589182 410614
rect 589418 410378 589502 410614
rect 589738 410378 590730 410614
rect -6806 410216 590730 410378
rect -4886 406954 588810 407116
rect -4886 406718 -3894 406954
rect -3658 406718 -3574 406954
rect -3338 406718 5546 406954
rect 5782 406718 5866 406954
rect 6102 406718 25546 406954
rect 25782 406718 25866 406954
rect 26102 406718 185546 406954
rect 185782 406718 185866 406954
rect 186102 406718 565546 406954
rect 565782 406718 565866 406954
rect 566102 406718 587262 406954
rect 587498 406718 587582 406954
rect 587818 406718 588810 406954
rect -4886 406556 588810 406718
rect -8726 404274 592650 404436
rect -8726 404038 -8694 404274
rect -8458 404038 -8374 404274
rect -8138 404038 22986 404274
rect 23222 404038 23306 404274
rect 23542 404038 182986 404274
rect 183222 404038 183306 404274
rect 183542 404038 562986 404274
rect 563222 404038 563306 404274
rect 563542 404038 592062 404274
rect 592298 404038 592382 404274
rect 592618 404038 592650 404274
rect -8726 403876 592650 404038
rect -2966 403294 586890 403456
rect -2966 403058 -1974 403294
rect -1738 403058 -1654 403294
rect -1418 403058 1826 403294
rect 2062 403058 2146 403294
rect 2382 403058 21826 403294
rect 22062 403058 22146 403294
rect 22382 403058 31008 403294
rect 31244 403058 165376 403294
rect 165612 403058 181826 403294
rect 182062 403058 182146 403294
rect 182382 403058 204250 403294
rect 204486 403058 234970 403294
rect 235206 403058 265690 403294
rect 265926 403058 296410 403294
rect 296646 403058 327130 403294
rect 327366 403058 357850 403294
rect 358086 403058 388570 403294
rect 388806 403058 419290 403294
rect 419526 403058 450010 403294
rect 450246 403058 480730 403294
rect 480966 403058 511450 403294
rect 511686 403058 542170 403294
rect 542406 403058 561826 403294
rect 562062 403058 562146 403294
rect 562382 403058 581826 403294
rect 582062 403058 582146 403294
rect 582382 403058 585342 403294
rect 585578 403058 585662 403294
rect 585898 403058 586890 403294
rect -2966 402896 586890 403058
rect -6806 400614 590730 400776
rect -6806 400378 -6774 400614
rect -6538 400378 -6454 400614
rect -6218 400378 19266 400614
rect 19502 400378 19586 400614
rect 19822 400378 179266 400614
rect 179502 400378 179586 400614
rect 179822 400378 559266 400614
rect 559502 400378 559586 400614
rect 559822 400378 579266 400614
rect 579502 400378 579586 400614
rect 579822 400378 590142 400614
rect 590378 400378 590462 400614
rect 590698 400378 590730 400614
rect -6806 400216 590730 400378
rect -4886 396954 588810 397116
rect -4886 396718 -4854 396954
rect -4618 396718 -4534 396954
rect -4298 396718 15546 396954
rect 15782 396718 15866 396954
rect 16102 396718 175546 396954
rect 175782 396718 175866 396954
rect 176102 396718 195546 396954
rect 195782 396718 195866 396954
rect 196102 396718 575546 396954
rect 575782 396718 575866 396954
rect 576102 396718 588222 396954
rect 588458 396718 588542 396954
rect 588778 396718 588810 396954
rect -4886 396556 588810 396718
rect -8726 394274 592650 394436
rect -8726 394038 -7734 394274
rect -7498 394038 -7414 394274
rect -7178 394038 12986 394274
rect 13222 394038 13306 394274
rect 13542 394038 172986 394274
rect 173222 394038 173306 394274
rect 173542 394038 192986 394274
rect 193222 394038 193306 394274
rect 193542 394038 572986 394274
rect 573222 394038 573306 394274
rect 573542 394038 591102 394274
rect 591338 394038 591422 394274
rect 591658 394038 592650 394274
rect -8726 393876 592650 394038
rect -2966 393294 586890 393456
rect -2966 393058 -2934 393294
rect -2698 393058 -2614 393294
rect -2378 393058 11826 393294
rect 12062 393058 12146 393294
rect 12382 393058 30328 393294
rect 30564 393058 166056 393294
rect 166292 393058 171826 393294
rect 172062 393058 172146 393294
rect 172382 393058 191826 393294
rect 192062 393058 192146 393294
rect 192382 393058 219610 393294
rect 219846 393058 250330 393294
rect 250566 393058 281050 393294
rect 281286 393058 311770 393294
rect 312006 393058 342490 393294
rect 342726 393058 373210 393294
rect 373446 393058 403930 393294
rect 404166 393058 434650 393294
rect 434886 393058 465370 393294
rect 465606 393058 496090 393294
rect 496326 393058 526810 393294
rect 527046 393058 571826 393294
rect 572062 393058 572146 393294
rect 572382 393058 586302 393294
rect 586538 393058 586622 393294
rect 586858 393058 586890 393294
rect -2966 392896 586890 393058
rect -6806 390614 590730 390776
rect -6806 390378 -5814 390614
rect -5578 390378 -5494 390614
rect -5258 390378 9266 390614
rect 9502 390378 9586 390614
rect 9822 390378 169266 390614
rect 169502 390378 169586 390614
rect 169822 390378 189266 390614
rect 189502 390378 189586 390614
rect 189822 390378 569266 390614
rect 569502 390378 569586 390614
rect 569822 390378 589182 390614
rect 589418 390378 589502 390614
rect 589738 390378 590730 390614
rect -6806 390216 590730 390378
rect -4886 386954 588810 387116
rect -4886 386718 -3894 386954
rect -3658 386718 -3574 386954
rect -3338 386718 5546 386954
rect 5782 386718 5866 386954
rect 6102 386718 25546 386954
rect 25782 386718 25866 386954
rect 26102 386718 185546 386954
rect 185782 386718 185866 386954
rect 186102 386718 565546 386954
rect 565782 386718 565866 386954
rect 566102 386718 587262 386954
rect 587498 386718 587582 386954
rect 587818 386718 588810 386954
rect -4886 386556 588810 386718
rect -8726 384274 592650 384436
rect -8726 384038 -8694 384274
rect -8458 384038 -8374 384274
rect -8138 384038 22986 384274
rect 23222 384038 23306 384274
rect 23542 384038 182986 384274
rect 183222 384038 183306 384274
rect 183542 384038 562986 384274
rect 563222 384038 563306 384274
rect 563542 384038 592062 384274
rect 592298 384038 592382 384274
rect 592618 384038 592650 384274
rect -8726 383876 592650 384038
rect -2966 383294 586890 383456
rect -2966 383058 -1974 383294
rect -1738 383058 -1654 383294
rect -1418 383058 1826 383294
rect 2062 383058 2146 383294
rect 2382 383058 21826 383294
rect 22062 383058 22146 383294
rect 22382 383058 31008 383294
rect 31244 383058 165376 383294
rect 165612 383058 181826 383294
rect 182062 383058 182146 383294
rect 182382 383058 204250 383294
rect 204486 383058 234970 383294
rect 235206 383058 265690 383294
rect 265926 383058 296410 383294
rect 296646 383058 327130 383294
rect 327366 383058 357850 383294
rect 358086 383058 388570 383294
rect 388806 383058 419290 383294
rect 419526 383058 450010 383294
rect 450246 383058 480730 383294
rect 480966 383058 511450 383294
rect 511686 383058 542170 383294
rect 542406 383058 561826 383294
rect 562062 383058 562146 383294
rect 562382 383058 581826 383294
rect 582062 383058 582146 383294
rect 582382 383058 585342 383294
rect 585578 383058 585662 383294
rect 585898 383058 586890 383294
rect -2966 382896 586890 383058
rect -6806 380614 590730 380776
rect -6806 380378 -6774 380614
rect -6538 380378 -6454 380614
rect -6218 380378 19266 380614
rect 19502 380378 19586 380614
rect 19822 380378 179266 380614
rect 179502 380378 179586 380614
rect 179822 380378 559266 380614
rect 559502 380378 559586 380614
rect 559822 380378 579266 380614
rect 579502 380378 579586 380614
rect 579822 380378 590142 380614
rect 590378 380378 590462 380614
rect 590698 380378 590730 380614
rect -6806 380216 590730 380378
rect -4886 376954 588810 377116
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15546 376954
rect 15782 376718 15866 376954
rect 16102 376718 175546 376954
rect 175782 376718 175866 376954
rect 176102 376718 195546 376954
rect 195782 376718 195866 376954
rect 196102 376718 575546 376954
rect 575782 376718 575866 376954
rect 576102 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect -4886 376556 588810 376718
rect -8726 374274 592650 374436
rect -8726 374038 -7734 374274
rect -7498 374038 -7414 374274
rect -7178 374038 12986 374274
rect 13222 374038 13306 374274
rect 13542 374038 172986 374274
rect 173222 374038 173306 374274
rect 173542 374038 192986 374274
rect 193222 374038 193306 374274
rect 193542 374038 572986 374274
rect 573222 374038 573306 374274
rect 573542 374038 591102 374274
rect 591338 374038 591422 374274
rect 591658 374038 592650 374274
rect -8726 373876 592650 374038
rect -2966 373294 586890 373456
rect -2966 373058 -2934 373294
rect -2698 373058 -2614 373294
rect -2378 373058 11826 373294
rect 12062 373058 12146 373294
rect 12382 373058 30328 373294
rect 30564 373058 166056 373294
rect 166292 373058 171826 373294
rect 172062 373058 172146 373294
rect 172382 373058 191826 373294
rect 192062 373058 192146 373294
rect 192382 373058 219610 373294
rect 219846 373058 250330 373294
rect 250566 373058 281050 373294
rect 281286 373058 311770 373294
rect 312006 373058 342490 373294
rect 342726 373058 373210 373294
rect 373446 373058 403930 373294
rect 404166 373058 434650 373294
rect 434886 373058 465370 373294
rect 465606 373058 496090 373294
rect 496326 373058 526810 373294
rect 527046 373058 571826 373294
rect 572062 373058 572146 373294
rect 572382 373058 586302 373294
rect 586538 373058 586622 373294
rect 586858 373058 586890 373294
rect -2966 372896 586890 373058
rect -6806 370614 590730 370776
rect -6806 370378 -5814 370614
rect -5578 370378 -5494 370614
rect -5258 370378 9266 370614
rect 9502 370378 9586 370614
rect 9822 370378 169266 370614
rect 169502 370378 169586 370614
rect 169822 370378 189266 370614
rect 189502 370378 189586 370614
rect 189822 370378 569266 370614
rect 569502 370378 569586 370614
rect 569822 370378 589182 370614
rect 589418 370378 589502 370614
rect 589738 370378 590730 370614
rect -6806 370216 590730 370378
rect -4886 366954 588810 367116
rect -4886 366718 -3894 366954
rect -3658 366718 -3574 366954
rect -3338 366718 5546 366954
rect 5782 366718 5866 366954
rect 6102 366718 25546 366954
rect 25782 366718 25866 366954
rect 26102 366718 185546 366954
rect 185782 366718 185866 366954
rect 186102 366718 565546 366954
rect 565782 366718 565866 366954
rect 566102 366718 587262 366954
rect 587498 366718 587582 366954
rect 587818 366718 588810 366954
rect -4886 366556 588810 366718
rect -8726 364274 592650 364436
rect -8726 364038 -8694 364274
rect -8458 364038 -8374 364274
rect -8138 364038 22986 364274
rect 23222 364038 23306 364274
rect 23542 364038 182986 364274
rect 183222 364038 183306 364274
rect 183542 364038 562986 364274
rect 563222 364038 563306 364274
rect 563542 364038 592062 364274
rect 592298 364038 592382 364274
rect 592618 364038 592650 364274
rect -8726 363876 592650 364038
rect -2966 363294 586890 363456
rect -2966 363058 -1974 363294
rect -1738 363058 -1654 363294
rect -1418 363058 1826 363294
rect 2062 363058 2146 363294
rect 2382 363058 21826 363294
rect 22062 363058 22146 363294
rect 22382 363058 41826 363294
rect 42062 363058 42146 363294
rect 42382 363058 61826 363294
rect 62062 363058 62146 363294
rect 62382 363058 81826 363294
rect 82062 363058 82146 363294
rect 82382 363058 101826 363294
rect 102062 363058 102146 363294
rect 102382 363058 121826 363294
rect 122062 363058 122146 363294
rect 122382 363058 141826 363294
rect 142062 363058 142146 363294
rect 142382 363058 161826 363294
rect 162062 363058 162146 363294
rect 162382 363058 181826 363294
rect 182062 363058 182146 363294
rect 182382 363058 204250 363294
rect 204486 363058 234970 363294
rect 235206 363058 265690 363294
rect 265926 363058 296410 363294
rect 296646 363058 327130 363294
rect 327366 363058 357850 363294
rect 358086 363058 388570 363294
rect 388806 363058 419290 363294
rect 419526 363058 450010 363294
rect 450246 363058 480730 363294
rect 480966 363058 511450 363294
rect 511686 363058 542170 363294
rect 542406 363058 561826 363294
rect 562062 363058 562146 363294
rect 562382 363058 581826 363294
rect 582062 363058 582146 363294
rect 582382 363058 585342 363294
rect 585578 363058 585662 363294
rect 585898 363058 586890 363294
rect -2966 362896 586890 363058
rect -6806 360614 590730 360776
rect -6806 360378 -6774 360614
rect -6538 360378 -6454 360614
rect -6218 360378 19266 360614
rect 19502 360378 19586 360614
rect 19822 360378 39266 360614
rect 39502 360378 39586 360614
rect 39822 360378 59266 360614
rect 59502 360378 59586 360614
rect 59822 360378 79266 360614
rect 79502 360378 79586 360614
rect 79822 360378 99266 360614
rect 99502 360378 99586 360614
rect 99822 360378 119266 360614
rect 119502 360378 119586 360614
rect 119822 360378 139266 360614
rect 139502 360378 139586 360614
rect 139822 360378 159266 360614
rect 159502 360378 159586 360614
rect 159822 360378 179266 360614
rect 179502 360378 179586 360614
rect 179822 360378 559266 360614
rect 559502 360378 559586 360614
rect 559822 360378 579266 360614
rect 579502 360378 579586 360614
rect 579822 360378 590142 360614
rect 590378 360378 590462 360614
rect 590698 360378 590730 360614
rect -6806 360216 590730 360378
rect -4886 356954 588810 357116
rect -4886 356718 -4854 356954
rect -4618 356718 -4534 356954
rect -4298 356718 15546 356954
rect 15782 356718 15866 356954
rect 16102 356718 35546 356954
rect 35782 356718 35866 356954
rect 36102 356718 55546 356954
rect 55782 356718 55866 356954
rect 56102 356718 75546 356954
rect 75782 356718 75866 356954
rect 76102 356718 95546 356954
rect 95782 356718 95866 356954
rect 96102 356718 115546 356954
rect 115782 356718 115866 356954
rect 116102 356718 135546 356954
rect 135782 356718 135866 356954
rect 136102 356718 155546 356954
rect 155782 356718 155866 356954
rect 156102 356718 175546 356954
rect 175782 356718 175866 356954
rect 176102 356718 195546 356954
rect 195782 356718 195866 356954
rect 196102 356718 575546 356954
rect 575782 356718 575866 356954
rect 576102 356718 588222 356954
rect 588458 356718 588542 356954
rect 588778 356718 588810 356954
rect -4886 356556 588810 356718
rect -8726 354274 592650 354436
rect -8726 354038 -7734 354274
rect -7498 354038 -7414 354274
rect -7178 354038 12986 354274
rect 13222 354038 13306 354274
rect 13542 354038 32986 354274
rect 33222 354038 33306 354274
rect 33542 354038 52986 354274
rect 53222 354038 53306 354274
rect 53542 354038 72986 354274
rect 73222 354038 73306 354274
rect 73542 354038 92986 354274
rect 93222 354038 93306 354274
rect 93542 354038 112986 354274
rect 113222 354038 113306 354274
rect 113542 354038 132986 354274
rect 133222 354038 133306 354274
rect 133542 354038 152986 354274
rect 153222 354038 153306 354274
rect 153542 354038 172986 354274
rect 173222 354038 173306 354274
rect 173542 354038 192986 354274
rect 193222 354038 193306 354274
rect 193542 354038 572986 354274
rect 573222 354038 573306 354274
rect 573542 354038 591102 354274
rect 591338 354038 591422 354274
rect 591658 354038 592650 354274
rect -8726 353876 592650 354038
rect -2966 353294 586890 353456
rect -2966 353058 -2934 353294
rect -2698 353058 -2614 353294
rect -2378 353058 11826 353294
rect 12062 353058 12146 353294
rect 12382 353058 31826 353294
rect 32062 353058 32146 353294
rect 32382 353058 51826 353294
rect 52062 353058 52146 353294
rect 52382 353058 71826 353294
rect 72062 353058 72146 353294
rect 72382 353058 91826 353294
rect 92062 353058 92146 353294
rect 92382 353058 111826 353294
rect 112062 353058 112146 353294
rect 112382 353058 131826 353294
rect 132062 353058 132146 353294
rect 132382 353058 151826 353294
rect 152062 353058 152146 353294
rect 152382 353058 171826 353294
rect 172062 353058 172146 353294
rect 172382 353058 191826 353294
rect 192062 353058 192146 353294
rect 192382 353058 219610 353294
rect 219846 353058 250330 353294
rect 250566 353058 281050 353294
rect 281286 353058 311770 353294
rect 312006 353058 342490 353294
rect 342726 353058 373210 353294
rect 373446 353058 403930 353294
rect 404166 353058 434650 353294
rect 434886 353058 465370 353294
rect 465606 353058 496090 353294
rect 496326 353058 526810 353294
rect 527046 353058 571826 353294
rect 572062 353058 572146 353294
rect 572382 353058 586302 353294
rect 586538 353058 586622 353294
rect 586858 353058 586890 353294
rect -2966 352896 586890 353058
rect -6806 350614 590730 350776
rect -6806 350378 -5814 350614
rect -5578 350378 -5494 350614
rect -5258 350378 9266 350614
rect 9502 350378 9586 350614
rect 9822 350378 29266 350614
rect 29502 350378 29586 350614
rect 29822 350378 49266 350614
rect 49502 350378 49586 350614
rect 49822 350378 69266 350614
rect 69502 350378 69586 350614
rect 69822 350378 89266 350614
rect 89502 350378 89586 350614
rect 89822 350378 109266 350614
rect 109502 350378 109586 350614
rect 109822 350378 129266 350614
rect 129502 350378 129586 350614
rect 129822 350378 149266 350614
rect 149502 350378 149586 350614
rect 149822 350378 169266 350614
rect 169502 350378 169586 350614
rect 169822 350378 189266 350614
rect 189502 350378 189586 350614
rect 189822 350378 569266 350614
rect 569502 350378 569586 350614
rect 569822 350378 589182 350614
rect 589418 350378 589502 350614
rect 589738 350378 590730 350614
rect -6806 350216 590730 350378
rect -4886 346954 588810 347116
rect -4886 346718 -3894 346954
rect -3658 346718 -3574 346954
rect -3338 346718 5546 346954
rect 5782 346718 5866 346954
rect 6102 346718 25546 346954
rect 25782 346718 25866 346954
rect 26102 346718 45546 346954
rect 45782 346718 45866 346954
rect 46102 346718 65546 346954
rect 65782 346718 65866 346954
rect 66102 346718 85546 346954
rect 85782 346718 85866 346954
rect 86102 346718 105546 346954
rect 105782 346718 105866 346954
rect 106102 346718 125546 346954
rect 125782 346718 125866 346954
rect 126102 346718 145546 346954
rect 145782 346718 145866 346954
rect 146102 346718 165546 346954
rect 165782 346718 165866 346954
rect 166102 346718 185546 346954
rect 185782 346718 185866 346954
rect 186102 346718 565546 346954
rect 565782 346718 565866 346954
rect 566102 346718 587262 346954
rect 587498 346718 587582 346954
rect 587818 346718 588810 346954
rect -4886 346556 588810 346718
rect -8726 344274 592650 344436
rect -8726 344038 -8694 344274
rect -8458 344038 -8374 344274
rect -8138 344038 22986 344274
rect 23222 344038 23306 344274
rect 23542 344038 42986 344274
rect 43222 344038 43306 344274
rect 43542 344038 62986 344274
rect 63222 344038 63306 344274
rect 63542 344038 82986 344274
rect 83222 344038 83306 344274
rect 83542 344038 102986 344274
rect 103222 344038 103306 344274
rect 103542 344038 122986 344274
rect 123222 344038 123306 344274
rect 123542 344038 142986 344274
rect 143222 344038 143306 344274
rect 143542 344038 162986 344274
rect 163222 344038 163306 344274
rect 163542 344038 182986 344274
rect 183222 344038 183306 344274
rect 183542 344038 562986 344274
rect 563222 344038 563306 344274
rect 563542 344038 592062 344274
rect 592298 344038 592382 344274
rect 592618 344038 592650 344274
rect -8726 343876 592650 344038
rect -2966 343294 586890 343456
rect -2966 343058 -1974 343294
rect -1738 343058 -1654 343294
rect -1418 343058 1826 343294
rect 2062 343058 2146 343294
rect 2382 343058 21826 343294
rect 22062 343058 22146 343294
rect 22382 343058 41826 343294
rect 42062 343058 42146 343294
rect 42382 343058 61826 343294
rect 62062 343058 62146 343294
rect 62382 343058 81826 343294
rect 82062 343058 82146 343294
rect 82382 343058 101826 343294
rect 102062 343058 102146 343294
rect 102382 343058 121826 343294
rect 122062 343058 122146 343294
rect 122382 343058 141826 343294
rect 142062 343058 142146 343294
rect 142382 343058 161826 343294
rect 162062 343058 162146 343294
rect 162382 343058 181826 343294
rect 182062 343058 182146 343294
rect 182382 343058 204250 343294
rect 204486 343058 234970 343294
rect 235206 343058 265690 343294
rect 265926 343058 296410 343294
rect 296646 343058 327130 343294
rect 327366 343058 357850 343294
rect 358086 343058 388570 343294
rect 388806 343058 419290 343294
rect 419526 343058 450010 343294
rect 450246 343058 480730 343294
rect 480966 343058 511450 343294
rect 511686 343058 542170 343294
rect 542406 343058 561826 343294
rect 562062 343058 562146 343294
rect 562382 343058 581826 343294
rect 582062 343058 582146 343294
rect 582382 343058 585342 343294
rect 585578 343058 585662 343294
rect 585898 343058 586890 343294
rect -2966 342896 586890 343058
rect -6806 340614 590730 340776
rect -6806 340378 -6774 340614
rect -6538 340378 -6454 340614
rect -6218 340378 19266 340614
rect 19502 340378 19586 340614
rect 19822 340378 39266 340614
rect 39502 340378 39586 340614
rect 39822 340378 59266 340614
rect 59502 340378 59586 340614
rect 59822 340378 79266 340614
rect 79502 340378 79586 340614
rect 79822 340378 99266 340614
rect 99502 340378 99586 340614
rect 99822 340378 119266 340614
rect 119502 340378 119586 340614
rect 119822 340378 139266 340614
rect 139502 340378 139586 340614
rect 139822 340378 159266 340614
rect 159502 340378 159586 340614
rect 159822 340378 179266 340614
rect 179502 340378 179586 340614
rect 179822 340378 559266 340614
rect 559502 340378 559586 340614
rect 559822 340378 579266 340614
rect 579502 340378 579586 340614
rect 579822 340378 590142 340614
rect 590378 340378 590462 340614
rect 590698 340378 590730 340614
rect -6806 340216 590730 340378
rect -4886 336954 588810 337116
rect -4886 336718 -4854 336954
rect -4618 336718 -4534 336954
rect -4298 336718 15546 336954
rect 15782 336718 15866 336954
rect 16102 336718 175546 336954
rect 175782 336718 175866 336954
rect 176102 336718 195546 336954
rect 195782 336718 195866 336954
rect 196102 336718 575546 336954
rect 575782 336718 575866 336954
rect 576102 336718 588222 336954
rect 588458 336718 588542 336954
rect 588778 336718 588810 336954
rect -4886 336556 588810 336718
rect -8726 334274 592650 334436
rect -8726 334038 -7734 334274
rect -7498 334038 -7414 334274
rect -7178 334038 12986 334274
rect 13222 334038 13306 334274
rect 13542 334038 172986 334274
rect 173222 334038 173306 334274
rect 173542 334038 192986 334274
rect 193222 334038 193306 334274
rect 193542 334038 572986 334274
rect 573222 334038 573306 334274
rect 573542 334038 591102 334274
rect 591338 334038 591422 334274
rect 591658 334038 592650 334274
rect -8726 333876 592650 334038
rect -2966 333294 586890 333456
rect -2966 333058 -2934 333294
rect -2698 333058 -2614 333294
rect -2378 333058 11826 333294
rect 12062 333058 12146 333294
rect 12382 333058 30328 333294
rect 30564 333058 166056 333294
rect 166292 333058 171826 333294
rect 172062 333058 172146 333294
rect 172382 333058 191826 333294
rect 192062 333058 192146 333294
rect 192382 333058 219610 333294
rect 219846 333058 250330 333294
rect 250566 333058 281050 333294
rect 281286 333058 311770 333294
rect 312006 333058 342490 333294
rect 342726 333058 373210 333294
rect 373446 333058 403930 333294
rect 404166 333058 434650 333294
rect 434886 333058 465370 333294
rect 465606 333058 496090 333294
rect 496326 333058 526810 333294
rect 527046 333058 571826 333294
rect 572062 333058 572146 333294
rect 572382 333058 586302 333294
rect 586538 333058 586622 333294
rect 586858 333058 586890 333294
rect -2966 332896 586890 333058
rect -6806 330614 590730 330776
rect -6806 330378 -5814 330614
rect -5578 330378 -5494 330614
rect -5258 330378 9266 330614
rect 9502 330378 9586 330614
rect 9822 330378 169266 330614
rect 169502 330378 169586 330614
rect 169822 330378 189266 330614
rect 189502 330378 189586 330614
rect 189822 330378 569266 330614
rect 569502 330378 569586 330614
rect 569822 330378 589182 330614
rect 589418 330378 589502 330614
rect 589738 330378 590730 330614
rect -6806 330216 590730 330378
rect -4886 326954 588810 327116
rect -4886 326718 -3894 326954
rect -3658 326718 -3574 326954
rect -3338 326718 5546 326954
rect 5782 326718 5866 326954
rect 6102 326718 25546 326954
rect 25782 326718 25866 326954
rect 26102 326718 185546 326954
rect 185782 326718 185866 326954
rect 186102 326718 565546 326954
rect 565782 326718 565866 326954
rect 566102 326718 587262 326954
rect 587498 326718 587582 326954
rect 587818 326718 588810 326954
rect -4886 326556 588810 326718
rect -8726 324274 592650 324436
rect -8726 324038 -8694 324274
rect -8458 324038 -8374 324274
rect -8138 324038 22986 324274
rect 23222 324038 23306 324274
rect 23542 324038 182986 324274
rect 183222 324038 183306 324274
rect 183542 324038 562986 324274
rect 563222 324038 563306 324274
rect 563542 324038 592062 324274
rect 592298 324038 592382 324274
rect 592618 324038 592650 324274
rect -8726 323876 592650 324038
rect -2966 323294 586890 323456
rect -2966 323058 -1974 323294
rect -1738 323058 -1654 323294
rect -1418 323058 1826 323294
rect 2062 323058 2146 323294
rect 2382 323058 21826 323294
rect 22062 323058 22146 323294
rect 22382 323058 31008 323294
rect 31244 323058 165376 323294
rect 165612 323058 181826 323294
rect 182062 323058 182146 323294
rect 182382 323058 204250 323294
rect 204486 323058 234970 323294
rect 235206 323058 265690 323294
rect 265926 323058 296410 323294
rect 296646 323058 327130 323294
rect 327366 323058 357850 323294
rect 358086 323058 388570 323294
rect 388806 323058 419290 323294
rect 419526 323058 450010 323294
rect 450246 323058 480730 323294
rect 480966 323058 511450 323294
rect 511686 323058 542170 323294
rect 542406 323058 561826 323294
rect 562062 323058 562146 323294
rect 562382 323058 581826 323294
rect 582062 323058 582146 323294
rect 582382 323058 585342 323294
rect 585578 323058 585662 323294
rect 585898 323058 586890 323294
rect -2966 322896 586890 323058
rect -6806 320614 590730 320776
rect -6806 320378 -6774 320614
rect -6538 320378 -6454 320614
rect -6218 320378 19266 320614
rect 19502 320378 19586 320614
rect 19822 320378 179266 320614
rect 179502 320378 179586 320614
rect 179822 320378 559266 320614
rect 559502 320378 559586 320614
rect 559822 320378 579266 320614
rect 579502 320378 579586 320614
rect 579822 320378 590142 320614
rect 590378 320378 590462 320614
rect 590698 320378 590730 320614
rect -6806 320216 590730 320378
rect -4886 316954 588810 317116
rect -4886 316718 -4854 316954
rect -4618 316718 -4534 316954
rect -4298 316718 15546 316954
rect 15782 316718 15866 316954
rect 16102 316718 175546 316954
rect 175782 316718 175866 316954
rect 176102 316718 195546 316954
rect 195782 316718 195866 316954
rect 196102 316718 575546 316954
rect 575782 316718 575866 316954
rect 576102 316718 588222 316954
rect 588458 316718 588542 316954
rect 588778 316718 588810 316954
rect -4886 316556 588810 316718
rect -8726 314274 592650 314436
rect -8726 314038 -7734 314274
rect -7498 314038 -7414 314274
rect -7178 314038 12986 314274
rect 13222 314038 13306 314274
rect 13542 314038 172986 314274
rect 173222 314038 173306 314274
rect 173542 314038 192986 314274
rect 193222 314038 193306 314274
rect 193542 314038 572986 314274
rect 573222 314038 573306 314274
rect 573542 314038 591102 314274
rect 591338 314038 591422 314274
rect 591658 314038 592650 314274
rect -8726 313876 592650 314038
rect -2966 313294 586890 313456
rect -2966 313058 -2934 313294
rect -2698 313058 -2614 313294
rect -2378 313058 11826 313294
rect 12062 313058 12146 313294
rect 12382 313058 30328 313294
rect 30564 313058 166056 313294
rect 166292 313058 171826 313294
rect 172062 313058 172146 313294
rect 172382 313058 191826 313294
rect 192062 313058 192146 313294
rect 192382 313058 219610 313294
rect 219846 313058 250330 313294
rect 250566 313058 281050 313294
rect 281286 313058 311770 313294
rect 312006 313058 342490 313294
rect 342726 313058 373210 313294
rect 373446 313058 403930 313294
rect 404166 313058 434650 313294
rect 434886 313058 465370 313294
rect 465606 313058 496090 313294
rect 496326 313058 526810 313294
rect 527046 313058 571826 313294
rect 572062 313058 572146 313294
rect 572382 313058 586302 313294
rect 586538 313058 586622 313294
rect 586858 313058 586890 313294
rect -2966 312896 586890 313058
rect -6806 310614 590730 310776
rect -6806 310378 -5814 310614
rect -5578 310378 -5494 310614
rect -5258 310378 9266 310614
rect 9502 310378 9586 310614
rect 9822 310378 169266 310614
rect 169502 310378 169586 310614
rect 169822 310378 189266 310614
rect 189502 310378 189586 310614
rect 189822 310378 569266 310614
rect 569502 310378 569586 310614
rect 569822 310378 589182 310614
rect 589418 310378 589502 310614
rect 589738 310378 590730 310614
rect -6806 310216 590730 310378
rect -4886 306954 588810 307116
rect -4886 306718 -3894 306954
rect -3658 306718 -3574 306954
rect -3338 306718 5546 306954
rect 5782 306718 5866 306954
rect 6102 306718 25546 306954
rect 25782 306718 25866 306954
rect 26102 306718 185546 306954
rect 185782 306718 185866 306954
rect 186102 306718 565546 306954
rect 565782 306718 565866 306954
rect 566102 306718 587262 306954
rect 587498 306718 587582 306954
rect 587818 306718 588810 306954
rect -4886 306556 588810 306718
rect -8726 304274 592650 304436
rect -8726 304038 -8694 304274
rect -8458 304038 -8374 304274
rect -8138 304038 22986 304274
rect 23222 304038 23306 304274
rect 23542 304038 182986 304274
rect 183222 304038 183306 304274
rect 183542 304038 562986 304274
rect 563222 304038 563306 304274
rect 563542 304038 592062 304274
rect 592298 304038 592382 304274
rect 592618 304038 592650 304274
rect -8726 303876 592650 304038
rect -2966 303294 586890 303456
rect -2966 303058 -1974 303294
rect -1738 303058 -1654 303294
rect -1418 303058 1826 303294
rect 2062 303058 2146 303294
rect 2382 303058 21826 303294
rect 22062 303058 22146 303294
rect 22382 303058 31008 303294
rect 31244 303058 165376 303294
rect 165612 303058 181826 303294
rect 182062 303058 182146 303294
rect 182382 303058 204250 303294
rect 204486 303058 234970 303294
rect 235206 303058 265690 303294
rect 265926 303058 296410 303294
rect 296646 303058 327130 303294
rect 327366 303058 357850 303294
rect 358086 303058 388570 303294
rect 388806 303058 419290 303294
rect 419526 303058 450010 303294
rect 450246 303058 480730 303294
rect 480966 303058 511450 303294
rect 511686 303058 542170 303294
rect 542406 303058 561826 303294
rect 562062 303058 562146 303294
rect 562382 303058 581826 303294
rect 582062 303058 582146 303294
rect 582382 303058 585342 303294
rect 585578 303058 585662 303294
rect 585898 303058 586890 303294
rect -2966 302896 586890 303058
rect -6806 300614 590730 300776
rect -6806 300378 -6774 300614
rect -6538 300378 -6454 300614
rect -6218 300378 19266 300614
rect 19502 300378 19586 300614
rect 19822 300378 179266 300614
rect 179502 300378 179586 300614
rect 179822 300378 559266 300614
rect 559502 300378 559586 300614
rect 559822 300378 579266 300614
rect 579502 300378 579586 300614
rect 579822 300378 590142 300614
rect 590378 300378 590462 300614
rect 590698 300378 590730 300614
rect -6806 300216 590730 300378
rect -4886 296954 588810 297116
rect -4886 296718 -4854 296954
rect -4618 296718 -4534 296954
rect -4298 296718 15546 296954
rect 15782 296718 15866 296954
rect 16102 296718 175546 296954
rect 175782 296718 175866 296954
rect 176102 296718 195546 296954
rect 195782 296718 195866 296954
rect 196102 296718 575546 296954
rect 575782 296718 575866 296954
rect 576102 296718 588222 296954
rect 588458 296718 588542 296954
rect 588778 296718 588810 296954
rect -4886 296556 588810 296718
rect -8726 294274 592650 294436
rect -8726 294038 -7734 294274
rect -7498 294038 -7414 294274
rect -7178 294038 12986 294274
rect 13222 294038 13306 294274
rect 13542 294038 172986 294274
rect 173222 294038 173306 294274
rect 173542 294038 192986 294274
rect 193222 294038 193306 294274
rect 193542 294038 572986 294274
rect 573222 294038 573306 294274
rect 573542 294038 591102 294274
rect 591338 294038 591422 294274
rect 591658 294038 592650 294274
rect -8726 293876 592650 294038
rect -2966 293294 586890 293456
rect -2966 293058 -2934 293294
rect -2698 293058 -2614 293294
rect -2378 293058 11826 293294
rect 12062 293058 12146 293294
rect 12382 293058 30328 293294
rect 30564 293058 166056 293294
rect 166292 293058 171826 293294
rect 172062 293058 172146 293294
rect 172382 293058 191826 293294
rect 192062 293058 192146 293294
rect 192382 293058 219610 293294
rect 219846 293058 250330 293294
rect 250566 293058 281050 293294
rect 281286 293058 311770 293294
rect 312006 293058 342490 293294
rect 342726 293058 373210 293294
rect 373446 293058 403930 293294
rect 404166 293058 434650 293294
rect 434886 293058 465370 293294
rect 465606 293058 496090 293294
rect 496326 293058 526810 293294
rect 527046 293058 571826 293294
rect 572062 293058 572146 293294
rect 572382 293058 586302 293294
rect 586538 293058 586622 293294
rect 586858 293058 586890 293294
rect -2966 292896 586890 293058
rect -6806 290614 590730 290776
rect -6806 290378 -5814 290614
rect -5578 290378 -5494 290614
rect -5258 290378 9266 290614
rect 9502 290378 9586 290614
rect 9822 290378 169266 290614
rect 169502 290378 169586 290614
rect 169822 290378 189266 290614
rect 189502 290378 189586 290614
rect 189822 290378 569266 290614
rect 569502 290378 569586 290614
rect 569822 290378 589182 290614
rect 589418 290378 589502 290614
rect 589738 290378 590730 290614
rect -6806 290216 590730 290378
rect -4886 286954 588810 287116
rect -4886 286718 -3894 286954
rect -3658 286718 -3574 286954
rect -3338 286718 5546 286954
rect 5782 286718 5866 286954
rect 6102 286718 25546 286954
rect 25782 286718 25866 286954
rect 26102 286718 185546 286954
rect 185782 286718 185866 286954
rect 186102 286718 565546 286954
rect 565782 286718 565866 286954
rect 566102 286718 587262 286954
rect 587498 286718 587582 286954
rect 587818 286718 588810 286954
rect -4886 286556 588810 286718
rect -8726 284274 592650 284436
rect -8726 284038 -8694 284274
rect -8458 284038 -8374 284274
rect -8138 284038 22986 284274
rect 23222 284038 23306 284274
rect 23542 284038 182986 284274
rect 183222 284038 183306 284274
rect 183542 284038 562986 284274
rect 563222 284038 563306 284274
rect 563542 284038 592062 284274
rect 592298 284038 592382 284274
rect 592618 284038 592650 284274
rect -8726 283876 592650 284038
rect -2966 283294 586890 283456
rect -2966 283058 -1974 283294
rect -1738 283058 -1654 283294
rect -1418 283058 1826 283294
rect 2062 283058 2146 283294
rect 2382 283058 21826 283294
rect 22062 283058 22146 283294
rect 22382 283058 31008 283294
rect 31244 283058 165376 283294
rect 165612 283058 181826 283294
rect 182062 283058 182146 283294
rect 182382 283058 204250 283294
rect 204486 283058 234970 283294
rect 235206 283058 265690 283294
rect 265926 283058 296410 283294
rect 296646 283058 327130 283294
rect 327366 283058 357850 283294
rect 358086 283058 388570 283294
rect 388806 283058 419290 283294
rect 419526 283058 450010 283294
rect 450246 283058 480730 283294
rect 480966 283058 511450 283294
rect 511686 283058 542170 283294
rect 542406 283058 561826 283294
rect 562062 283058 562146 283294
rect 562382 283058 581826 283294
rect 582062 283058 582146 283294
rect 582382 283058 585342 283294
rect 585578 283058 585662 283294
rect 585898 283058 586890 283294
rect -2966 282896 586890 283058
rect -6806 280614 590730 280776
rect -6806 280378 -6774 280614
rect -6538 280378 -6454 280614
rect -6218 280378 19266 280614
rect 19502 280378 19586 280614
rect 19822 280378 179266 280614
rect 179502 280378 179586 280614
rect 179822 280378 559266 280614
rect 559502 280378 559586 280614
rect 559822 280378 579266 280614
rect 579502 280378 579586 280614
rect 579822 280378 590142 280614
rect 590378 280378 590462 280614
rect 590698 280378 590730 280614
rect -6806 280216 590730 280378
rect -4886 276954 588810 277116
rect -4886 276718 -4854 276954
rect -4618 276718 -4534 276954
rect -4298 276718 15546 276954
rect 15782 276718 15866 276954
rect 16102 276718 175546 276954
rect 175782 276718 175866 276954
rect 176102 276718 195546 276954
rect 195782 276718 195866 276954
rect 196102 276718 575546 276954
rect 575782 276718 575866 276954
rect 576102 276718 588222 276954
rect 588458 276718 588542 276954
rect 588778 276718 588810 276954
rect -4886 276556 588810 276718
rect -8726 274274 592650 274436
rect -8726 274038 -7734 274274
rect -7498 274038 -7414 274274
rect -7178 274038 12986 274274
rect 13222 274038 13306 274274
rect 13542 274038 172986 274274
rect 173222 274038 173306 274274
rect 173542 274038 192986 274274
rect 193222 274038 193306 274274
rect 193542 274038 572986 274274
rect 573222 274038 573306 274274
rect 573542 274038 591102 274274
rect 591338 274038 591422 274274
rect 591658 274038 592650 274274
rect -8726 273876 592650 274038
rect -2966 273294 586890 273456
rect -2966 273058 -2934 273294
rect -2698 273058 -2614 273294
rect -2378 273058 11826 273294
rect 12062 273058 12146 273294
rect 12382 273058 30328 273294
rect 30564 273058 166056 273294
rect 166292 273058 171826 273294
rect 172062 273058 172146 273294
rect 172382 273058 191826 273294
rect 192062 273058 192146 273294
rect 192382 273058 219610 273294
rect 219846 273058 250330 273294
rect 250566 273058 281050 273294
rect 281286 273058 311770 273294
rect 312006 273058 342490 273294
rect 342726 273058 373210 273294
rect 373446 273058 403930 273294
rect 404166 273058 434650 273294
rect 434886 273058 465370 273294
rect 465606 273058 496090 273294
rect 496326 273058 526810 273294
rect 527046 273058 571826 273294
rect 572062 273058 572146 273294
rect 572382 273058 586302 273294
rect 586538 273058 586622 273294
rect 586858 273058 586890 273294
rect -2966 272896 586890 273058
rect -6806 270614 590730 270776
rect -6806 270378 -5814 270614
rect -5578 270378 -5494 270614
rect -5258 270378 9266 270614
rect 9502 270378 9586 270614
rect 9822 270378 169266 270614
rect 169502 270378 169586 270614
rect 169822 270378 189266 270614
rect 189502 270378 189586 270614
rect 189822 270378 569266 270614
rect 569502 270378 569586 270614
rect 569822 270378 589182 270614
rect 589418 270378 589502 270614
rect 589738 270378 590730 270614
rect -6806 270216 590730 270378
rect -4886 266954 588810 267116
rect -4886 266718 -3894 266954
rect -3658 266718 -3574 266954
rect -3338 266718 5546 266954
rect 5782 266718 5866 266954
rect 6102 266718 25546 266954
rect 25782 266718 25866 266954
rect 26102 266718 185546 266954
rect 185782 266718 185866 266954
rect 186102 266718 565546 266954
rect 565782 266718 565866 266954
rect 566102 266718 587262 266954
rect 587498 266718 587582 266954
rect 587818 266718 588810 266954
rect -4886 266556 588810 266718
rect -8726 264274 592650 264436
rect -8726 264038 -8694 264274
rect -8458 264038 -8374 264274
rect -8138 264038 22986 264274
rect 23222 264038 23306 264274
rect 23542 264038 182986 264274
rect 183222 264038 183306 264274
rect 183542 264038 562986 264274
rect 563222 264038 563306 264274
rect 563542 264038 592062 264274
rect 592298 264038 592382 264274
rect 592618 264038 592650 264274
rect -8726 263876 592650 264038
rect -2966 263294 586890 263456
rect -2966 263058 -1974 263294
rect -1738 263058 -1654 263294
rect -1418 263058 1826 263294
rect 2062 263058 2146 263294
rect 2382 263058 21826 263294
rect 22062 263058 22146 263294
rect 22382 263058 31008 263294
rect 31244 263058 165376 263294
rect 165612 263058 181826 263294
rect 182062 263058 182146 263294
rect 182382 263058 204250 263294
rect 204486 263058 234970 263294
rect 235206 263058 265690 263294
rect 265926 263058 296410 263294
rect 296646 263058 327130 263294
rect 327366 263058 357850 263294
rect 358086 263058 388570 263294
rect 388806 263058 419290 263294
rect 419526 263058 450010 263294
rect 450246 263058 480730 263294
rect 480966 263058 511450 263294
rect 511686 263058 542170 263294
rect 542406 263058 561826 263294
rect 562062 263058 562146 263294
rect 562382 263058 581826 263294
rect 582062 263058 582146 263294
rect 582382 263058 585342 263294
rect 585578 263058 585662 263294
rect 585898 263058 586890 263294
rect -2966 262896 586890 263058
rect -6806 260614 590730 260776
rect -6806 260378 -6774 260614
rect -6538 260378 -6454 260614
rect -6218 260378 19266 260614
rect 19502 260378 19586 260614
rect 19822 260378 179266 260614
rect 179502 260378 179586 260614
rect 179822 260378 559266 260614
rect 559502 260378 559586 260614
rect 559822 260378 579266 260614
rect 579502 260378 579586 260614
rect 579822 260378 590142 260614
rect 590378 260378 590462 260614
rect 590698 260378 590730 260614
rect -6806 260216 590730 260378
rect -4886 256954 588810 257116
rect -4886 256718 -4854 256954
rect -4618 256718 -4534 256954
rect -4298 256718 15546 256954
rect 15782 256718 15866 256954
rect 16102 256718 175546 256954
rect 175782 256718 175866 256954
rect 176102 256718 195546 256954
rect 195782 256718 195866 256954
rect 196102 256718 575546 256954
rect 575782 256718 575866 256954
rect 576102 256718 588222 256954
rect 588458 256718 588542 256954
rect 588778 256718 588810 256954
rect -4886 256556 588810 256718
rect -8726 254274 592650 254436
rect -8726 254038 -7734 254274
rect -7498 254038 -7414 254274
rect -7178 254038 12986 254274
rect 13222 254038 13306 254274
rect 13542 254038 172986 254274
rect 173222 254038 173306 254274
rect 173542 254038 192986 254274
rect 193222 254038 193306 254274
rect 193542 254038 572986 254274
rect 573222 254038 573306 254274
rect 573542 254038 591102 254274
rect 591338 254038 591422 254274
rect 591658 254038 592650 254274
rect -8726 253876 592650 254038
rect -2966 253294 586890 253456
rect -2966 253058 -2934 253294
rect -2698 253058 -2614 253294
rect -2378 253058 11826 253294
rect 12062 253058 12146 253294
rect 12382 253058 171826 253294
rect 172062 253058 172146 253294
rect 172382 253058 191826 253294
rect 192062 253058 192146 253294
rect 192382 253058 219610 253294
rect 219846 253058 250330 253294
rect 250566 253058 281050 253294
rect 281286 253058 311770 253294
rect 312006 253058 342490 253294
rect 342726 253058 373210 253294
rect 373446 253058 403930 253294
rect 404166 253058 434650 253294
rect 434886 253058 465370 253294
rect 465606 253058 496090 253294
rect 496326 253058 526810 253294
rect 527046 253058 571826 253294
rect 572062 253058 572146 253294
rect 572382 253058 586302 253294
rect 586538 253058 586622 253294
rect 586858 253058 586890 253294
rect -2966 252896 586890 253058
rect -6806 250614 590730 250776
rect -6806 250378 -5814 250614
rect -5578 250378 -5494 250614
rect -5258 250378 9266 250614
rect 9502 250378 9586 250614
rect 9822 250378 29266 250614
rect 29502 250378 29586 250614
rect 29822 250378 49266 250614
rect 49502 250378 49586 250614
rect 49822 250378 69266 250614
rect 69502 250378 69586 250614
rect 69822 250378 89266 250614
rect 89502 250378 89586 250614
rect 89822 250378 109266 250614
rect 109502 250378 109586 250614
rect 109822 250378 129266 250614
rect 129502 250378 129586 250614
rect 129822 250378 149266 250614
rect 149502 250378 149586 250614
rect 149822 250378 169266 250614
rect 169502 250378 169586 250614
rect 169822 250378 189266 250614
rect 189502 250378 189586 250614
rect 189822 250378 569266 250614
rect 569502 250378 569586 250614
rect 569822 250378 589182 250614
rect 589418 250378 589502 250614
rect 589738 250378 590730 250614
rect -6806 250216 590730 250378
rect -4886 246954 588810 247116
rect -4886 246718 -3894 246954
rect -3658 246718 -3574 246954
rect -3338 246718 5546 246954
rect 5782 246718 5866 246954
rect 6102 246718 25546 246954
rect 25782 246718 25866 246954
rect 26102 246718 45546 246954
rect 45782 246718 45866 246954
rect 46102 246718 65546 246954
rect 65782 246718 65866 246954
rect 66102 246718 85546 246954
rect 85782 246718 85866 246954
rect 86102 246718 105546 246954
rect 105782 246718 105866 246954
rect 106102 246718 125546 246954
rect 125782 246718 125866 246954
rect 126102 246718 145546 246954
rect 145782 246718 145866 246954
rect 146102 246718 165546 246954
rect 165782 246718 165866 246954
rect 166102 246718 185546 246954
rect 185782 246718 185866 246954
rect 186102 246718 565546 246954
rect 565782 246718 565866 246954
rect 566102 246718 587262 246954
rect 587498 246718 587582 246954
rect 587818 246718 588810 246954
rect -4886 246556 588810 246718
rect -8726 244274 592650 244436
rect -8726 244038 -8694 244274
rect -8458 244038 -8374 244274
rect -8138 244038 22986 244274
rect 23222 244038 23306 244274
rect 23542 244038 42986 244274
rect 43222 244038 43306 244274
rect 43542 244038 62986 244274
rect 63222 244038 63306 244274
rect 63542 244038 82986 244274
rect 83222 244038 83306 244274
rect 83542 244038 102986 244274
rect 103222 244038 103306 244274
rect 103542 244038 122986 244274
rect 123222 244038 123306 244274
rect 123542 244038 142986 244274
rect 143222 244038 143306 244274
rect 143542 244038 162986 244274
rect 163222 244038 163306 244274
rect 163542 244038 182986 244274
rect 183222 244038 183306 244274
rect 183542 244038 562986 244274
rect 563222 244038 563306 244274
rect 563542 244038 592062 244274
rect 592298 244038 592382 244274
rect 592618 244038 592650 244274
rect -8726 243876 592650 244038
rect -2966 243294 586890 243456
rect -2966 243058 -1974 243294
rect -1738 243058 -1654 243294
rect -1418 243058 1826 243294
rect 2062 243058 2146 243294
rect 2382 243058 21826 243294
rect 22062 243058 22146 243294
rect 22382 243058 41826 243294
rect 42062 243058 42146 243294
rect 42382 243058 61826 243294
rect 62062 243058 62146 243294
rect 62382 243058 81826 243294
rect 82062 243058 82146 243294
rect 82382 243058 101826 243294
rect 102062 243058 102146 243294
rect 102382 243058 121826 243294
rect 122062 243058 122146 243294
rect 122382 243058 141826 243294
rect 142062 243058 142146 243294
rect 142382 243058 161826 243294
rect 162062 243058 162146 243294
rect 162382 243058 181826 243294
rect 182062 243058 182146 243294
rect 182382 243058 204250 243294
rect 204486 243058 234970 243294
rect 235206 243058 265690 243294
rect 265926 243058 296410 243294
rect 296646 243058 327130 243294
rect 327366 243058 357850 243294
rect 358086 243058 388570 243294
rect 388806 243058 419290 243294
rect 419526 243058 450010 243294
rect 450246 243058 480730 243294
rect 480966 243058 511450 243294
rect 511686 243058 542170 243294
rect 542406 243058 561826 243294
rect 562062 243058 562146 243294
rect 562382 243058 581826 243294
rect 582062 243058 582146 243294
rect 582382 243058 585342 243294
rect 585578 243058 585662 243294
rect 585898 243058 586890 243294
rect -2966 242896 586890 243058
rect -6806 240614 590730 240776
rect -6806 240378 -6774 240614
rect -6538 240378 -6454 240614
rect -6218 240378 19266 240614
rect 19502 240378 19586 240614
rect 19822 240378 39266 240614
rect 39502 240378 39586 240614
rect 39822 240378 59266 240614
rect 59502 240378 59586 240614
rect 59822 240378 79266 240614
rect 79502 240378 79586 240614
rect 79822 240378 99266 240614
rect 99502 240378 99586 240614
rect 99822 240378 119266 240614
rect 119502 240378 119586 240614
rect 119822 240378 139266 240614
rect 139502 240378 139586 240614
rect 139822 240378 159266 240614
rect 159502 240378 159586 240614
rect 159822 240378 179266 240614
rect 179502 240378 179586 240614
rect 179822 240378 559266 240614
rect 559502 240378 559586 240614
rect 559822 240378 579266 240614
rect 579502 240378 579586 240614
rect 579822 240378 590142 240614
rect 590378 240378 590462 240614
rect 590698 240378 590730 240614
rect -6806 240216 590730 240378
rect -4886 236954 588810 237116
rect -4886 236718 -4854 236954
rect -4618 236718 -4534 236954
rect -4298 236718 15546 236954
rect 15782 236718 15866 236954
rect 16102 236718 35546 236954
rect 35782 236718 35866 236954
rect 36102 236718 55546 236954
rect 55782 236718 55866 236954
rect 56102 236718 75546 236954
rect 75782 236718 75866 236954
rect 76102 236718 95546 236954
rect 95782 236718 95866 236954
rect 96102 236718 115546 236954
rect 115782 236718 115866 236954
rect 116102 236718 135546 236954
rect 135782 236718 135866 236954
rect 136102 236718 155546 236954
rect 155782 236718 155866 236954
rect 156102 236718 175546 236954
rect 175782 236718 175866 236954
rect 176102 236718 195546 236954
rect 195782 236718 195866 236954
rect 196102 236718 575546 236954
rect 575782 236718 575866 236954
rect 576102 236718 588222 236954
rect 588458 236718 588542 236954
rect 588778 236718 588810 236954
rect -4886 236556 588810 236718
rect -8726 234274 592650 234436
rect -8726 234038 -7734 234274
rect -7498 234038 -7414 234274
rect -7178 234038 12986 234274
rect 13222 234038 13306 234274
rect 13542 234038 32986 234274
rect 33222 234038 33306 234274
rect 33542 234038 52986 234274
rect 53222 234038 53306 234274
rect 53542 234038 72986 234274
rect 73222 234038 73306 234274
rect 73542 234038 92986 234274
rect 93222 234038 93306 234274
rect 93542 234038 112986 234274
rect 113222 234038 113306 234274
rect 113542 234038 132986 234274
rect 133222 234038 133306 234274
rect 133542 234038 152986 234274
rect 153222 234038 153306 234274
rect 153542 234038 172986 234274
rect 173222 234038 173306 234274
rect 173542 234038 192986 234274
rect 193222 234038 193306 234274
rect 193542 234038 572986 234274
rect 573222 234038 573306 234274
rect 573542 234038 591102 234274
rect 591338 234038 591422 234274
rect 591658 234038 592650 234274
rect -8726 233876 592650 234038
rect -2966 233294 586890 233456
rect -2966 233058 -2934 233294
rect -2698 233058 -2614 233294
rect -2378 233058 11826 233294
rect 12062 233058 12146 233294
rect 12382 233058 31826 233294
rect 32062 233058 32146 233294
rect 32382 233058 51826 233294
rect 52062 233058 52146 233294
rect 52382 233058 71826 233294
rect 72062 233058 72146 233294
rect 72382 233058 91826 233294
rect 92062 233058 92146 233294
rect 92382 233058 111826 233294
rect 112062 233058 112146 233294
rect 112382 233058 131826 233294
rect 132062 233058 132146 233294
rect 132382 233058 151826 233294
rect 152062 233058 152146 233294
rect 152382 233058 171826 233294
rect 172062 233058 172146 233294
rect 172382 233058 191826 233294
rect 192062 233058 192146 233294
rect 192382 233058 219610 233294
rect 219846 233058 250330 233294
rect 250566 233058 281050 233294
rect 281286 233058 311770 233294
rect 312006 233058 342490 233294
rect 342726 233058 373210 233294
rect 373446 233058 403930 233294
rect 404166 233058 434650 233294
rect 434886 233058 465370 233294
rect 465606 233058 496090 233294
rect 496326 233058 526810 233294
rect 527046 233058 571826 233294
rect 572062 233058 572146 233294
rect 572382 233058 586302 233294
rect 586538 233058 586622 233294
rect 586858 233058 586890 233294
rect -2966 232896 586890 233058
rect -6806 230614 590730 230776
rect -6806 230378 -5814 230614
rect -5578 230378 -5494 230614
rect -5258 230378 9266 230614
rect 9502 230378 9586 230614
rect 9822 230378 29266 230614
rect 29502 230378 29586 230614
rect 29822 230378 49266 230614
rect 49502 230378 49586 230614
rect 49822 230378 69266 230614
rect 69502 230378 69586 230614
rect 69822 230378 89266 230614
rect 89502 230378 89586 230614
rect 89822 230378 109266 230614
rect 109502 230378 109586 230614
rect 109822 230378 129266 230614
rect 129502 230378 129586 230614
rect 129822 230378 149266 230614
rect 149502 230378 149586 230614
rect 149822 230378 169266 230614
rect 169502 230378 169586 230614
rect 169822 230378 189266 230614
rect 189502 230378 189586 230614
rect 189822 230378 569266 230614
rect 569502 230378 569586 230614
rect 569822 230378 589182 230614
rect 589418 230378 589502 230614
rect 589738 230378 590730 230614
rect -6806 230216 590730 230378
rect -4886 226954 588810 227116
rect -4886 226718 -3894 226954
rect -3658 226718 -3574 226954
rect -3338 226718 5546 226954
rect 5782 226718 5866 226954
rect 6102 226718 25546 226954
rect 25782 226718 25866 226954
rect 26102 226718 185546 226954
rect 185782 226718 185866 226954
rect 186102 226718 565546 226954
rect 565782 226718 565866 226954
rect 566102 226718 587262 226954
rect 587498 226718 587582 226954
rect 587818 226718 588810 226954
rect -4886 226556 588810 226718
rect -8726 224274 592650 224436
rect -8726 224038 -8694 224274
rect -8458 224038 -8374 224274
rect -8138 224038 22986 224274
rect 23222 224038 23306 224274
rect 23542 224038 182986 224274
rect 183222 224038 183306 224274
rect 183542 224038 562986 224274
rect 563222 224038 563306 224274
rect 563542 224038 592062 224274
rect 592298 224038 592382 224274
rect 592618 224038 592650 224274
rect -8726 223876 592650 224038
rect -2966 223294 586890 223456
rect -2966 223058 -1974 223294
rect -1738 223058 -1654 223294
rect -1418 223058 1826 223294
rect 2062 223058 2146 223294
rect 2382 223058 21826 223294
rect 22062 223058 22146 223294
rect 22382 223058 31008 223294
rect 31244 223058 165376 223294
rect 165612 223058 181826 223294
rect 182062 223058 182146 223294
rect 182382 223058 204250 223294
rect 204486 223058 234970 223294
rect 235206 223058 265690 223294
rect 265926 223058 296410 223294
rect 296646 223058 327130 223294
rect 327366 223058 357850 223294
rect 358086 223058 388570 223294
rect 388806 223058 419290 223294
rect 419526 223058 450010 223294
rect 450246 223058 480730 223294
rect 480966 223058 511450 223294
rect 511686 223058 542170 223294
rect 542406 223058 561826 223294
rect 562062 223058 562146 223294
rect 562382 223058 581826 223294
rect 582062 223058 582146 223294
rect 582382 223058 585342 223294
rect 585578 223058 585662 223294
rect 585898 223058 586890 223294
rect -2966 222896 586890 223058
rect -6806 220614 590730 220776
rect -6806 220378 -6774 220614
rect -6538 220378 -6454 220614
rect -6218 220378 19266 220614
rect 19502 220378 19586 220614
rect 19822 220378 179266 220614
rect 179502 220378 179586 220614
rect 179822 220378 559266 220614
rect 559502 220378 559586 220614
rect 559822 220378 579266 220614
rect 579502 220378 579586 220614
rect 579822 220378 590142 220614
rect 590378 220378 590462 220614
rect 590698 220378 590730 220614
rect -6806 220216 590730 220378
rect -4886 216954 588810 217116
rect -4886 216718 -4854 216954
rect -4618 216718 -4534 216954
rect -4298 216718 15546 216954
rect 15782 216718 15866 216954
rect 16102 216718 175546 216954
rect 175782 216718 175866 216954
rect 176102 216718 195546 216954
rect 195782 216718 195866 216954
rect 196102 216718 575546 216954
rect 575782 216718 575866 216954
rect 576102 216718 588222 216954
rect 588458 216718 588542 216954
rect 588778 216718 588810 216954
rect -4886 216556 588810 216718
rect -8726 214274 592650 214436
rect -8726 214038 -7734 214274
rect -7498 214038 -7414 214274
rect -7178 214038 12986 214274
rect 13222 214038 13306 214274
rect 13542 214038 172986 214274
rect 173222 214038 173306 214274
rect 173542 214038 192986 214274
rect 193222 214038 193306 214274
rect 193542 214038 572986 214274
rect 573222 214038 573306 214274
rect 573542 214038 591102 214274
rect 591338 214038 591422 214274
rect 591658 214038 592650 214274
rect -8726 213876 592650 214038
rect -2966 213294 586890 213456
rect -2966 213058 -2934 213294
rect -2698 213058 -2614 213294
rect -2378 213058 11826 213294
rect 12062 213058 12146 213294
rect 12382 213058 30328 213294
rect 30564 213058 166056 213294
rect 166292 213058 171826 213294
rect 172062 213058 172146 213294
rect 172382 213058 191826 213294
rect 192062 213058 192146 213294
rect 192382 213058 219610 213294
rect 219846 213058 250330 213294
rect 250566 213058 281050 213294
rect 281286 213058 311770 213294
rect 312006 213058 342490 213294
rect 342726 213058 373210 213294
rect 373446 213058 403930 213294
rect 404166 213058 434650 213294
rect 434886 213058 465370 213294
rect 465606 213058 496090 213294
rect 496326 213058 526810 213294
rect 527046 213058 571826 213294
rect 572062 213058 572146 213294
rect 572382 213058 586302 213294
rect 586538 213058 586622 213294
rect 586858 213058 586890 213294
rect -2966 212896 586890 213058
rect -6806 210614 590730 210776
rect -6806 210378 -5814 210614
rect -5578 210378 -5494 210614
rect -5258 210378 9266 210614
rect 9502 210378 9586 210614
rect 9822 210378 169266 210614
rect 169502 210378 169586 210614
rect 169822 210378 189266 210614
rect 189502 210378 189586 210614
rect 189822 210378 569266 210614
rect 569502 210378 569586 210614
rect 569822 210378 589182 210614
rect 589418 210378 589502 210614
rect 589738 210378 590730 210614
rect -6806 210216 590730 210378
rect -4886 206954 588810 207116
rect -4886 206718 -3894 206954
rect -3658 206718 -3574 206954
rect -3338 206718 5546 206954
rect 5782 206718 5866 206954
rect 6102 206718 25546 206954
rect 25782 206718 25866 206954
rect 26102 206718 185546 206954
rect 185782 206718 185866 206954
rect 186102 206718 565546 206954
rect 565782 206718 565866 206954
rect 566102 206718 587262 206954
rect 587498 206718 587582 206954
rect 587818 206718 588810 206954
rect -4886 206556 588810 206718
rect -8726 204274 592650 204436
rect -8726 204038 -8694 204274
rect -8458 204038 -8374 204274
rect -8138 204038 22986 204274
rect 23222 204038 23306 204274
rect 23542 204038 182986 204274
rect 183222 204038 183306 204274
rect 183542 204038 562986 204274
rect 563222 204038 563306 204274
rect 563542 204038 592062 204274
rect 592298 204038 592382 204274
rect 592618 204038 592650 204274
rect -8726 203876 592650 204038
rect -2966 203294 586890 203456
rect -2966 203058 -1974 203294
rect -1738 203058 -1654 203294
rect -1418 203058 1826 203294
rect 2062 203058 2146 203294
rect 2382 203058 21826 203294
rect 22062 203058 22146 203294
rect 22382 203058 31008 203294
rect 31244 203058 165376 203294
rect 165612 203058 181826 203294
rect 182062 203058 182146 203294
rect 182382 203058 204250 203294
rect 204486 203058 234970 203294
rect 235206 203058 265690 203294
rect 265926 203058 296410 203294
rect 296646 203058 327130 203294
rect 327366 203058 357850 203294
rect 358086 203058 388570 203294
rect 388806 203058 419290 203294
rect 419526 203058 450010 203294
rect 450246 203058 480730 203294
rect 480966 203058 511450 203294
rect 511686 203058 542170 203294
rect 542406 203058 561826 203294
rect 562062 203058 562146 203294
rect 562382 203058 581826 203294
rect 582062 203058 582146 203294
rect 582382 203058 585342 203294
rect 585578 203058 585662 203294
rect 585898 203058 586890 203294
rect -2966 202896 586890 203058
rect -6806 200614 590730 200776
rect -6806 200378 -6774 200614
rect -6538 200378 -6454 200614
rect -6218 200378 19266 200614
rect 19502 200378 19586 200614
rect 19822 200378 179266 200614
rect 179502 200378 179586 200614
rect 179822 200378 559266 200614
rect 559502 200378 559586 200614
rect 559822 200378 579266 200614
rect 579502 200378 579586 200614
rect 579822 200378 590142 200614
rect 590378 200378 590462 200614
rect 590698 200378 590730 200614
rect -6806 200216 590730 200378
rect -4886 196954 588810 197116
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15546 196954
rect 15782 196718 15866 196954
rect 16102 196718 175546 196954
rect 175782 196718 175866 196954
rect 176102 196718 195546 196954
rect 195782 196718 195866 196954
rect 196102 196718 575546 196954
rect 575782 196718 575866 196954
rect 576102 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect -4886 196556 588810 196718
rect -8726 194274 592650 194436
rect -8726 194038 -7734 194274
rect -7498 194038 -7414 194274
rect -7178 194038 12986 194274
rect 13222 194038 13306 194274
rect 13542 194038 172986 194274
rect 173222 194038 173306 194274
rect 173542 194038 192986 194274
rect 193222 194038 193306 194274
rect 193542 194038 572986 194274
rect 573222 194038 573306 194274
rect 573542 194038 591102 194274
rect 591338 194038 591422 194274
rect 591658 194038 592650 194274
rect -8726 193876 592650 194038
rect -2966 193294 586890 193456
rect -2966 193058 -2934 193294
rect -2698 193058 -2614 193294
rect -2378 193058 11826 193294
rect 12062 193058 12146 193294
rect 12382 193058 30328 193294
rect 30564 193058 166056 193294
rect 166292 193058 171826 193294
rect 172062 193058 172146 193294
rect 172382 193058 191826 193294
rect 192062 193058 192146 193294
rect 192382 193058 219610 193294
rect 219846 193058 250330 193294
rect 250566 193058 281050 193294
rect 281286 193058 311770 193294
rect 312006 193058 342490 193294
rect 342726 193058 373210 193294
rect 373446 193058 403930 193294
rect 404166 193058 434650 193294
rect 434886 193058 465370 193294
rect 465606 193058 496090 193294
rect 496326 193058 526810 193294
rect 527046 193058 571826 193294
rect 572062 193058 572146 193294
rect 572382 193058 586302 193294
rect 586538 193058 586622 193294
rect 586858 193058 586890 193294
rect -2966 192896 586890 193058
rect -6806 190614 590730 190776
rect -6806 190378 -5814 190614
rect -5578 190378 -5494 190614
rect -5258 190378 9266 190614
rect 9502 190378 9586 190614
rect 9822 190378 169266 190614
rect 169502 190378 169586 190614
rect 169822 190378 189266 190614
rect 189502 190378 189586 190614
rect 189822 190378 569266 190614
rect 569502 190378 569586 190614
rect 569822 190378 589182 190614
rect 589418 190378 589502 190614
rect 589738 190378 590730 190614
rect -6806 190216 590730 190378
rect -4886 186954 588810 187116
rect -4886 186718 -3894 186954
rect -3658 186718 -3574 186954
rect -3338 186718 5546 186954
rect 5782 186718 5866 186954
rect 6102 186718 25546 186954
rect 25782 186718 25866 186954
rect 26102 186718 185546 186954
rect 185782 186718 185866 186954
rect 186102 186718 565546 186954
rect 565782 186718 565866 186954
rect 566102 186718 587262 186954
rect 587498 186718 587582 186954
rect 587818 186718 588810 186954
rect -4886 186556 588810 186718
rect -8726 184274 592650 184436
rect -8726 184038 -8694 184274
rect -8458 184038 -8374 184274
rect -8138 184038 22986 184274
rect 23222 184038 23306 184274
rect 23542 184038 182986 184274
rect 183222 184038 183306 184274
rect 183542 184038 562986 184274
rect 563222 184038 563306 184274
rect 563542 184038 592062 184274
rect 592298 184038 592382 184274
rect 592618 184038 592650 184274
rect -8726 183876 592650 184038
rect -2966 183294 586890 183456
rect -2966 183058 -1974 183294
rect -1738 183058 -1654 183294
rect -1418 183058 1826 183294
rect 2062 183058 2146 183294
rect 2382 183058 21826 183294
rect 22062 183058 22146 183294
rect 22382 183058 31008 183294
rect 31244 183058 165376 183294
rect 165612 183058 181826 183294
rect 182062 183058 182146 183294
rect 182382 183058 204250 183294
rect 204486 183058 234970 183294
rect 235206 183058 265690 183294
rect 265926 183058 296410 183294
rect 296646 183058 327130 183294
rect 327366 183058 357850 183294
rect 358086 183058 388570 183294
rect 388806 183058 419290 183294
rect 419526 183058 450010 183294
rect 450246 183058 480730 183294
rect 480966 183058 511450 183294
rect 511686 183058 542170 183294
rect 542406 183058 561826 183294
rect 562062 183058 562146 183294
rect 562382 183058 581826 183294
rect 582062 183058 582146 183294
rect 582382 183058 585342 183294
rect 585578 183058 585662 183294
rect 585898 183058 586890 183294
rect -2966 182896 586890 183058
rect -6806 180614 590730 180776
rect -6806 180378 -6774 180614
rect -6538 180378 -6454 180614
rect -6218 180378 19266 180614
rect 19502 180378 19586 180614
rect 19822 180378 179266 180614
rect 179502 180378 179586 180614
rect 179822 180378 559266 180614
rect 559502 180378 559586 180614
rect 559822 180378 579266 180614
rect 579502 180378 579586 180614
rect 579822 180378 590142 180614
rect 590378 180378 590462 180614
rect 590698 180378 590730 180614
rect -6806 180216 590730 180378
rect -4886 176954 588810 177116
rect -4886 176718 -4854 176954
rect -4618 176718 -4534 176954
rect -4298 176718 15546 176954
rect 15782 176718 15866 176954
rect 16102 176718 175546 176954
rect 175782 176718 175866 176954
rect 176102 176718 195546 176954
rect 195782 176718 195866 176954
rect 196102 176718 575546 176954
rect 575782 176718 575866 176954
rect 576102 176718 588222 176954
rect 588458 176718 588542 176954
rect 588778 176718 588810 176954
rect -4886 176556 588810 176718
rect -8726 174274 592650 174436
rect -8726 174038 -7734 174274
rect -7498 174038 -7414 174274
rect -7178 174038 12986 174274
rect 13222 174038 13306 174274
rect 13542 174038 172986 174274
rect 173222 174038 173306 174274
rect 173542 174038 192986 174274
rect 193222 174038 193306 174274
rect 193542 174038 572986 174274
rect 573222 174038 573306 174274
rect 573542 174038 591102 174274
rect 591338 174038 591422 174274
rect 591658 174038 592650 174274
rect -8726 173876 592650 174038
rect -2966 173294 586890 173456
rect -2966 173058 -2934 173294
rect -2698 173058 -2614 173294
rect -2378 173058 11826 173294
rect 12062 173058 12146 173294
rect 12382 173058 30328 173294
rect 30564 173058 166056 173294
rect 166292 173058 171826 173294
rect 172062 173058 172146 173294
rect 172382 173058 191826 173294
rect 192062 173058 192146 173294
rect 192382 173058 219610 173294
rect 219846 173058 250330 173294
rect 250566 173058 281050 173294
rect 281286 173058 311770 173294
rect 312006 173058 342490 173294
rect 342726 173058 373210 173294
rect 373446 173058 403930 173294
rect 404166 173058 434650 173294
rect 434886 173058 465370 173294
rect 465606 173058 496090 173294
rect 496326 173058 526810 173294
rect 527046 173058 571826 173294
rect 572062 173058 572146 173294
rect 572382 173058 586302 173294
rect 586538 173058 586622 173294
rect 586858 173058 586890 173294
rect -2966 172896 586890 173058
rect -6806 170614 590730 170776
rect -6806 170378 -5814 170614
rect -5578 170378 -5494 170614
rect -5258 170378 9266 170614
rect 9502 170378 9586 170614
rect 9822 170378 169266 170614
rect 169502 170378 169586 170614
rect 169822 170378 189266 170614
rect 189502 170378 189586 170614
rect 189822 170378 569266 170614
rect 569502 170378 569586 170614
rect 569822 170378 589182 170614
rect 589418 170378 589502 170614
rect 589738 170378 590730 170614
rect -6806 170216 590730 170378
rect -4886 166954 588810 167116
rect -4886 166718 -3894 166954
rect -3658 166718 -3574 166954
rect -3338 166718 5546 166954
rect 5782 166718 5866 166954
rect 6102 166718 25546 166954
rect 25782 166718 25866 166954
rect 26102 166718 185546 166954
rect 185782 166718 185866 166954
rect 186102 166718 565546 166954
rect 565782 166718 565866 166954
rect 566102 166718 587262 166954
rect 587498 166718 587582 166954
rect 587818 166718 588810 166954
rect -4886 166556 588810 166718
rect -8726 164274 592650 164436
rect -8726 164038 -8694 164274
rect -8458 164038 -8374 164274
rect -8138 164038 22986 164274
rect 23222 164038 23306 164274
rect 23542 164038 182986 164274
rect 183222 164038 183306 164274
rect 183542 164038 562986 164274
rect 563222 164038 563306 164274
rect 563542 164038 592062 164274
rect 592298 164038 592382 164274
rect 592618 164038 592650 164274
rect -8726 163876 592650 164038
rect -2966 163294 586890 163456
rect -2966 163058 -1974 163294
rect -1738 163058 -1654 163294
rect -1418 163058 1826 163294
rect 2062 163058 2146 163294
rect 2382 163058 21826 163294
rect 22062 163058 22146 163294
rect 22382 163058 31008 163294
rect 31244 163058 165376 163294
rect 165612 163058 181826 163294
rect 182062 163058 182146 163294
rect 182382 163058 204250 163294
rect 204486 163058 234970 163294
rect 235206 163058 265690 163294
rect 265926 163058 296410 163294
rect 296646 163058 327130 163294
rect 327366 163058 357850 163294
rect 358086 163058 388570 163294
rect 388806 163058 419290 163294
rect 419526 163058 450010 163294
rect 450246 163058 480730 163294
rect 480966 163058 511450 163294
rect 511686 163058 542170 163294
rect 542406 163058 561826 163294
rect 562062 163058 562146 163294
rect 562382 163058 581826 163294
rect 582062 163058 582146 163294
rect 582382 163058 585342 163294
rect 585578 163058 585662 163294
rect 585898 163058 586890 163294
rect -2966 162896 586890 163058
rect -6806 160614 590730 160776
rect -6806 160378 -6774 160614
rect -6538 160378 -6454 160614
rect -6218 160378 19266 160614
rect 19502 160378 19586 160614
rect 19822 160378 179266 160614
rect 179502 160378 179586 160614
rect 179822 160378 559266 160614
rect 559502 160378 559586 160614
rect 559822 160378 579266 160614
rect 579502 160378 579586 160614
rect 579822 160378 590142 160614
rect 590378 160378 590462 160614
rect 590698 160378 590730 160614
rect -6806 160216 590730 160378
rect -4886 156954 588810 157116
rect -4886 156718 -4854 156954
rect -4618 156718 -4534 156954
rect -4298 156718 15546 156954
rect 15782 156718 15866 156954
rect 16102 156718 175546 156954
rect 175782 156718 175866 156954
rect 176102 156718 195546 156954
rect 195782 156718 195866 156954
rect 196102 156718 575546 156954
rect 575782 156718 575866 156954
rect 576102 156718 588222 156954
rect 588458 156718 588542 156954
rect 588778 156718 588810 156954
rect -4886 156556 588810 156718
rect -8726 154274 592650 154436
rect -8726 154038 -7734 154274
rect -7498 154038 -7414 154274
rect -7178 154038 12986 154274
rect 13222 154038 13306 154274
rect 13542 154038 172986 154274
rect 173222 154038 173306 154274
rect 173542 154038 192986 154274
rect 193222 154038 193306 154274
rect 193542 154038 572986 154274
rect 573222 154038 573306 154274
rect 573542 154038 591102 154274
rect 591338 154038 591422 154274
rect 591658 154038 592650 154274
rect -8726 153876 592650 154038
rect -2966 153294 586890 153456
rect -2966 153058 -2934 153294
rect -2698 153058 -2614 153294
rect -2378 153058 11826 153294
rect 12062 153058 12146 153294
rect 12382 153058 30328 153294
rect 30564 153058 166056 153294
rect 166292 153058 171826 153294
rect 172062 153058 172146 153294
rect 172382 153058 191826 153294
rect 192062 153058 192146 153294
rect 192382 153058 219610 153294
rect 219846 153058 250330 153294
rect 250566 153058 281050 153294
rect 281286 153058 311770 153294
rect 312006 153058 342490 153294
rect 342726 153058 373210 153294
rect 373446 153058 403930 153294
rect 404166 153058 434650 153294
rect 434886 153058 465370 153294
rect 465606 153058 496090 153294
rect 496326 153058 526810 153294
rect 527046 153058 571826 153294
rect 572062 153058 572146 153294
rect 572382 153058 586302 153294
rect 586538 153058 586622 153294
rect 586858 153058 586890 153294
rect -2966 152896 586890 153058
rect -6806 150614 590730 150776
rect -6806 150378 -5814 150614
rect -5578 150378 -5494 150614
rect -5258 150378 9266 150614
rect 9502 150378 9586 150614
rect 9822 150378 169266 150614
rect 169502 150378 169586 150614
rect 169822 150378 189266 150614
rect 189502 150378 189586 150614
rect 189822 150378 569266 150614
rect 569502 150378 569586 150614
rect 569822 150378 589182 150614
rect 589418 150378 589502 150614
rect 589738 150378 590730 150614
rect -6806 150216 590730 150378
rect -4886 146954 588810 147116
rect -4886 146718 -3894 146954
rect -3658 146718 -3574 146954
rect -3338 146718 5546 146954
rect 5782 146718 5866 146954
rect 6102 146718 25546 146954
rect 25782 146718 25866 146954
rect 26102 146718 185546 146954
rect 185782 146718 185866 146954
rect 186102 146718 565546 146954
rect 565782 146718 565866 146954
rect 566102 146718 587262 146954
rect 587498 146718 587582 146954
rect 587818 146718 588810 146954
rect -4886 146556 588810 146718
rect -8726 144274 592650 144436
rect -8726 144038 -8694 144274
rect -8458 144038 -8374 144274
rect -8138 144038 22986 144274
rect 23222 144038 23306 144274
rect 23542 144038 182986 144274
rect 183222 144038 183306 144274
rect 183542 144038 562986 144274
rect 563222 144038 563306 144274
rect 563542 144038 592062 144274
rect 592298 144038 592382 144274
rect 592618 144038 592650 144274
rect -8726 143876 592650 144038
rect -2966 143294 586890 143456
rect -2966 143058 -1974 143294
rect -1738 143058 -1654 143294
rect -1418 143058 1826 143294
rect 2062 143058 2146 143294
rect 2382 143058 21826 143294
rect 22062 143058 22146 143294
rect 22382 143058 181826 143294
rect 182062 143058 182146 143294
rect 182382 143058 204250 143294
rect 204486 143058 234970 143294
rect 235206 143058 265690 143294
rect 265926 143058 296410 143294
rect 296646 143058 327130 143294
rect 327366 143058 357850 143294
rect 358086 143058 388570 143294
rect 388806 143058 419290 143294
rect 419526 143058 450010 143294
rect 450246 143058 480730 143294
rect 480966 143058 511450 143294
rect 511686 143058 542170 143294
rect 542406 143058 561826 143294
rect 562062 143058 562146 143294
rect 562382 143058 581826 143294
rect 582062 143058 582146 143294
rect 582382 143058 585342 143294
rect 585578 143058 585662 143294
rect 585898 143058 586890 143294
rect -2966 142896 586890 143058
rect -6806 140614 590730 140776
rect -6806 140378 -6774 140614
rect -6538 140378 -6454 140614
rect -6218 140378 19266 140614
rect 19502 140378 19586 140614
rect 19822 140378 179266 140614
rect 179502 140378 179586 140614
rect 179822 140378 559266 140614
rect 559502 140378 559586 140614
rect 559822 140378 579266 140614
rect 579502 140378 579586 140614
rect 579822 140378 590142 140614
rect 590378 140378 590462 140614
rect 590698 140378 590730 140614
rect -6806 140216 590730 140378
rect -4886 136954 588810 137116
rect -4886 136718 -4854 136954
rect -4618 136718 -4534 136954
rect -4298 136718 15546 136954
rect 15782 136718 15866 136954
rect 16102 136718 35546 136954
rect 35782 136718 35866 136954
rect 36102 136718 55546 136954
rect 55782 136718 55866 136954
rect 56102 136718 75546 136954
rect 75782 136718 75866 136954
rect 76102 136718 95546 136954
rect 95782 136718 95866 136954
rect 96102 136718 115546 136954
rect 115782 136718 115866 136954
rect 116102 136718 135546 136954
rect 135782 136718 135866 136954
rect 136102 136718 155546 136954
rect 155782 136718 155866 136954
rect 156102 136718 175546 136954
rect 175782 136718 175866 136954
rect 176102 136718 195546 136954
rect 195782 136718 195866 136954
rect 196102 136718 575546 136954
rect 575782 136718 575866 136954
rect 576102 136718 588222 136954
rect 588458 136718 588542 136954
rect 588778 136718 588810 136954
rect -4886 136556 588810 136718
rect -8726 134274 592650 134436
rect -8726 134038 -7734 134274
rect -7498 134038 -7414 134274
rect -7178 134038 12986 134274
rect 13222 134038 13306 134274
rect 13542 134038 32986 134274
rect 33222 134038 33306 134274
rect 33542 134038 52986 134274
rect 53222 134038 53306 134274
rect 53542 134038 72986 134274
rect 73222 134038 73306 134274
rect 73542 134038 92986 134274
rect 93222 134038 93306 134274
rect 93542 134038 112986 134274
rect 113222 134038 113306 134274
rect 113542 134038 132986 134274
rect 133222 134038 133306 134274
rect 133542 134038 152986 134274
rect 153222 134038 153306 134274
rect 153542 134038 172986 134274
rect 173222 134038 173306 134274
rect 173542 134038 192986 134274
rect 193222 134038 193306 134274
rect 193542 134038 572986 134274
rect 573222 134038 573306 134274
rect 573542 134038 591102 134274
rect 591338 134038 591422 134274
rect 591658 134038 592650 134274
rect -8726 133876 592650 134038
rect -2966 133294 586890 133456
rect -2966 133058 -2934 133294
rect -2698 133058 -2614 133294
rect -2378 133058 11826 133294
rect 12062 133058 12146 133294
rect 12382 133058 31826 133294
rect 32062 133058 32146 133294
rect 32382 133058 51826 133294
rect 52062 133058 52146 133294
rect 52382 133058 71826 133294
rect 72062 133058 72146 133294
rect 72382 133058 91826 133294
rect 92062 133058 92146 133294
rect 92382 133058 111826 133294
rect 112062 133058 112146 133294
rect 112382 133058 131826 133294
rect 132062 133058 132146 133294
rect 132382 133058 151826 133294
rect 152062 133058 152146 133294
rect 152382 133058 171826 133294
rect 172062 133058 172146 133294
rect 172382 133058 191826 133294
rect 192062 133058 192146 133294
rect 192382 133058 219610 133294
rect 219846 133058 250330 133294
rect 250566 133058 281050 133294
rect 281286 133058 311770 133294
rect 312006 133058 342490 133294
rect 342726 133058 373210 133294
rect 373446 133058 403930 133294
rect 404166 133058 434650 133294
rect 434886 133058 465370 133294
rect 465606 133058 496090 133294
rect 496326 133058 526810 133294
rect 527046 133058 571826 133294
rect 572062 133058 572146 133294
rect 572382 133058 586302 133294
rect 586538 133058 586622 133294
rect 586858 133058 586890 133294
rect -2966 132896 586890 133058
rect -6806 130614 590730 130776
rect -6806 130378 -5814 130614
rect -5578 130378 -5494 130614
rect -5258 130378 9266 130614
rect 9502 130378 9586 130614
rect 9822 130378 29266 130614
rect 29502 130378 29586 130614
rect 29822 130378 49266 130614
rect 49502 130378 49586 130614
rect 49822 130378 69266 130614
rect 69502 130378 69586 130614
rect 69822 130378 89266 130614
rect 89502 130378 89586 130614
rect 89822 130378 109266 130614
rect 109502 130378 109586 130614
rect 109822 130378 129266 130614
rect 129502 130378 129586 130614
rect 129822 130378 149266 130614
rect 149502 130378 149586 130614
rect 149822 130378 169266 130614
rect 169502 130378 169586 130614
rect 169822 130378 189266 130614
rect 189502 130378 189586 130614
rect 189822 130378 569266 130614
rect 569502 130378 569586 130614
rect 569822 130378 589182 130614
rect 589418 130378 589502 130614
rect 589738 130378 590730 130614
rect -6806 130216 590730 130378
rect -4886 126954 588810 127116
rect -4886 126718 -3894 126954
rect -3658 126718 -3574 126954
rect -3338 126718 5546 126954
rect 5782 126718 5866 126954
rect 6102 126718 25546 126954
rect 25782 126718 25866 126954
rect 26102 126718 45546 126954
rect 45782 126718 45866 126954
rect 46102 126718 65546 126954
rect 65782 126718 65866 126954
rect 66102 126718 85546 126954
rect 85782 126718 85866 126954
rect 86102 126718 105546 126954
rect 105782 126718 105866 126954
rect 106102 126718 125546 126954
rect 125782 126718 125866 126954
rect 126102 126718 145546 126954
rect 145782 126718 145866 126954
rect 146102 126718 165546 126954
rect 165782 126718 165866 126954
rect 166102 126718 185546 126954
rect 185782 126718 185866 126954
rect 186102 126718 565546 126954
rect 565782 126718 565866 126954
rect 566102 126718 587262 126954
rect 587498 126718 587582 126954
rect 587818 126718 588810 126954
rect -4886 126556 588810 126718
rect -8726 124274 592650 124436
rect -8726 124038 -8694 124274
rect -8458 124038 -8374 124274
rect -8138 124038 22986 124274
rect 23222 124038 23306 124274
rect 23542 124038 42986 124274
rect 43222 124038 43306 124274
rect 43542 124038 62986 124274
rect 63222 124038 63306 124274
rect 63542 124038 82986 124274
rect 83222 124038 83306 124274
rect 83542 124038 102986 124274
rect 103222 124038 103306 124274
rect 103542 124038 122986 124274
rect 123222 124038 123306 124274
rect 123542 124038 142986 124274
rect 143222 124038 143306 124274
rect 143542 124038 162986 124274
rect 163222 124038 163306 124274
rect 163542 124038 182986 124274
rect 183222 124038 183306 124274
rect 183542 124038 562986 124274
rect 563222 124038 563306 124274
rect 563542 124038 592062 124274
rect 592298 124038 592382 124274
rect 592618 124038 592650 124274
rect -8726 123876 592650 124038
rect -2966 123294 586890 123456
rect -2966 123058 -1974 123294
rect -1738 123058 -1654 123294
rect -1418 123058 1826 123294
rect 2062 123058 2146 123294
rect 2382 123058 21826 123294
rect 22062 123058 22146 123294
rect 22382 123058 41826 123294
rect 42062 123058 42146 123294
rect 42382 123058 61826 123294
rect 62062 123058 62146 123294
rect 62382 123058 81826 123294
rect 82062 123058 82146 123294
rect 82382 123058 101826 123294
rect 102062 123058 102146 123294
rect 102382 123058 121826 123294
rect 122062 123058 122146 123294
rect 122382 123058 141826 123294
rect 142062 123058 142146 123294
rect 142382 123058 161826 123294
rect 162062 123058 162146 123294
rect 162382 123058 181826 123294
rect 182062 123058 182146 123294
rect 182382 123058 204250 123294
rect 204486 123058 234970 123294
rect 235206 123058 265690 123294
rect 265926 123058 296410 123294
rect 296646 123058 327130 123294
rect 327366 123058 357850 123294
rect 358086 123058 388570 123294
rect 388806 123058 419290 123294
rect 419526 123058 450010 123294
rect 450246 123058 480730 123294
rect 480966 123058 511450 123294
rect 511686 123058 542170 123294
rect 542406 123058 561826 123294
rect 562062 123058 562146 123294
rect 562382 123058 581826 123294
rect 582062 123058 582146 123294
rect 582382 123058 585342 123294
rect 585578 123058 585662 123294
rect 585898 123058 586890 123294
rect -2966 122896 586890 123058
rect -6806 120614 590730 120776
rect -6806 120378 -6774 120614
rect -6538 120378 -6454 120614
rect -6218 120378 19266 120614
rect 19502 120378 19586 120614
rect 19822 120378 39266 120614
rect 39502 120378 39586 120614
rect 39822 120378 59266 120614
rect 59502 120378 59586 120614
rect 59822 120378 79266 120614
rect 79502 120378 79586 120614
rect 79822 120378 99266 120614
rect 99502 120378 99586 120614
rect 99822 120378 119266 120614
rect 119502 120378 119586 120614
rect 119822 120378 139266 120614
rect 139502 120378 139586 120614
rect 139822 120378 159266 120614
rect 159502 120378 159586 120614
rect 159822 120378 179266 120614
rect 179502 120378 179586 120614
rect 179822 120378 559266 120614
rect 559502 120378 559586 120614
rect 559822 120378 579266 120614
rect 579502 120378 579586 120614
rect 579822 120378 590142 120614
rect 590378 120378 590462 120614
rect 590698 120378 590730 120614
rect -6806 120216 590730 120378
rect -4886 116954 588810 117116
rect -4886 116718 -4854 116954
rect -4618 116718 -4534 116954
rect -4298 116718 15546 116954
rect 15782 116718 15866 116954
rect 16102 116718 35546 116954
rect 35782 116718 35866 116954
rect 36102 116718 55546 116954
rect 55782 116718 55866 116954
rect 56102 116718 75546 116954
rect 75782 116718 75866 116954
rect 76102 116718 95546 116954
rect 95782 116718 95866 116954
rect 96102 116718 115546 116954
rect 115782 116718 115866 116954
rect 116102 116718 135546 116954
rect 135782 116718 135866 116954
rect 136102 116718 155546 116954
rect 155782 116718 155866 116954
rect 156102 116718 175546 116954
rect 175782 116718 175866 116954
rect 176102 116718 195546 116954
rect 195782 116718 195866 116954
rect 196102 116718 575546 116954
rect 575782 116718 575866 116954
rect 576102 116718 588222 116954
rect 588458 116718 588542 116954
rect 588778 116718 588810 116954
rect -4886 116556 588810 116718
rect -8726 114274 592650 114436
rect -8726 114038 -7734 114274
rect -7498 114038 -7414 114274
rect -7178 114038 12986 114274
rect 13222 114038 13306 114274
rect 13542 114038 172986 114274
rect 173222 114038 173306 114274
rect 173542 114038 192986 114274
rect 193222 114038 193306 114274
rect 193542 114038 572986 114274
rect 573222 114038 573306 114274
rect 573542 114038 591102 114274
rect 591338 114038 591422 114274
rect 591658 114038 592650 114274
rect -8726 113876 592650 114038
rect -2966 113294 586890 113456
rect -2966 113058 -2934 113294
rect -2698 113058 -2614 113294
rect -2378 113058 11826 113294
rect 12062 113058 12146 113294
rect 12382 113058 171826 113294
rect 172062 113058 172146 113294
rect 172382 113058 191826 113294
rect 192062 113058 192146 113294
rect 192382 113058 219610 113294
rect 219846 113058 250330 113294
rect 250566 113058 281050 113294
rect 281286 113058 311770 113294
rect 312006 113058 342490 113294
rect 342726 113058 373210 113294
rect 373446 113058 403930 113294
rect 404166 113058 434650 113294
rect 434886 113058 465370 113294
rect 465606 113058 496090 113294
rect 496326 113058 526810 113294
rect 527046 113058 571826 113294
rect 572062 113058 572146 113294
rect 572382 113058 586302 113294
rect 586538 113058 586622 113294
rect 586858 113058 586890 113294
rect -2966 112896 586890 113058
rect -6806 110614 590730 110776
rect -6806 110378 -5814 110614
rect -5578 110378 -5494 110614
rect -5258 110378 9266 110614
rect 9502 110378 9586 110614
rect 9822 110378 169266 110614
rect 169502 110378 169586 110614
rect 169822 110378 189266 110614
rect 189502 110378 189586 110614
rect 189822 110378 569266 110614
rect 569502 110378 569586 110614
rect 569822 110378 589182 110614
rect 589418 110378 589502 110614
rect 589738 110378 590730 110614
rect -6806 110216 590730 110378
rect -4886 106954 588810 107116
rect -4886 106718 -3894 106954
rect -3658 106718 -3574 106954
rect -3338 106718 5546 106954
rect 5782 106718 5866 106954
rect 6102 106718 25546 106954
rect 25782 106718 25866 106954
rect 26102 106718 185546 106954
rect 185782 106718 185866 106954
rect 186102 106718 565546 106954
rect 565782 106718 565866 106954
rect 566102 106718 587262 106954
rect 587498 106718 587582 106954
rect 587818 106718 588810 106954
rect -4886 106556 588810 106718
rect -8726 104274 592650 104436
rect -8726 104038 -8694 104274
rect -8458 104038 -8374 104274
rect -8138 104038 22986 104274
rect 23222 104038 23306 104274
rect 23542 104038 182986 104274
rect 183222 104038 183306 104274
rect 183542 104038 562986 104274
rect 563222 104038 563306 104274
rect 563542 104038 592062 104274
rect 592298 104038 592382 104274
rect 592618 104038 592650 104274
rect -8726 103876 592650 104038
rect -2966 103294 586890 103456
rect -2966 103058 -1974 103294
rect -1738 103058 -1654 103294
rect -1418 103058 1826 103294
rect 2062 103058 2146 103294
rect 2382 103058 21826 103294
rect 22062 103058 22146 103294
rect 22382 103058 31008 103294
rect 31244 103058 165376 103294
rect 165612 103058 181826 103294
rect 182062 103058 182146 103294
rect 182382 103058 204250 103294
rect 204486 103058 234970 103294
rect 235206 103058 265690 103294
rect 265926 103058 296410 103294
rect 296646 103058 327130 103294
rect 327366 103058 357850 103294
rect 358086 103058 388570 103294
rect 388806 103058 419290 103294
rect 419526 103058 450010 103294
rect 450246 103058 480730 103294
rect 480966 103058 511450 103294
rect 511686 103058 542170 103294
rect 542406 103058 561826 103294
rect 562062 103058 562146 103294
rect 562382 103058 581826 103294
rect 582062 103058 582146 103294
rect 582382 103058 585342 103294
rect 585578 103058 585662 103294
rect 585898 103058 586890 103294
rect -2966 102896 586890 103058
rect -6806 100614 590730 100776
rect -6806 100378 -6774 100614
rect -6538 100378 -6454 100614
rect -6218 100378 19266 100614
rect 19502 100378 19586 100614
rect 19822 100378 179266 100614
rect 179502 100378 179586 100614
rect 179822 100378 559266 100614
rect 559502 100378 559586 100614
rect 559822 100378 579266 100614
rect 579502 100378 579586 100614
rect 579822 100378 590142 100614
rect 590378 100378 590462 100614
rect 590698 100378 590730 100614
rect -6806 100216 590730 100378
rect -4886 96954 588810 97116
rect -4886 96718 -4854 96954
rect -4618 96718 -4534 96954
rect -4298 96718 15546 96954
rect 15782 96718 15866 96954
rect 16102 96718 175546 96954
rect 175782 96718 175866 96954
rect 176102 96718 195546 96954
rect 195782 96718 195866 96954
rect 196102 96718 575546 96954
rect 575782 96718 575866 96954
rect 576102 96718 588222 96954
rect 588458 96718 588542 96954
rect 588778 96718 588810 96954
rect -4886 96556 588810 96718
rect -8726 94274 592650 94436
rect -8726 94038 -7734 94274
rect -7498 94038 -7414 94274
rect -7178 94038 12986 94274
rect 13222 94038 13306 94274
rect 13542 94038 172986 94274
rect 173222 94038 173306 94274
rect 173542 94038 192986 94274
rect 193222 94038 193306 94274
rect 193542 94038 572986 94274
rect 573222 94038 573306 94274
rect 573542 94038 591102 94274
rect 591338 94038 591422 94274
rect 591658 94038 592650 94274
rect -8726 93876 592650 94038
rect -2966 93294 586890 93456
rect -2966 93058 -2934 93294
rect -2698 93058 -2614 93294
rect -2378 93058 11826 93294
rect 12062 93058 12146 93294
rect 12382 93058 30328 93294
rect 30564 93058 166056 93294
rect 166292 93058 171826 93294
rect 172062 93058 172146 93294
rect 172382 93058 191826 93294
rect 192062 93058 192146 93294
rect 192382 93058 219610 93294
rect 219846 93058 250330 93294
rect 250566 93058 281050 93294
rect 281286 93058 311770 93294
rect 312006 93058 342490 93294
rect 342726 93058 373210 93294
rect 373446 93058 403930 93294
rect 404166 93058 434650 93294
rect 434886 93058 465370 93294
rect 465606 93058 496090 93294
rect 496326 93058 526810 93294
rect 527046 93058 571826 93294
rect 572062 93058 572146 93294
rect 572382 93058 586302 93294
rect 586538 93058 586622 93294
rect 586858 93058 586890 93294
rect -2966 92896 586890 93058
rect -6806 90614 590730 90776
rect -6806 90378 -5814 90614
rect -5578 90378 -5494 90614
rect -5258 90378 9266 90614
rect 9502 90378 9586 90614
rect 9822 90378 169266 90614
rect 169502 90378 169586 90614
rect 169822 90378 189266 90614
rect 189502 90378 189586 90614
rect 189822 90378 569266 90614
rect 569502 90378 569586 90614
rect 569822 90378 589182 90614
rect 589418 90378 589502 90614
rect 589738 90378 590730 90614
rect -6806 90216 590730 90378
rect -4886 86954 588810 87116
rect -4886 86718 -3894 86954
rect -3658 86718 -3574 86954
rect -3338 86718 5546 86954
rect 5782 86718 5866 86954
rect 6102 86718 25546 86954
rect 25782 86718 25866 86954
rect 26102 86718 185546 86954
rect 185782 86718 185866 86954
rect 186102 86718 565546 86954
rect 565782 86718 565866 86954
rect 566102 86718 587262 86954
rect 587498 86718 587582 86954
rect 587818 86718 588810 86954
rect -4886 86556 588810 86718
rect -8726 84274 592650 84436
rect -8726 84038 -8694 84274
rect -8458 84038 -8374 84274
rect -8138 84038 22986 84274
rect 23222 84038 23306 84274
rect 23542 84038 182986 84274
rect 183222 84038 183306 84274
rect 183542 84038 562986 84274
rect 563222 84038 563306 84274
rect 563542 84038 592062 84274
rect 592298 84038 592382 84274
rect 592618 84038 592650 84274
rect -8726 83876 592650 84038
rect -2966 83294 586890 83456
rect -2966 83058 -1974 83294
rect -1738 83058 -1654 83294
rect -1418 83058 1826 83294
rect 2062 83058 2146 83294
rect 2382 83058 21826 83294
rect 22062 83058 22146 83294
rect 22382 83058 31008 83294
rect 31244 83058 165376 83294
rect 165612 83058 181826 83294
rect 182062 83058 182146 83294
rect 182382 83058 204250 83294
rect 204486 83058 234970 83294
rect 235206 83058 265690 83294
rect 265926 83058 296410 83294
rect 296646 83058 327130 83294
rect 327366 83058 357850 83294
rect 358086 83058 388570 83294
rect 388806 83058 419290 83294
rect 419526 83058 450010 83294
rect 450246 83058 480730 83294
rect 480966 83058 511450 83294
rect 511686 83058 542170 83294
rect 542406 83058 561826 83294
rect 562062 83058 562146 83294
rect 562382 83058 581826 83294
rect 582062 83058 582146 83294
rect 582382 83058 585342 83294
rect 585578 83058 585662 83294
rect 585898 83058 586890 83294
rect -2966 82896 586890 83058
rect -6806 80614 590730 80776
rect -6806 80378 -6774 80614
rect -6538 80378 -6454 80614
rect -6218 80378 19266 80614
rect 19502 80378 19586 80614
rect 19822 80378 179266 80614
rect 179502 80378 179586 80614
rect 179822 80378 559266 80614
rect 559502 80378 559586 80614
rect 559822 80378 579266 80614
rect 579502 80378 579586 80614
rect 579822 80378 590142 80614
rect 590378 80378 590462 80614
rect 590698 80378 590730 80614
rect -6806 80216 590730 80378
rect -4886 76954 588810 77116
rect -4886 76718 -4854 76954
rect -4618 76718 -4534 76954
rect -4298 76718 15546 76954
rect 15782 76718 15866 76954
rect 16102 76718 175546 76954
rect 175782 76718 175866 76954
rect 176102 76718 195546 76954
rect 195782 76718 195866 76954
rect 196102 76718 575546 76954
rect 575782 76718 575866 76954
rect 576102 76718 588222 76954
rect 588458 76718 588542 76954
rect 588778 76718 588810 76954
rect -4886 76556 588810 76718
rect -8726 74274 592650 74436
rect -8726 74038 -7734 74274
rect -7498 74038 -7414 74274
rect -7178 74038 12986 74274
rect 13222 74038 13306 74274
rect 13542 74038 172986 74274
rect 173222 74038 173306 74274
rect 173542 74038 192986 74274
rect 193222 74038 193306 74274
rect 193542 74038 572986 74274
rect 573222 74038 573306 74274
rect 573542 74038 591102 74274
rect 591338 74038 591422 74274
rect 591658 74038 592650 74274
rect -8726 73876 592650 74038
rect -2966 73294 586890 73456
rect -2966 73058 -2934 73294
rect -2698 73058 -2614 73294
rect -2378 73058 11826 73294
rect 12062 73058 12146 73294
rect 12382 73058 30328 73294
rect 30564 73058 166056 73294
rect 166292 73058 171826 73294
rect 172062 73058 172146 73294
rect 172382 73058 191826 73294
rect 192062 73058 192146 73294
rect 192382 73058 219610 73294
rect 219846 73058 250330 73294
rect 250566 73058 281050 73294
rect 281286 73058 311770 73294
rect 312006 73058 342490 73294
rect 342726 73058 373210 73294
rect 373446 73058 403930 73294
rect 404166 73058 434650 73294
rect 434886 73058 465370 73294
rect 465606 73058 496090 73294
rect 496326 73058 526810 73294
rect 527046 73058 571826 73294
rect 572062 73058 572146 73294
rect 572382 73058 586302 73294
rect 586538 73058 586622 73294
rect 586858 73058 586890 73294
rect -2966 72896 586890 73058
rect -6806 70614 590730 70776
rect -6806 70378 -5814 70614
rect -5578 70378 -5494 70614
rect -5258 70378 9266 70614
rect 9502 70378 9586 70614
rect 9822 70378 169266 70614
rect 169502 70378 169586 70614
rect 169822 70378 189266 70614
rect 189502 70378 189586 70614
rect 189822 70378 569266 70614
rect 569502 70378 569586 70614
rect 569822 70378 589182 70614
rect 589418 70378 589502 70614
rect 589738 70378 590730 70614
rect -6806 70216 590730 70378
rect -4886 66954 588810 67116
rect -4886 66718 -3894 66954
rect -3658 66718 -3574 66954
rect -3338 66718 5546 66954
rect 5782 66718 5866 66954
rect 6102 66718 25546 66954
rect 25782 66718 25866 66954
rect 26102 66718 185546 66954
rect 185782 66718 185866 66954
rect 186102 66718 565546 66954
rect 565782 66718 565866 66954
rect 566102 66718 587262 66954
rect 587498 66718 587582 66954
rect 587818 66718 588810 66954
rect -4886 66556 588810 66718
rect -8726 64274 592650 64436
rect -8726 64038 -8694 64274
rect -8458 64038 -8374 64274
rect -8138 64038 22986 64274
rect 23222 64038 23306 64274
rect 23542 64038 182986 64274
rect 183222 64038 183306 64274
rect 183542 64038 562986 64274
rect 563222 64038 563306 64274
rect 563542 64038 592062 64274
rect 592298 64038 592382 64274
rect 592618 64038 592650 64274
rect -8726 63876 592650 64038
rect -2966 63294 586890 63456
rect -2966 63058 -1974 63294
rect -1738 63058 -1654 63294
rect -1418 63058 1826 63294
rect 2062 63058 2146 63294
rect 2382 63058 21826 63294
rect 22062 63058 22146 63294
rect 22382 63058 31008 63294
rect 31244 63058 165376 63294
rect 165612 63058 181826 63294
rect 182062 63058 182146 63294
rect 182382 63058 204250 63294
rect 204486 63058 234970 63294
rect 235206 63058 265690 63294
rect 265926 63058 296410 63294
rect 296646 63058 327130 63294
rect 327366 63058 357850 63294
rect 358086 63058 388570 63294
rect 388806 63058 419290 63294
rect 419526 63058 450010 63294
rect 450246 63058 480730 63294
rect 480966 63058 511450 63294
rect 511686 63058 542170 63294
rect 542406 63058 561826 63294
rect 562062 63058 562146 63294
rect 562382 63058 581826 63294
rect 582062 63058 582146 63294
rect 582382 63058 585342 63294
rect 585578 63058 585662 63294
rect 585898 63058 586890 63294
rect -2966 62896 586890 63058
rect -6806 60614 590730 60776
rect -6806 60378 -6774 60614
rect -6538 60378 -6454 60614
rect -6218 60378 19266 60614
rect 19502 60378 19586 60614
rect 19822 60378 179266 60614
rect 179502 60378 179586 60614
rect 179822 60378 559266 60614
rect 559502 60378 559586 60614
rect 559822 60378 579266 60614
rect 579502 60378 579586 60614
rect 579822 60378 590142 60614
rect 590378 60378 590462 60614
rect 590698 60378 590730 60614
rect -6806 60216 590730 60378
rect -4886 56954 588810 57116
rect -4886 56718 -4854 56954
rect -4618 56718 -4534 56954
rect -4298 56718 15546 56954
rect 15782 56718 15866 56954
rect 16102 56718 175546 56954
rect 175782 56718 175866 56954
rect 176102 56718 195546 56954
rect 195782 56718 195866 56954
rect 196102 56718 215546 56954
rect 215782 56718 215866 56954
rect 216102 56718 235546 56954
rect 235782 56718 235866 56954
rect 236102 56718 255546 56954
rect 255782 56718 255866 56954
rect 256102 56718 275546 56954
rect 275782 56718 275866 56954
rect 276102 56718 295546 56954
rect 295782 56718 295866 56954
rect 296102 56718 315546 56954
rect 315782 56718 315866 56954
rect 316102 56718 335546 56954
rect 335782 56718 335866 56954
rect 336102 56718 355546 56954
rect 355782 56718 355866 56954
rect 356102 56718 375546 56954
rect 375782 56718 375866 56954
rect 376102 56718 395546 56954
rect 395782 56718 395866 56954
rect 396102 56718 415546 56954
rect 415782 56718 415866 56954
rect 416102 56718 435546 56954
rect 435782 56718 435866 56954
rect 436102 56718 455546 56954
rect 455782 56718 455866 56954
rect 456102 56718 475546 56954
rect 475782 56718 475866 56954
rect 476102 56718 495546 56954
rect 495782 56718 495866 56954
rect 496102 56718 515546 56954
rect 515782 56718 515866 56954
rect 516102 56718 535546 56954
rect 535782 56718 535866 56954
rect 536102 56718 555546 56954
rect 555782 56718 555866 56954
rect 556102 56718 575546 56954
rect 575782 56718 575866 56954
rect 576102 56718 588222 56954
rect 588458 56718 588542 56954
rect 588778 56718 588810 56954
rect -4886 56556 588810 56718
rect -8726 54274 592650 54436
rect -8726 54038 -7734 54274
rect -7498 54038 -7414 54274
rect -7178 54038 12986 54274
rect 13222 54038 13306 54274
rect 13542 54038 172986 54274
rect 173222 54038 173306 54274
rect 173542 54038 192986 54274
rect 193222 54038 193306 54274
rect 193542 54038 212986 54274
rect 213222 54038 213306 54274
rect 213542 54038 232986 54274
rect 233222 54038 233306 54274
rect 233542 54038 252986 54274
rect 253222 54038 253306 54274
rect 253542 54038 272986 54274
rect 273222 54038 273306 54274
rect 273542 54038 292986 54274
rect 293222 54038 293306 54274
rect 293542 54038 312986 54274
rect 313222 54038 313306 54274
rect 313542 54038 332986 54274
rect 333222 54038 333306 54274
rect 333542 54038 352986 54274
rect 353222 54038 353306 54274
rect 353542 54038 372986 54274
rect 373222 54038 373306 54274
rect 373542 54038 392986 54274
rect 393222 54038 393306 54274
rect 393542 54038 412986 54274
rect 413222 54038 413306 54274
rect 413542 54038 432986 54274
rect 433222 54038 433306 54274
rect 433542 54038 452986 54274
rect 453222 54038 453306 54274
rect 453542 54038 472986 54274
rect 473222 54038 473306 54274
rect 473542 54038 492986 54274
rect 493222 54038 493306 54274
rect 493542 54038 512986 54274
rect 513222 54038 513306 54274
rect 513542 54038 532986 54274
rect 533222 54038 533306 54274
rect 533542 54038 552986 54274
rect 553222 54038 553306 54274
rect 553542 54038 572986 54274
rect 573222 54038 573306 54274
rect 573542 54038 591102 54274
rect 591338 54038 591422 54274
rect 591658 54038 592650 54274
rect -8726 53876 592650 54038
rect -2966 53294 586890 53456
rect -2966 53058 -2934 53294
rect -2698 53058 -2614 53294
rect -2378 53058 11826 53294
rect 12062 53058 12146 53294
rect 12382 53058 30328 53294
rect 30564 53058 166056 53294
rect 166292 53058 171826 53294
rect 172062 53058 172146 53294
rect 172382 53058 191826 53294
rect 192062 53058 192146 53294
rect 192382 53058 211826 53294
rect 212062 53058 212146 53294
rect 212382 53058 231826 53294
rect 232062 53058 232146 53294
rect 232382 53058 251826 53294
rect 252062 53058 252146 53294
rect 252382 53058 271826 53294
rect 272062 53058 272146 53294
rect 272382 53058 291826 53294
rect 292062 53058 292146 53294
rect 292382 53058 311826 53294
rect 312062 53058 312146 53294
rect 312382 53058 331826 53294
rect 332062 53058 332146 53294
rect 332382 53058 351826 53294
rect 352062 53058 352146 53294
rect 352382 53058 371826 53294
rect 372062 53058 372146 53294
rect 372382 53058 391826 53294
rect 392062 53058 392146 53294
rect 392382 53058 411826 53294
rect 412062 53058 412146 53294
rect 412382 53058 431826 53294
rect 432062 53058 432146 53294
rect 432382 53058 451826 53294
rect 452062 53058 452146 53294
rect 452382 53058 471826 53294
rect 472062 53058 472146 53294
rect 472382 53058 491826 53294
rect 492062 53058 492146 53294
rect 492382 53058 511826 53294
rect 512062 53058 512146 53294
rect 512382 53058 531826 53294
rect 532062 53058 532146 53294
rect 532382 53058 551826 53294
rect 552062 53058 552146 53294
rect 552382 53058 571826 53294
rect 572062 53058 572146 53294
rect 572382 53058 586302 53294
rect 586538 53058 586622 53294
rect 586858 53058 586890 53294
rect -2966 52896 586890 53058
rect -6806 50614 590730 50776
rect -6806 50378 -5814 50614
rect -5578 50378 -5494 50614
rect -5258 50378 9266 50614
rect 9502 50378 9586 50614
rect 9822 50378 169266 50614
rect 169502 50378 169586 50614
rect 169822 50378 189266 50614
rect 189502 50378 189586 50614
rect 189822 50378 209266 50614
rect 209502 50378 209586 50614
rect 209822 50378 229266 50614
rect 229502 50378 229586 50614
rect 229822 50378 249266 50614
rect 249502 50378 249586 50614
rect 249822 50378 269266 50614
rect 269502 50378 269586 50614
rect 269822 50378 289266 50614
rect 289502 50378 289586 50614
rect 289822 50378 309266 50614
rect 309502 50378 309586 50614
rect 309822 50378 329266 50614
rect 329502 50378 329586 50614
rect 329822 50378 349266 50614
rect 349502 50378 349586 50614
rect 349822 50378 369266 50614
rect 369502 50378 369586 50614
rect 369822 50378 389266 50614
rect 389502 50378 389586 50614
rect 389822 50378 409266 50614
rect 409502 50378 409586 50614
rect 409822 50378 429266 50614
rect 429502 50378 429586 50614
rect 429822 50378 449266 50614
rect 449502 50378 449586 50614
rect 449822 50378 469266 50614
rect 469502 50378 469586 50614
rect 469822 50378 489266 50614
rect 489502 50378 489586 50614
rect 489822 50378 509266 50614
rect 509502 50378 509586 50614
rect 509822 50378 529266 50614
rect 529502 50378 529586 50614
rect 529822 50378 549266 50614
rect 549502 50378 549586 50614
rect 549822 50378 569266 50614
rect 569502 50378 569586 50614
rect 569822 50378 589182 50614
rect 589418 50378 589502 50614
rect 589738 50378 590730 50614
rect -6806 50216 590730 50378
rect -4886 46954 588810 47116
rect -4886 46718 -3894 46954
rect -3658 46718 -3574 46954
rect -3338 46718 5546 46954
rect 5782 46718 5866 46954
rect 6102 46718 25546 46954
rect 25782 46718 25866 46954
rect 26102 46718 185546 46954
rect 185782 46718 185866 46954
rect 186102 46718 205546 46954
rect 205782 46718 205866 46954
rect 206102 46718 225546 46954
rect 225782 46718 225866 46954
rect 226102 46718 245546 46954
rect 245782 46718 245866 46954
rect 246102 46718 265546 46954
rect 265782 46718 265866 46954
rect 266102 46718 285546 46954
rect 285782 46718 285866 46954
rect 286102 46718 305546 46954
rect 305782 46718 305866 46954
rect 306102 46718 325546 46954
rect 325782 46718 325866 46954
rect 326102 46718 345546 46954
rect 345782 46718 345866 46954
rect 346102 46718 365546 46954
rect 365782 46718 365866 46954
rect 366102 46718 385546 46954
rect 385782 46718 385866 46954
rect 386102 46718 405546 46954
rect 405782 46718 405866 46954
rect 406102 46718 425546 46954
rect 425782 46718 425866 46954
rect 426102 46718 445546 46954
rect 445782 46718 445866 46954
rect 446102 46718 465546 46954
rect 465782 46718 465866 46954
rect 466102 46718 485546 46954
rect 485782 46718 485866 46954
rect 486102 46718 505546 46954
rect 505782 46718 505866 46954
rect 506102 46718 525546 46954
rect 525782 46718 525866 46954
rect 526102 46718 545546 46954
rect 545782 46718 545866 46954
rect 546102 46718 565546 46954
rect 565782 46718 565866 46954
rect 566102 46718 587262 46954
rect 587498 46718 587582 46954
rect 587818 46718 588810 46954
rect -4886 46556 588810 46718
rect -8726 44274 592650 44436
rect -8726 44038 -8694 44274
rect -8458 44038 -8374 44274
rect -8138 44038 22986 44274
rect 23222 44038 23306 44274
rect 23542 44038 182986 44274
rect 183222 44038 183306 44274
rect 183542 44038 202986 44274
rect 203222 44038 203306 44274
rect 203542 44038 222986 44274
rect 223222 44038 223306 44274
rect 223542 44038 242986 44274
rect 243222 44038 243306 44274
rect 243542 44038 262986 44274
rect 263222 44038 263306 44274
rect 263542 44038 282986 44274
rect 283222 44038 283306 44274
rect 283542 44038 302986 44274
rect 303222 44038 303306 44274
rect 303542 44038 322986 44274
rect 323222 44038 323306 44274
rect 323542 44038 342986 44274
rect 343222 44038 343306 44274
rect 343542 44038 362986 44274
rect 363222 44038 363306 44274
rect 363542 44038 382986 44274
rect 383222 44038 383306 44274
rect 383542 44038 402986 44274
rect 403222 44038 403306 44274
rect 403542 44038 422986 44274
rect 423222 44038 423306 44274
rect 423542 44038 442986 44274
rect 443222 44038 443306 44274
rect 443542 44038 462986 44274
rect 463222 44038 463306 44274
rect 463542 44038 482986 44274
rect 483222 44038 483306 44274
rect 483542 44038 502986 44274
rect 503222 44038 503306 44274
rect 503542 44038 522986 44274
rect 523222 44038 523306 44274
rect 523542 44038 542986 44274
rect 543222 44038 543306 44274
rect 543542 44038 562986 44274
rect 563222 44038 563306 44274
rect 563542 44038 592062 44274
rect 592298 44038 592382 44274
rect 592618 44038 592650 44274
rect -8726 43876 592650 44038
rect -2966 43294 586890 43456
rect -2966 43058 -1974 43294
rect -1738 43058 -1654 43294
rect -1418 43058 1826 43294
rect 2062 43058 2146 43294
rect 2382 43058 21826 43294
rect 22062 43058 22146 43294
rect 22382 43058 31008 43294
rect 31244 43058 165376 43294
rect 165612 43058 181826 43294
rect 182062 43058 182146 43294
rect 182382 43058 201826 43294
rect 202062 43058 202146 43294
rect 202382 43058 221826 43294
rect 222062 43058 222146 43294
rect 222382 43058 241826 43294
rect 242062 43058 242146 43294
rect 242382 43058 261826 43294
rect 262062 43058 262146 43294
rect 262382 43058 281826 43294
rect 282062 43058 282146 43294
rect 282382 43058 301826 43294
rect 302062 43058 302146 43294
rect 302382 43058 321826 43294
rect 322062 43058 322146 43294
rect 322382 43058 341826 43294
rect 342062 43058 342146 43294
rect 342382 43058 361826 43294
rect 362062 43058 362146 43294
rect 362382 43058 381826 43294
rect 382062 43058 382146 43294
rect 382382 43058 401826 43294
rect 402062 43058 402146 43294
rect 402382 43058 421826 43294
rect 422062 43058 422146 43294
rect 422382 43058 441826 43294
rect 442062 43058 442146 43294
rect 442382 43058 461826 43294
rect 462062 43058 462146 43294
rect 462382 43058 481826 43294
rect 482062 43058 482146 43294
rect 482382 43058 501826 43294
rect 502062 43058 502146 43294
rect 502382 43058 521826 43294
rect 522062 43058 522146 43294
rect 522382 43058 541826 43294
rect 542062 43058 542146 43294
rect 542382 43058 561826 43294
rect 562062 43058 562146 43294
rect 562382 43058 581826 43294
rect 582062 43058 582146 43294
rect 582382 43058 585342 43294
rect 585578 43058 585662 43294
rect 585898 43058 586890 43294
rect -2966 42896 586890 43058
rect -6806 40614 590730 40776
rect -6806 40378 -6774 40614
rect -6538 40378 -6454 40614
rect -6218 40378 19266 40614
rect 19502 40378 19586 40614
rect 19822 40378 179266 40614
rect 179502 40378 179586 40614
rect 179822 40378 199266 40614
rect 199502 40378 199586 40614
rect 199822 40378 219266 40614
rect 219502 40378 219586 40614
rect 219822 40378 239266 40614
rect 239502 40378 239586 40614
rect 239822 40378 259266 40614
rect 259502 40378 259586 40614
rect 259822 40378 279266 40614
rect 279502 40378 279586 40614
rect 279822 40378 299266 40614
rect 299502 40378 299586 40614
rect 299822 40378 319266 40614
rect 319502 40378 319586 40614
rect 319822 40378 339266 40614
rect 339502 40378 339586 40614
rect 339822 40378 359266 40614
rect 359502 40378 359586 40614
rect 359822 40378 379266 40614
rect 379502 40378 379586 40614
rect 379822 40378 399266 40614
rect 399502 40378 399586 40614
rect 399822 40378 419266 40614
rect 419502 40378 419586 40614
rect 419822 40378 439266 40614
rect 439502 40378 439586 40614
rect 439822 40378 459266 40614
rect 459502 40378 459586 40614
rect 459822 40378 479266 40614
rect 479502 40378 479586 40614
rect 479822 40378 499266 40614
rect 499502 40378 499586 40614
rect 499822 40378 519266 40614
rect 519502 40378 519586 40614
rect 519822 40378 539266 40614
rect 539502 40378 539586 40614
rect 539822 40378 559266 40614
rect 559502 40378 559586 40614
rect 559822 40378 579266 40614
rect 579502 40378 579586 40614
rect 579822 40378 590142 40614
rect 590378 40378 590462 40614
rect 590698 40378 590730 40614
rect -6806 40216 590730 40378
rect -4886 36954 588810 37116
rect -4886 36718 -4854 36954
rect -4618 36718 -4534 36954
rect -4298 36718 15546 36954
rect 15782 36718 15866 36954
rect 16102 36718 175546 36954
rect 175782 36718 175866 36954
rect 176102 36718 195546 36954
rect 195782 36718 195866 36954
rect 196102 36718 215546 36954
rect 215782 36718 215866 36954
rect 216102 36718 235546 36954
rect 235782 36718 235866 36954
rect 236102 36718 255546 36954
rect 255782 36718 255866 36954
rect 256102 36718 275546 36954
rect 275782 36718 275866 36954
rect 276102 36718 295546 36954
rect 295782 36718 295866 36954
rect 296102 36718 315546 36954
rect 315782 36718 315866 36954
rect 316102 36718 335546 36954
rect 335782 36718 335866 36954
rect 336102 36718 355546 36954
rect 355782 36718 355866 36954
rect 356102 36718 375546 36954
rect 375782 36718 375866 36954
rect 376102 36718 395546 36954
rect 395782 36718 395866 36954
rect 396102 36718 415546 36954
rect 415782 36718 415866 36954
rect 416102 36718 435546 36954
rect 435782 36718 435866 36954
rect 436102 36718 455546 36954
rect 455782 36718 455866 36954
rect 456102 36718 475546 36954
rect 475782 36718 475866 36954
rect 476102 36718 495546 36954
rect 495782 36718 495866 36954
rect 496102 36718 515546 36954
rect 515782 36718 515866 36954
rect 516102 36718 535546 36954
rect 535782 36718 535866 36954
rect 536102 36718 555546 36954
rect 555782 36718 555866 36954
rect 556102 36718 575546 36954
rect 575782 36718 575866 36954
rect 576102 36718 588222 36954
rect 588458 36718 588542 36954
rect 588778 36718 588810 36954
rect -4886 36556 588810 36718
rect -8726 34274 592650 34436
rect -8726 34038 -7734 34274
rect -7498 34038 -7414 34274
rect -7178 34038 12986 34274
rect 13222 34038 13306 34274
rect 13542 34038 172986 34274
rect 173222 34038 173306 34274
rect 173542 34038 192986 34274
rect 193222 34038 193306 34274
rect 193542 34038 212986 34274
rect 213222 34038 213306 34274
rect 213542 34038 232986 34274
rect 233222 34038 233306 34274
rect 233542 34038 252986 34274
rect 253222 34038 253306 34274
rect 253542 34038 272986 34274
rect 273222 34038 273306 34274
rect 273542 34038 292986 34274
rect 293222 34038 293306 34274
rect 293542 34038 312986 34274
rect 313222 34038 313306 34274
rect 313542 34038 332986 34274
rect 333222 34038 333306 34274
rect 333542 34038 352986 34274
rect 353222 34038 353306 34274
rect 353542 34038 372986 34274
rect 373222 34038 373306 34274
rect 373542 34038 392986 34274
rect 393222 34038 393306 34274
rect 393542 34038 412986 34274
rect 413222 34038 413306 34274
rect 413542 34038 432986 34274
rect 433222 34038 433306 34274
rect 433542 34038 452986 34274
rect 453222 34038 453306 34274
rect 453542 34038 472986 34274
rect 473222 34038 473306 34274
rect 473542 34038 492986 34274
rect 493222 34038 493306 34274
rect 493542 34038 512986 34274
rect 513222 34038 513306 34274
rect 513542 34038 532986 34274
rect 533222 34038 533306 34274
rect 533542 34038 552986 34274
rect 553222 34038 553306 34274
rect 553542 34038 572986 34274
rect 573222 34038 573306 34274
rect 573542 34038 591102 34274
rect 591338 34038 591422 34274
rect 591658 34038 592650 34274
rect -8726 33876 592650 34038
rect -2966 33294 586890 33456
rect -2966 33058 -2934 33294
rect -2698 33058 -2614 33294
rect -2378 33058 11826 33294
rect 12062 33058 12146 33294
rect 12382 33058 30328 33294
rect 30564 33058 166056 33294
rect 166292 33058 171826 33294
rect 172062 33058 172146 33294
rect 172382 33058 191826 33294
rect 192062 33058 192146 33294
rect 192382 33058 211826 33294
rect 212062 33058 212146 33294
rect 212382 33058 231826 33294
rect 232062 33058 232146 33294
rect 232382 33058 251826 33294
rect 252062 33058 252146 33294
rect 252382 33058 271826 33294
rect 272062 33058 272146 33294
rect 272382 33058 291826 33294
rect 292062 33058 292146 33294
rect 292382 33058 311826 33294
rect 312062 33058 312146 33294
rect 312382 33058 331826 33294
rect 332062 33058 332146 33294
rect 332382 33058 351826 33294
rect 352062 33058 352146 33294
rect 352382 33058 371826 33294
rect 372062 33058 372146 33294
rect 372382 33058 391826 33294
rect 392062 33058 392146 33294
rect 392382 33058 411826 33294
rect 412062 33058 412146 33294
rect 412382 33058 431826 33294
rect 432062 33058 432146 33294
rect 432382 33058 451826 33294
rect 452062 33058 452146 33294
rect 452382 33058 471826 33294
rect 472062 33058 472146 33294
rect 472382 33058 491826 33294
rect 492062 33058 492146 33294
rect 492382 33058 511826 33294
rect 512062 33058 512146 33294
rect 512382 33058 531826 33294
rect 532062 33058 532146 33294
rect 532382 33058 551826 33294
rect 552062 33058 552146 33294
rect 552382 33058 571826 33294
rect 572062 33058 572146 33294
rect 572382 33058 586302 33294
rect 586538 33058 586622 33294
rect 586858 33058 586890 33294
rect -2966 32896 586890 33058
rect -6806 30614 590730 30776
rect -6806 30378 -5814 30614
rect -5578 30378 -5494 30614
rect -5258 30378 9266 30614
rect 9502 30378 9586 30614
rect 9822 30378 169266 30614
rect 169502 30378 169586 30614
rect 169822 30378 189266 30614
rect 189502 30378 189586 30614
rect 189822 30378 209266 30614
rect 209502 30378 209586 30614
rect 209822 30378 229266 30614
rect 229502 30378 229586 30614
rect 229822 30378 249266 30614
rect 249502 30378 249586 30614
rect 249822 30378 269266 30614
rect 269502 30378 269586 30614
rect 269822 30378 289266 30614
rect 289502 30378 289586 30614
rect 289822 30378 309266 30614
rect 309502 30378 309586 30614
rect 309822 30378 329266 30614
rect 329502 30378 329586 30614
rect 329822 30378 349266 30614
rect 349502 30378 349586 30614
rect 349822 30378 369266 30614
rect 369502 30378 369586 30614
rect 369822 30378 389266 30614
rect 389502 30378 389586 30614
rect 389822 30378 409266 30614
rect 409502 30378 409586 30614
rect 409822 30378 429266 30614
rect 429502 30378 429586 30614
rect 429822 30378 449266 30614
rect 449502 30378 449586 30614
rect 449822 30378 469266 30614
rect 469502 30378 469586 30614
rect 469822 30378 489266 30614
rect 489502 30378 489586 30614
rect 489822 30378 509266 30614
rect 509502 30378 509586 30614
rect 509822 30378 529266 30614
rect 529502 30378 529586 30614
rect 529822 30378 549266 30614
rect 549502 30378 549586 30614
rect 549822 30378 569266 30614
rect 569502 30378 569586 30614
rect 569822 30378 589182 30614
rect 589418 30378 589502 30614
rect 589738 30378 590730 30614
rect -6806 30216 590730 30378
rect -4886 26954 588810 27116
rect -4886 26718 -3894 26954
rect -3658 26718 -3574 26954
rect -3338 26718 5546 26954
rect 5782 26718 5866 26954
rect 6102 26718 25546 26954
rect 25782 26718 25866 26954
rect 26102 26718 45546 26954
rect 45782 26718 45866 26954
rect 46102 26718 65546 26954
rect 65782 26718 65866 26954
rect 66102 26718 85546 26954
rect 85782 26718 85866 26954
rect 86102 26718 105546 26954
rect 105782 26718 105866 26954
rect 106102 26718 125546 26954
rect 125782 26718 125866 26954
rect 126102 26718 145546 26954
rect 145782 26718 145866 26954
rect 146102 26718 165546 26954
rect 165782 26718 165866 26954
rect 166102 26718 185546 26954
rect 185782 26718 185866 26954
rect 186102 26718 205546 26954
rect 205782 26718 205866 26954
rect 206102 26718 225546 26954
rect 225782 26718 225866 26954
rect 226102 26718 245546 26954
rect 245782 26718 245866 26954
rect 246102 26718 265546 26954
rect 265782 26718 265866 26954
rect 266102 26718 285546 26954
rect 285782 26718 285866 26954
rect 286102 26718 305546 26954
rect 305782 26718 305866 26954
rect 306102 26718 325546 26954
rect 325782 26718 325866 26954
rect 326102 26718 345546 26954
rect 345782 26718 345866 26954
rect 346102 26718 365546 26954
rect 365782 26718 365866 26954
rect 366102 26718 385546 26954
rect 385782 26718 385866 26954
rect 386102 26718 405546 26954
rect 405782 26718 405866 26954
rect 406102 26718 425546 26954
rect 425782 26718 425866 26954
rect 426102 26718 445546 26954
rect 445782 26718 445866 26954
rect 446102 26718 465546 26954
rect 465782 26718 465866 26954
rect 466102 26718 485546 26954
rect 485782 26718 485866 26954
rect 486102 26718 505546 26954
rect 505782 26718 505866 26954
rect 506102 26718 525546 26954
rect 525782 26718 525866 26954
rect 526102 26718 545546 26954
rect 545782 26718 545866 26954
rect 546102 26718 565546 26954
rect 565782 26718 565866 26954
rect 566102 26718 587262 26954
rect 587498 26718 587582 26954
rect 587818 26718 588810 26954
rect -4886 26556 588810 26718
rect -8726 24274 592650 24436
rect -8726 24038 -8694 24274
rect -8458 24038 -8374 24274
rect -8138 24038 22986 24274
rect 23222 24038 23306 24274
rect 23542 24038 42986 24274
rect 43222 24038 43306 24274
rect 43542 24038 62986 24274
rect 63222 24038 63306 24274
rect 63542 24038 82986 24274
rect 83222 24038 83306 24274
rect 83542 24038 102986 24274
rect 103222 24038 103306 24274
rect 103542 24038 122986 24274
rect 123222 24038 123306 24274
rect 123542 24038 142986 24274
rect 143222 24038 143306 24274
rect 143542 24038 162986 24274
rect 163222 24038 163306 24274
rect 163542 24038 182986 24274
rect 183222 24038 183306 24274
rect 183542 24038 202986 24274
rect 203222 24038 203306 24274
rect 203542 24038 222986 24274
rect 223222 24038 223306 24274
rect 223542 24038 242986 24274
rect 243222 24038 243306 24274
rect 243542 24038 262986 24274
rect 263222 24038 263306 24274
rect 263542 24038 282986 24274
rect 283222 24038 283306 24274
rect 283542 24038 302986 24274
rect 303222 24038 303306 24274
rect 303542 24038 322986 24274
rect 323222 24038 323306 24274
rect 323542 24038 342986 24274
rect 343222 24038 343306 24274
rect 343542 24038 362986 24274
rect 363222 24038 363306 24274
rect 363542 24038 382986 24274
rect 383222 24038 383306 24274
rect 383542 24038 402986 24274
rect 403222 24038 403306 24274
rect 403542 24038 422986 24274
rect 423222 24038 423306 24274
rect 423542 24038 442986 24274
rect 443222 24038 443306 24274
rect 443542 24038 462986 24274
rect 463222 24038 463306 24274
rect 463542 24038 482986 24274
rect 483222 24038 483306 24274
rect 483542 24038 502986 24274
rect 503222 24038 503306 24274
rect 503542 24038 522986 24274
rect 523222 24038 523306 24274
rect 523542 24038 542986 24274
rect 543222 24038 543306 24274
rect 543542 24038 562986 24274
rect 563222 24038 563306 24274
rect 563542 24038 592062 24274
rect 592298 24038 592382 24274
rect 592618 24038 592650 24274
rect -8726 23876 592650 24038
rect -2966 23294 586890 23456
rect -2966 23058 -1974 23294
rect -1738 23058 -1654 23294
rect -1418 23058 1826 23294
rect 2062 23058 2146 23294
rect 2382 23058 21826 23294
rect 22062 23058 22146 23294
rect 22382 23058 41826 23294
rect 42062 23058 42146 23294
rect 42382 23058 61826 23294
rect 62062 23058 62146 23294
rect 62382 23058 81826 23294
rect 82062 23058 82146 23294
rect 82382 23058 101826 23294
rect 102062 23058 102146 23294
rect 102382 23058 121826 23294
rect 122062 23058 122146 23294
rect 122382 23058 141826 23294
rect 142062 23058 142146 23294
rect 142382 23058 161826 23294
rect 162062 23058 162146 23294
rect 162382 23058 181826 23294
rect 182062 23058 182146 23294
rect 182382 23058 201826 23294
rect 202062 23058 202146 23294
rect 202382 23058 221826 23294
rect 222062 23058 222146 23294
rect 222382 23058 241826 23294
rect 242062 23058 242146 23294
rect 242382 23058 261826 23294
rect 262062 23058 262146 23294
rect 262382 23058 281826 23294
rect 282062 23058 282146 23294
rect 282382 23058 301826 23294
rect 302062 23058 302146 23294
rect 302382 23058 321826 23294
rect 322062 23058 322146 23294
rect 322382 23058 341826 23294
rect 342062 23058 342146 23294
rect 342382 23058 361826 23294
rect 362062 23058 362146 23294
rect 362382 23058 381826 23294
rect 382062 23058 382146 23294
rect 382382 23058 401826 23294
rect 402062 23058 402146 23294
rect 402382 23058 421826 23294
rect 422062 23058 422146 23294
rect 422382 23058 441826 23294
rect 442062 23058 442146 23294
rect 442382 23058 461826 23294
rect 462062 23058 462146 23294
rect 462382 23058 481826 23294
rect 482062 23058 482146 23294
rect 482382 23058 501826 23294
rect 502062 23058 502146 23294
rect 502382 23058 521826 23294
rect 522062 23058 522146 23294
rect 522382 23058 541826 23294
rect 542062 23058 542146 23294
rect 542382 23058 561826 23294
rect 562062 23058 562146 23294
rect 562382 23058 581826 23294
rect 582062 23058 582146 23294
rect 582382 23058 585342 23294
rect 585578 23058 585662 23294
rect 585898 23058 586890 23294
rect -2966 22896 586890 23058
rect -6806 20614 590730 20776
rect -6806 20378 -6774 20614
rect -6538 20378 -6454 20614
rect -6218 20378 19266 20614
rect 19502 20378 19586 20614
rect 19822 20378 39266 20614
rect 39502 20378 39586 20614
rect 39822 20378 59266 20614
rect 59502 20378 59586 20614
rect 59822 20378 79266 20614
rect 79502 20378 79586 20614
rect 79822 20378 99266 20614
rect 99502 20378 99586 20614
rect 99822 20378 119266 20614
rect 119502 20378 119586 20614
rect 119822 20378 139266 20614
rect 139502 20378 139586 20614
rect 139822 20378 159266 20614
rect 159502 20378 159586 20614
rect 159822 20378 179266 20614
rect 179502 20378 179586 20614
rect 179822 20378 199266 20614
rect 199502 20378 199586 20614
rect 199822 20378 219266 20614
rect 219502 20378 219586 20614
rect 219822 20378 239266 20614
rect 239502 20378 239586 20614
rect 239822 20378 259266 20614
rect 259502 20378 259586 20614
rect 259822 20378 279266 20614
rect 279502 20378 279586 20614
rect 279822 20378 299266 20614
rect 299502 20378 299586 20614
rect 299822 20378 319266 20614
rect 319502 20378 319586 20614
rect 319822 20378 339266 20614
rect 339502 20378 339586 20614
rect 339822 20378 359266 20614
rect 359502 20378 359586 20614
rect 359822 20378 379266 20614
rect 379502 20378 379586 20614
rect 379822 20378 399266 20614
rect 399502 20378 399586 20614
rect 399822 20378 419266 20614
rect 419502 20378 419586 20614
rect 419822 20378 439266 20614
rect 439502 20378 439586 20614
rect 439822 20378 459266 20614
rect 459502 20378 459586 20614
rect 459822 20378 479266 20614
rect 479502 20378 479586 20614
rect 479822 20378 499266 20614
rect 499502 20378 499586 20614
rect 499822 20378 519266 20614
rect 519502 20378 519586 20614
rect 519822 20378 539266 20614
rect 539502 20378 539586 20614
rect 539822 20378 559266 20614
rect 559502 20378 559586 20614
rect 559822 20378 579266 20614
rect 579502 20378 579586 20614
rect 579822 20378 590142 20614
rect 590378 20378 590462 20614
rect 590698 20378 590730 20614
rect -6806 20216 590730 20378
rect -4886 16954 588810 17116
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15546 16954
rect 15782 16718 15866 16954
rect 16102 16718 35546 16954
rect 35782 16718 35866 16954
rect 36102 16718 55546 16954
rect 55782 16718 55866 16954
rect 56102 16718 75546 16954
rect 75782 16718 75866 16954
rect 76102 16718 95546 16954
rect 95782 16718 95866 16954
rect 96102 16718 115546 16954
rect 115782 16718 115866 16954
rect 116102 16718 135546 16954
rect 135782 16718 135866 16954
rect 136102 16718 155546 16954
rect 155782 16718 155866 16954
rect 156102 16718 175546 16954
rect 175782 16718 175866 16954
rect 176102 16718 195546 16954
rect 195782 16718 195866 16954
rect 196102 16718 215546 16954
rect 215782 16718 215866 16954
rect 216102 16718 235546 16954
rect 235782 16718 235866 16954
rect 236102 16718 255546 16954
rect 255782 16718 255866 16954
rect 256102 16718 275546 16954
rect 275782 16718 275866 16954
rect 276102 16718 295546 16954
rect 295782 16718 295866 16954
rect 296102 16718 315546 16954
rect 315782 16718 315866 16954
rect 316102 16718 335546 16954
rect 335782 16718 335866 16954
rect 336102 16718 355546 16954
rect 355782 16718 355866 16954
rect 356102 16718 375546 16954
rect 375782 16718 375866 16954
rect 376102 16718 395546 16954
rect 395782 16718 395866 16954
rect 396102 16718 415546 16954
rect 415782 16718 415866 16954
rect 416102 16718 435546 16954
rect 435782 16718 435866 16954
rect 436102 16718 455546 16954
rect 455782 16718 455866 16954
rect 456102 16718 475546 16954
rect 475782 16718 475866 16954
rect 476102 16718 495546 16954
rect 495782 16718 495866 16954
rect 496102 16718 515546 16954
rect 515782 16718 515866 16954
rect 516102 16718 535546 16954
rect 535782 16718 535866 16954
rect 536102 16718 555546 16954
rect 555782 16718 555866 16954
rect 556102 16718 575546 16954
rect 575782 16718 575866 16954
rect 576102 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect -4886 16556 588810 16718
rect -8726 14274 592650 14436
rect -8726 14038 -7734 14274
rect -7498 14038 -7414 14274
rect -7178 14038 12986 14274
rect 13222 14038 13306 14274
rect 13542 14038 32986 14274
rect 33222 14038 33306 14274
rect 33542 14038 52986 14274
rect 53222 14038 53306 14274
rect 53542 14038 72986 14274
rect 73222 14038 73306 14274
rect 73542 14038 92986 14274
rect 93222 14038 93306 14274
rect 93542 14038 112986 14274
rect 113222 14038 113306 14274
rect 113542 14038 132986 14274
rect 133222 14038 133306 14274
rect 133542 14038 152986 14274
rect 153222 14038 153306 14274
rect 153542 14038 172986 14274
rect 173222 14038 173306 14274
rect 173542 14038 192986 14274
rect 193222 14038 193306 14274
rect 193542 14038 212986 14274
rect 213222 14038 213306 14274
rect 213542 14038 232986 14274
rect 233222 14038 233306 14274
rect 233542 14038 252986 14274
rect 253222 14038 253306 14274
rect 253542 14038 272986 14274
rect 273222 14038 273306 14274
rect 273542 14038 292986 14274
rect 293222 14038 293306 14274
rect 293542 14038 312986 14274
rect 313222 14038 313306 14274
rect 313542 14038 332986 14274
rect 333222 14038 333306 14274
rect 333542 14038 352986 14274
rect 353222 14038 353306 14274
rect 353542 14038 372986 14274
rect 373222 14038 373306 14274
rect 373542 14038 392986 14274
rect 393222 14038 393306 14274
rect 393542 14038 412986 14274
rect 413222 14038 413306 14274
rect 413542 14038 432986 14274
rect 433222 14038 433306 14274
rect 433542 14038 452986 14274
rect 453222 14038 453306 14274
rect 453542 14038 472986 14274
rect 473222 14038 473306 14274
rect 473542 14038 492986 14274
rect 493222 14038 493306 14274
rect 493542 14038 512986 14274
rect 513222 14038 513306 14274
rect 513542 14038 532986 14274
rect 533222 14038 533306 14274
rect 533542 14038 552986 14274
rect 553222 14038 553306 14274
rect 553542 14038 572986 14274
rect 573222 14038 573306 14274
rect 573542 14038 591102 14274
rect 591338 14038 591422 14274
rect 591658 14038 592650 14274
rect -8726 13876 592650 14038
rect -2966 13294 586890 13456
rect -2966 13058 -2934 13294
rect -2698 13058 -2614 13294
rect -2378 13058 11826 13294
rect 12062 13058 12146 13294
rect 12382 13058 31826 13294
rect 32062 13058 32146 13294
rect 32382 13058 51826 13294
rect 52062 13058 52146 13294
rect 52382 13058 71826 13294
rect 72062 13058 72146 13294
rect 72382 13058 91826 13294
rect 92062 13058 92146 13294
rect 92382 13058 111826 13294
rect 112062 13058 112146 13294
rect 112382 13058 131826 13294
rect 132062 13058 132146 13294
rect 132382 13058 151826 13294
rect 152062 13058 152146 13294
rect 152382 13058 171826 13294
rect 172062 13058 172146 13294
rect 172382 13058 191826 13294
rect 192062 13058 192146 13294
rect 192382 13058 211826 13294
rect 212062 13058 212146 13294
rect 212382 13058 231826 13294
rect 232062 13058 232146 13294
rect 232382 13058 251826 13294
rect 252062 13058 252146 13294
rect 252382 13058 271826 13294
rect 272062 13058 272146 13294
rect 272382 13058 291826 13294
rect 292062 13058 292146 13294
rect 292382 13058 311826 13294
rect 312062 13058 312146 13294
rect 312382 13058 331826 13294
rect 332062 13058 332146 13294
rect 332382 13058 351826 13294
rect 352062 13058 352146 13294
rect 352382 13058 371826 13294
rect 372062 13058 372146 13294
rect 372382 13058 391826 13294
rect 392062 13058 392146 13294
rect 392382 13058 411826 13294
rect 412062 13058 412146 13294
rect 412382 13058 431826 13294
rect 432062 13058 432146 13294
rect 432382 13058 451826 13294
rect 452062 13058 452146 13294
rect 452382 13058 471826 13294
rect 472062 13058 472146 13294
rect 472382 13058 491826 13294
rect 492062 13058 492146 13294
rect 492382 13058 511826 13294
rect 512062 13058 512146 13294
rect 512382 13058 531826 13294
rect 532062 13058 532146 13294
rect 532382 13058 551826 13294
rect 552062 13058 552146 13294
rect 552382 13058 571826 13294
rect 572062 13058 572146 13294
rect 572382 13058 586302 13294
rect 586538 13058 586622 13294
rect 586858 13058 586890 13294
rect -2966 12896 586890 13058
rect -6806 10614 590730 10776
rect -6806 10378 -5814 10614
rect -5578 10378 -5494 10614
rect -5258 10378 9266 10614
rect 9502 10378 9586 10614
rect 9822 10378 29266 10614
rect 29502 10378 29586 10614
rect 29822 10378 49266 10614
rect 49502 10378 49586 10614
rect 49822 10378 69266 10614
rect 69502 10378 69586 10614
rect 69822 10378 89266 10614
rect 89502 10378 89586 10614
rect 89822 10378 109266 10614
rect 109502 10378 109586 10614
rect 109822 10378 129266 10614
rect 129502 10378 129586 10614
rect 129822 10378 149266 10614
rect 149502 10378 149586 10614
rect 149822 10378 169266 10614
rect 169502 10378 169586 10614
rect 169822 10378 189266 10614
rect 189502 10378 189586 10614
rect 189822 10378 209266 10614
rect 209502 10378 209586 10614
rect 209822 10378 229266 10614
rect 229502 10378 229586 10614
rect 229822 10378 249266 10614
rect 249502 10378 249586 10614
rect 249822 10378 269266 10614
rect 269502 10378 269586 10614
rect 269822 10378 289266 10614
rect 289502 10378 289586 10614
rect 289822 10378 309266 10614
rect 309502 10378 309586 10614
rect 309822 10378 329266 10614
rect 329502 10378 329586 10614
rect 329822 10378 349266 10614
rect 349502 10378 349586 10614
rect 349822 10378 369266 10614
rect 369502 10378 369586 10614
rect 369822 10378 389266 10614
rect 389502 10378 389586 10614
rect 389822 10378 409266 10614
rect 409502 10378 409586 10614
rect 409822 10378 429266 10614
rect 429502 10378 429586 10614
rect 429822 10378 449266 10614
rect 449502 10378 449586 10614
rect 449822 10378 469266 10614
rect 469502 10378 469586 10614
rect 469822 10378 489266 10614
rect 489502 10378 489586 10614
rect 489822 10378 509266 10614
rect 509502 10378 509586 10614
rect 509822 10378 529266 10614
rect 529502 10378 529586 10614
rect 529822 10378 549266 10614
rect 549502 10378 549586 10614
rect 549822 10378 569266 10614
rect 569502 10378 569586 10614
rect 569822 10378 589182 10614
rect 589418 10378 589502 10614
rect 589738 10378 590730 10614
rect -6806 10216 590730 10378
rect -4886 6954 588810 7116
rect -4886 6718 -3894 6954
rect -3658 6718 -3574 6954
rect -3338 6718 5546 6954
rect 5782 6718 5866 6954
rect 6102 6718 25546 6954
rect 25782 6718 25866 6954
rect 26102 6718 45546 6954
rect 45782 6718 45866 6954
rect 46102 6718 65546 6954
rect 65782 6718 65866 6954
rect 66102 6718 85546 6954
rect 85782 6718 85866 6954
rect 86102 6718 105546 6954
rect 105782 6718 105866 6954
rect 106102 6718 125546 6954
rect 125782 6718 125866 6954
rect 126102 6718 145546 6954
rect 145782 6718 145866 6954
rect 146102 6718 165546 6954
rect 165782 6718 165866 6954
rect 166102 6718 185546 6954
rect 185782 6718 185866 6954
rect 186102 6718 205546 6954
rect 205782 6718 205866 6954
rect 206102 6718 225546 6954
rect 225782 6718 225866 6954
rect 226102 6718 245546 6954
rect 245782 6718 245866 6954
rect 246102 6718 265546 6954
rect 265782 6718 265866 6954
rect 266102 6718 285546 6954
rect 285782 6718 285866 6954
rect 286102 6718 305546 6954
rect 305782 6718 305866 6954
rect 306102 6718 325546 6954
rect 325782 6718 325866 6954
rect 326102 6718 345546 6954
rect 345782 6718 345866 6954
rect 346102 6718 365546 6954
rect 365782 6718 365866 6954
rect 366102 6718 385546 6954
rect 385782 6718 385866 6954
rect 386102 6718 405546 6954
rect 405782 6718 405866 6954
rect 406102 6718 425546 6954
rect 425782 6718 425866 6954
rect 426102 6718 445546 6954
rect 445782 6718 445866 6954
rect 446102 6718 465546 6954
rect 465782 6718 465866 6954
rect 466102 6718 485546 6954
rect 485782 6718 485866 6954
rect 486102 6718 505546 6954
rect 505782 6718 505866 6954
rect 506102 6718 525546 6954
rect 525782 6718 525866 6954
rect 526102 6718 545546 6954
rect 545782 6718 545866 6954
rect 546102 6718 565546 6954
rect 565782 6718 565866 6954
rect 566102 6718 587262 6954
rect 587498 6718 587582 6954
rect 587818 6718 588810 6954
rect -4886 6556 588810 6718
rect -2966 3294 586890 3456
rect -2966 3058 -1974 3294
rect -1738 3058 -1654 3294
rect -1418 3058 1826 3294
rect 2062 3058 2146 3294
rect 2382 3058 21826 3294
rect 22062 3058 22146 3294
rect 22382 3058 41826 3294
rect 42062 3058 42146 3294
rect 42382 3058 61826 3294
rect 62062 3058 62146 3294
rect 62382 3058 81826 3294
rect 82062 3058 82146 3294
rect 82382 3058 101826 3294
rect 102062 3058 102146 3294
rect 102382 3058 121826 3294
rect 122062 3058 122146 3294
rect 122382 3058 141826 3294
rect 142062 3058 142146 3294
rect 142382 3058 161826 3294
rect 162062 3058 162146 3294
rect 162382 3058 181826 3294
rect 182062 3058 182146 3294
rect 182382 3058 201826 3294
rect 202062 3058 202146 3294
rect 202382 3058 221826 3294
rect 222062 3058 222146 3294
rect 222382 3058 241826 3294
rect 242062 3058 242146 3294
rect 242382 3058 261826 3294
rect 262062 3058 262146 3294
rect 262382 3058 281826 3294
rect 282062 3058 282146 3294
rect 282382 3058 301826 3294
rect 302062 3058 302146 3294
rect 302382 3058 321826 3294
rect 322062 3058 322146 3294
rect 322382 3058 341826 3294
rect 342062 3058 342146 3294
rect 342382 3058 361826 3294
rect 362062 3058 362146 3294
rect 362382 3058 381826 3294
rect 382062 3058 382146 3294
rect 382382 3058 401826 3294
rect 402062 3058 402146 3294
rect 402382 3058 421826 3294
rect 422062 3058 422146 3294
rect 422382 3058 441826 3294
rect 442062 3058 442146 3294
rect 442382 3058 461826 3294
rect 462062 3058 462146 3294
rect 462382 3058 481826 3294
rect 482062 3058 482146 3294
rect 482382 3058 501826 3294
rect 502062 3058 502146 3294
rect 502382 3058 521826 3294
rect 522062 3058 522146 3294
rect 522382 3058 541826 3294
rect 542062 3058 542146 3294
rect 542382 3058 561826 3294
rect 562062 3058 562146 3294
rect 562382 3058 581826 3294
rect 582062 3058 582146 3294
rect 582382 3058 585342 3294
rect 585578 3058 585662 3294
rect 585898 3058 586890 3294
rect -2966 2896 586890 3058
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 21826 -346
rect 22062 -582 22146 -346
rect 22382 -582 41826 -346
rect 42062 -582 42146 -346
rect 42382 -582 61826 -346
rect 62062 -582 62146 -346
rect 62382 -582 81826 -346
rect 82062 -582 82146 -346
rect 82382 -582 101826 -346
rect 102062 -582 102146 -346
rect 102382 -582 121826 -346
rect 122062 -582 122146 -346
rect 122382 -582 141826 -346
rect 142062 -582 142146 -346
rect 142382 -582 161826 -346
rect 162062 -582 162146 -346
rect 162382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 201826 -346
rect 202062 -582 202146 -346
rect 202382 -582 221826 -346
rect 222062 -582 222146 -346
rect 222382 -582 241826 -346
rect 242062 -582 242146 -346
rect 242382 -582 261826 -346
rect 262062 -582 262146 -346
rect 262382 -582 281826 -346
rect 282062 -582 282146 -346
rect 282382 -582 301826 -346
rect 302062 -582 302146 -346
rect 302382 -582 321826 -346
rect 322062 -582 322146 -346
rect 322382 -582 341826 -346
rect 342062 -582 342146 -346
rect 342382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 381826 -346
rect 382062 -582 382146 -346
rect 382382 -582 401826 -346
rect 402062 -582 402146 -346
rect 402382 -582 421826 -346
rect 422062 -582 422146 -346
rect 422382 -582 441826 -346
rect 442062 -582 442146 -346
rect 442382 -582 461826 -346
rect 462062 -582 462146 -346
rect 462382 -582 481826 -346
rect 482062 -582 482146 -346
rect 482382 -582 501826 -346
rect 502062 -582 502146 -346
rect 502382 -582 521826 -346
rect 522062 -582 522146 -346
rect 522382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 561826 -346
rect 562062 -582 562146 -346
rect 562382 -582 581826 -346
rect 582062 -582 582146 -346
rect 582382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 21826 -666
rect 22062 -902 22146 -666
rect 22382 -902 41826 -666
rect 42062 -902 42146 -666
rect 42382 -902 61826 -666
rect 62062 -902 62146 -666
rect 62382 -902 81826 -666
rect 82062 -902 82146 -666
rect 82382 -902 101826 -666
rect 102062 -902 102146 -666
rect 102382 -902 121826 -666
rect 122062 -902 122146 -666
rect 122382 -902 141826 -666
rect 142062 -902 142146 -666
rect 142382 -902 161826 -666
rect 162062 -902 162146 -666
rect 162382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 201826 -666
rect 202062 -902 202146 -666
rect 202382 -902 221826 -666
rect 222062 -902 222146 -666
rect 222382 -902 241826 -666
rect 242062 -902 242146 -666
rect 242382 -902 261826 -666
rect 262062 -902 262146 -666
rect 262382 -902 281826 -666
rect 282062 -902 282146 -666
rect 282382 -902 301826 -666
rect 302062 -902 302146 -666
rect 302382 -902 321826 -666
rect 322062 -902 322146 -666
rect 322382 -902 341826 -666
rect 342062 -902 342146 -666
rect 342382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 381826 -666
rect 382062 -902 382146 -666
rect 382382 -902 401826 -666
rect 402062 -902 402146 -666
rect 402382 -902 421826 -666
rect 422062 -902 422146 -666
rect 422382 -902 441826 -666
rect 442062 -902 442146 -666
rect 442382 -902 461826 -666
rect 462062 -902 462146 -666
rect 462382 -902 481826 -666
rect 482062 -902 482146 -666
rect 482382 -902 501826 -666
rect 502062 -902 502146 -666
rect 502382 -902 521826 -666
rect 522062 -902 522146 -666
rect 522382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 561826 -666
rect 562062 -902 562146 -666
rect 562382 -902 581826 -666
rect 582062 -902 582146 -666
rect 582382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 11826 -1306
rect 12062 -1542 12146 -1306
rect 12382 -1542 31826 -1306
rect 32062 -1542 32146 -1306
rect 32382 -1542 51826 -1306
rect 52062 -1542 52146 -1306
rect 52382 -1542 71826 -1306
rect 72062 -1542 72146 -1306
rect 72382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 111826 -1306
rect 112062 -1542 112146 -1306
rect 112382 -1542 131826 -1306
rect 132062 -1542 132146 -1306
rect 132382 -1542 151826 -1306
rect 152062 -1542 152146 -1306
rect 152382 -1542 171826 -1306
rect 172062 -1542 172146 -1306
rect 172382 -1542 191826 -1306
rect 192062 -1542 192146 -1306
rect 192382 -1542 211826 -1306
rect 212062 -1542 212146 -1306
rect 212382 -1542 231826 -1306
rect 232062 -1542 232146 -1306
rect 232382 -1542 251826 -1306
rect 252062 -1542 252146 -1306
rect 252382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 291826 -1306
rect 292062 -1542 292146 -1306
rect 292382 -1542 311826 -1306
rect 312062 -1542 312146 -1306
rect 312382 -1542 331826 -1306
rect 332062 -1542 332146 -1306
rect 332382 -1542 351826 -1306
rect 352062 -1542 352146 -1306
rect 352382 -1542 371826 -1306
rect 372062 -1542 372146 -1306
rect 372382 -1542 391826 -1306
rect 392062 -1542 392146 -1306
rect 392382 -1542 411826 -1306
rect 412062 -1542 412146 -1306
rect 412382 -1542 431826 -1306
rect 432062 -1542 432146 -1306
rect 432382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 471826 -1306
rect 472062 -1542 472146 -1306
rect 472382 -1542 491826 -1306
rect 492062 -1542 492146 -1306
rect 492382 -1542 511826 -1306
rect 512062 -1542 512146 -1306
rect 512382 -1542 531826 -1306
rect 532062 -1542 532146 -1306
rect 532382 -1542 551826 -1306
rect 552062 -1542 552146 -1306
rect 552382 -1542 571826 -1306
rect 572062 -1542 572146 -1306
rect 572382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 11826 -1626
rect 12062 -1862 12146 -1626
rect 12382 -1862 31826 -1626
rect 32062 -1862 32146 -1626
rect 32382 -1862 51826 -1626
rect 52062 -1862 52146 -1626
rect 52382 -1862 71826 -1626
rect 72062 -1862 72146 -1626
rect 72382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 111826 -1626
rect 112062 -1862 112146 -1626
rect 112382 -1862 131826 -1626
rect 132062 -1862 132146 -1626
rect 132382 -1862 151826 -1626
rect 152062 -1862 152146 -1626
rect 152382 -1862 171826 -1626
rect 172062 -1862 172146 -1626
rect 172382 -1862 191826 -1626
rect 192062 -1862 192146 -1626
rect 192382 -1862 211826 -1626
rect 212062 -1862 212146 -1626
rect 212382 -1862 231826 -1626
rect 232062 -1862 232146 -1626
rect 232382 -1862 251826 -1626
rect 252062 -1862 252146 -1626
rect 252382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 291826 -1626
rect 292062 -1862 292146 -1626
rect 292382 -1862 311826 -1626
rect 312062 -1862 312146 -1626
rect 312382 -1862 331826 -1626
rect 332062 -1862 332146 -1626
rect 332382 -1862 351826 -1626
rect 352062 -1862 352146 -1626
rect 352382 -1862 371826 -1626
rect 372062 -1862 372146 -1626
rect 372382 -1862 391826 -1626
rect 392062 -1862 392146 -1626
rect 392382 -1862 411826 -1626
rect 412062 -1862 412146 -1626
rect 412382 -1862 431826 -1626
rect 432062 -1862 432146 -1626
rect 432382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 471826 -1626
rect 472062 -1862 472146 -1626
rect 472382 -1862 491826 -1626
rect 492062 -1862 492146 -1626
rect 492382 -1862 511826 -1626
rect 512062 -1862 512146 -1626
rect 512382 -1862 531826 -1626
rect 532062 -1862 532146 -1626
rect 532382 -1862 551826 -1626
rect 552062 -1862 552146 -1626
rect 552382 -1862 571826 -1626
rect 572062 -1862 572146 -1626
rect 572382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 25546 -2266
rect 25782 -2502 25866 -2266
rect 26102 -2502 45546 -2266
rect 45782 -2502 45866 -2266
rect 46102 -2502 65546 -2266
rect 65782 -2502 65866 -2266
rect 66102 -2502 85546 -2266
rect 85782 -2502 85866 -2266
rect 86102 -2502 105546 -2266
rect 105782 -2502 105866 -2266
rect 106102 -2502 125546 -2266
rect 125782 -2502 125866 -2266
rect 126102 -2502 145546 -2266
rect 145782 -2502 145866 -2266
rect 146102 -2502 165546 -2266
rect 165782 -2502 165866 -2266
rect 166102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 205546 -2266
rect 205782 -2502 205866 -2266
rect 206102 -2502 225546 -2266
rect 225782 -2502 225866 -2266
rect 226102 -2502 245546 -2266
rect 245782 -2502 245866 -2266
rect 246102 -2502 265546 -2266
rect 265782 -2502 265866 -2266
rect 266102 -2502 285546 -2266
rect 285782 -2502 285866 -2266
rect 286102 -2502 305546 -2266
rect 305782 -2502 305866 -2266
rect 306102 -2502 325546 -2266
rect 325782 -2502 325866 -2266
rect 326102 -2502 345546 -2266
rect 345782 -2502 345866 -2266
rect 346102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 385546 -2266
rect 385782 -2502 385866 -2266
rect 386102 -2502 405546 -2266
rect 405782 -2502 405866 -2266
rect 406102 -2502 425546 -2266
rect 425782 -2502 425866 -2266
rect 426102 -2502 445546 -2266
rect 445782 -2502 445866 -2266
rect 446102 -2502 465546 -2266
rect 465782 -2502 465866 -2266
rect 466102 -2502 485546 -2266
rect 485782 -2502 485866 -2266
rect 486102 -2502 505546 -2266
rect 505782 -2502 505866 -2266
rect 506102 -2502 525546 -2266
rect 525782 -2502 525866 -2266
rect 526102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 565546 -2266
rect 565782 -2502 565866 -2266
rect 566102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 25546 -2586
rect 25782 -2822 25866 -2586
rect 26102 -2822 45546 -2586
rect 45782 -2822 45866 -2586
rect 46102 -2822 65546 -2586
rect 65782 -2822 65866 -2586
rect 66102 -2822 85546 -2586
rect 85782 -2822 85866 -2586
rect 86102 -2822 105546 -2586
rect 105782 -2822 105866 -2586
rect 106102 -2822 125546 -2586
rect 125782 -2822 125866 -2586
rect 126102 -2822 145546 -2586
rect 145782 -2822 145866 -2586
rect 146102 -2822 165546 -2586
rect 165782 -2822 165866 -2586
rect 166102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 205546 -2586
rect 205782 -2822 205866 -2586
rect 206102 -2822 225546 -2586
rect 225782 -2822 225866 -2586
rect 226102 -2822 245546 -2586
rect 245782 -2822 245866 -2586
rect 246102 -2822 265546 -2586
rect 265782 -2822 265866 -2586
rect 266102 -2822 285546 -2586
rect 285782 -2822 285866 -2586
rect 286102 -2822 305546 -2586
rect 305782 -2822 305866 -2586
rect 306102 -2822 325546 -2586
rect 325782 -2822 325866 -2586
rect 326102 -2822 345546 -2586
rect 345782 -2822 345866 -2586
rect 346102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 385546 -2586
rect 385782 -2822 385866 -2586
rect 386102 -2822 405546 -2586
rect 405782 -2822 405866 -2586
rect 406102 -2822 425546 -2586
rect 425782 -2822 425866 -2586
rect 426102 -2822 445546 -2586
rect 445782 -2822 445866 -2586
rect 446102 -2822 465546 -2586
rect 465782 -2822 465866 -2586
rect 466102 -2822 485546 -2586
rect 485782 -2822 485866 -2586
rect 486102 -2822 505546 -2586
rect 505782 -2822 505866 -2586
rect 506102 -2822 525546 -2586
rect 525782 -2822 525866 -2586
rect 526102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 565546 -2586
rect 565782 -2822 565866 -2586
rect 566102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15546 -3226
rect 15782 -3462 15866 -3226
rect 16102 -3462 35546 -3226
rect 35782 -3462 35866 -3226
rect 36102 -3462 55546 -3226
rect 55782 -3462 55866 -3226
rect 56102 -3462 75546 -3226
rect 75782 -3462 75866 -3226
rect 76102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 115546 -3226
rect 115782 -3462 115866 -3226
rect 116102 -3462 135546 -3226
rect 135782 -3462 135866 -3226
rect 136102 -3462 155546 -3226
rect 155782 -3462 155866 -3226
rect 156102 -3462 175546 -3226
rect 175782 -3462 175866 -3226
rect 176102 -3462 195546 -3226
rect 195782 -3462 195866 -3226
rect 196102 -3462 215546 -3226
rect 215782 -3462 215866 -3226
rect 216102 -3462 235546 -3226
rect 235782 -3462 235866 -3226
rect 236102 -3462 255546 -3226
rect 255782 -3462 255866 -3226
rect 256102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 295546 -3226
rect 295782 -3462 295866 -3226
rect 296102 -3462 315546 -3226
rect 315782 -3462 315866 -3226
rect 316102 -3462 335546 -3226
rect 335782 -3462 335866 -3226
rect 336102 -3462 355546 -3226
rect 355782 -3462 355866 -3226
rect 356102 -3462 375546 -3226
rect 375782 -3462 375866 -3226
rect 376102 -3462 395546 -3226
rect 395782 -3462 395866 -3226
rect 396102 -3462 415546 -3226
rect 415782 -3462 415866 -3226
rect 416102 -3462 435546 -3226
rect 435782 -3462 435866 -3226
rect 436102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 475546 -3226
rect 475782 -3462 475866 -3226
rect 476102 -3462 495546 -3226
rect 495782 -3462 495866 -3226
rect 496102 -3462 515546 -3226
rect 515782 -3462 515866 -3226
rect 516102 -3462 535546 -3226
rect 535782 -3462 535866 -3226
rect 536102 -3462 555546 -3226
rect 555782 -3462 555866 -3226
rect 556102 -3462 575546 -3226
rect 575782 -3462 575866 -3226
rect 576102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15546 -3546
rect 15782 -3782 15866 -3546
rect 16102 -3782 35546 -3546
rect 35782 -3782 35866 -3546
rect 36102 -3782 55546 -3546
rect 55782 -3782 55866 -3546
rect 56102 -3782 75546 -3546
rect 75782 -3782 75866 -3546
rect 76102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 115546 -3546
rect 115782 -3782 115866 -3546
rect 116102 -3782 135546 -3546
rect 135782 -3782 135866 -3546
rect 136102 -3782 155546 -3546
rect 155782 -3782 155866 -3546
rect 156102 -3782 175546 -3546
rect 175782 -3782 175866 -3546
rect 176102 -3782 195546 -3546
rect 195782 -3782 195866 -3546
rect 196102 -3782 215546 -3546
rect 215782 -3782 215866 -3546
rect 216102 -3782 235546 -3546
rect 235782 -3782 235866 -3546
rect 236102 -3782 255546 -3546
rect 255782 -3782 255866 -3546
rect 256102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 295546 -3546
rect 295782 -3782 295866 -3546
rect 296102 -3782 315546 -3546
rect 315782 -3782 315866 -3546
rect 316102 -3782 335546 -3546
rect 335782 -3782 335866 -3546
rect 336102 -3782 355546 -3546
rect 355782 -3782 355866 -3546
rect 356102 -3782 375546 -3546
rect 375782 -3782 375866 -3546
rect 376102 -3782 395546 -3546
rect 395782 -3782 395866 -3546
rect 396102 -3782 415546 -3546
rect 415782 -3782 415866 -3546
rect 416102 -3782 435546 -3546
rect 435782 -3782 435866 -3546
rect 436102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 475546 -3546
rect 475782 -3782 475866 -3546
rect 476102 -3782 495546 -3546
rect 495782 -3782 495866 -3546
rect 496102 -3782 515546 -3546
rect 515782 -3782 515866 -3546
rect 516102 -3782 535546 -3546
rect 535782 -3782 535866 -3546
rect 536102 -3782 555546 -3546
rect 555782 -3782 555866 -3546
rect 556102 -3782 575546 -3546
rect 575782 -3782 575866 -3546
rect 576102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 29266 -4186
rect 29502 -4422 29586 -4186
rect 29822 -4422 49266 -4186
rect 49502 -4422 49586 -4186
rect 49822 -4422 69266 -4186
rect 69502 -4422 69586 -4186
rect 69822 -4422 89266 -4186
rect 89502 -4422 89586 -4186
rect 89822 -4422 109266 -4186
rect 109502 -4422 109586 -4186
rect 109822 -4422 129266 -4186
rect 129502 -4422 129586 -4186
rect 129822 -4422 149266 -4186
rect 149502 -4422 149586 -4186
rect 149822 -4422 169266 -4186
rect 169502 -4422 169586 -4186
rect 169822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 209266 -4186
rect 209502 -4422 209586 -4186
rect 209822 -4422 229266 -4186
rect 229502 -4422 229586 -4186
rect 229822 -4422 249266 -4186
rect 249502 -4422 249586 -4186
rect 249822 -4422 269266 -4186
rect 269502 -4422 269586 -4186
rect 269822 -4422 289266 -4186
rect 289502 -4422 289586 -4186
rect 289822 -4422 309266 -4186
rect 309502 -4422 309586 -4186
rect 309822 -4422 329266 -4186
rect 329502 -4422 329586 -4186
rect 329822 -4422 349266 -4186
rect 349502 -4422 349586 -4186
rect 349822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 389266 -4186
rect 389502 -4422 389586 -4186
rect 389822 -4422 409266 -4186
rect 409502 -4422 409586 -4186
rect 409822 -4422 429266 -4186
rect 429502 -4422 429586 -4186
rect 429822 -4422 449266 -4186
rect 449502 -4422 449586 -4186
rect 449822 -4422 469266 -4186
rect 469502 -4422 469586 -4186
rect 469822 -4422 489266 -4186
rect 489502 -4422 489586 -4186
rect 489822 -4422 509266 -4186
rect 509502 -4422 509586 -4186
rect 509822 -4422 529266 -4186
rect 529502 -4422 529586 -4186
rect 529822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 569266 -4186
rect 569502 -4422 569586 -4186
rect 569822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 29266 -4506
rect 29502 -4742 29586 -4506
rect 29822 -4742 49266 -4506
rect 49502 -4742 49586 -4506
rect 49822 -4742 69266 -4506
rect 69502 -4742 69586 -4506
rect 69822 -4742 89266 -4506
rect 89502 -4742 89586 -4506
rect 89822 -4742 109266 -4506
rect 109502 -4742 109586 -4506
rect 109822 -4742 129266 -4506
rect 129502 -4742 129586 -4506
rect 129822 -4742 149266 -4506
rect 149502 -4742 149586 -4506
rect 149822 -4742 169266 -4506
rect 169502 -4742 169586 -4506
rect 169822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 209266 -4506
rect 209502 -4742 209586 -4506
rect 209822 -4742 229266 -4506
rect 229502 -4742 229586 -4506
rect 229822 -4742 249266 -4506
rect 249502 -4742 249586 -4506
rect 249822 -4742 269266 -4506
rect 269502 -4742 269586 -4506
rect 269822 -4742 289266 -4506
rect 289502 -4742 289586 -4506
rect 289822 -4742 309266 -4506
rect 309502 -4742 309586 -4506
rect 309822 -4742 329266 -4506
rect 329502 -4742 329586 -4506
rect 329822 -4742 349266 -4506
rect 349502 -4742 349586 -4506
rect 349822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 389266 -4506
rect 389502 -4742 389586 -4506
rect 389822 -4742 409266 -4506
rect 409502 -4742 409586 -4506
rect 409822 -4742 429266 -4506
rect 429502 -4742 429586 -4506
rect 429822 -4742 449266 -4506
rect 449502 -4742 449586 -4506
rect 449822 -4742 469266 -4506
rect 469502 -4742 469586 -4506
rect 469822 -4742 489266 -4506
rect 489502 -4742 489586 -4506
rect 489822 -4742 509266 -4506
rect 509502 -4742 509586 -4506
rect 509822 -4742 529266 -4506
rect 529502 -4742 529586 -4506
rect 529822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 569266 -4506
rect 569502 -4742 569586 -4506
rect 569822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 19266 -5146
rect 19502 -5382 19586 -5146
rect 19822 -5382 39266 -5146
rect 39502 -5382 39586 -5146
rect 39822 -5382 59266 -5146
rect 59502 -5382 59586 -5146
rect 59822 -5382 79266 -5146
rect 79502 -5382 79586 -5146
rect 79822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 119266 -5146
rect 119502 -5382 119586 -5146
rect 119822 -5382 139266 -5146
rect 139502 -5382 139586 -5146
rect 139822 -5382 159266 -5146
rect 159502 -5382 159586 -5146
rect 159822 -5382 179266 -5146
rect 179502 -5382 179586 -5146
rect 179822 -5382 199266 -5146
rect 199502 -5382 199586 -5146
rect 199822 -5382 219266 -5146
rect 219502 -5382 219586 -5146
rect 219822 -5382 239266 -5146
rect 239502 -5382 239586 -5146
rect 239822 -5382 259266 -5146
rect 259502 -5382 259586 -5146
rect 259822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 299266 -5146
rect 299502 -5382 299586 -5146
rect 299822 -5382 319266 -5146
rect 319502 -5382 319586 -5146
rect 319822 -5382 339266 -5146
rect 339502 -5382 339586 -5146
rect 339822 -5382 359266 -5146
rect 359502 -5382 359586 -5146
rect 359822 -5382 379266 -5146
rect 379502 -5382 379586 -5146
rect 379822 -5382 399266 -5146
rect 399502 -5382 399586 -5146
rect 399822 -5382 419266 -5146
rect 419502 -5382 419586 -5146
rect 419822 -5382 439266 -5146
rect 439502 -5382 439586 -5146
rect 439822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 479266 -5146
rect 479502 -5382 479586 -5146
rect 479822 -5382 499266 -5146
rect 499502 -5382 499586 -5146
rect 499822 -5382 519266 -5146
rect 519502 -5382 519586 -5146
rect 519822 -5382 539266 -5146
rect 539502 -5382 539586 -5146
rect 539822 -5382 559266 -5146
rect 559502 -5382 559586 -5146
rect 559822 -5382 579266 -5146
rect 579502 -5382 579586 -5146
rect 579822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 19266 -5466
rect 19502 -5702 19586 -5466
rect 19822 -5702 39266 -5466
rect 39502 -5702 39586 -5466
rect 39822 -5702 59266 -5466
rect 59502 -5702 59586 -5466
rect 59822 -5702 79266 -5466
rect 79502 -5702 79586 -5466
rect 79822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 119266 -5466
rect 119502 -5702 119586 -5466
rect 119822 -5702 139266 -5466
rect 139502 -5702 139586 -5466
rect 139822 -5702 159266 -5466
rect 159502 -5702 159586 -5466
rect 159822 -5702 179266 -5466
rect 179502 -5702 179586 -5466
rect 179822 -5702 199266 -5466
rect 199502 -5702 199586 -5466
rect 199822 -5702 219266 -5466
rect 219502 -5702 219586 -5466
rect 219822 -5702 239266 -5466
rect 239502 -5702 239586 -5466
rect 239822 -5702 259266 -5466
rect 259502 -5702 259586 -5466
rect 259822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 299266 -5466
rect 299502 -5702 299586 -5466
rect 299822 -5702 319266 -5466
rect 319502 -5702 319586 -5466
rect 319822 -5702 339266 -5466
rect 339502 -5702 339586 -5466
rect 339822 -5702 359266 -5466
rect 359502 -5702 359586 -5466
rect 359822 -5702 379266 -5466
rect 379502 -5702 379586 -5466
rect 379822 -5702 399266 -5466
rect 399502 -5702 399586 -5466
rect 399822 -5702 419266 -5466
rect 419502 -5702 419586 -5466
rect 419822 -5702 439266 -5466
rect 439502 -5702 439586 -5466
rect 439822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 479266 -5466
rect 479502 -5702 479586 -5466
rect 479822 -5702 499266 -5466
rect 499502 -5702 499586 -5466
rect 499822 -5702 519266 -5466
rect 519502 -5702 519586 -5466
rect 519822 -5702 539266 -5466
rect 539502 -5702 539586 -5466
rect 539822 -5702 559266 -5466
rect 559502 -5702 559586 -5466
rect 559822 -5702 579266 -5466
rect 579502 -5702 579586 -5466
rect 579822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 32986 -6106
rect 33222 -6342 33306 -6106
rect 33542 -6342 52986 -6106
rect 53222 -6342 53306 -6106
rect 53542 -6342 72986 -6106
rect 73222 -6342 73306 -6106
rect 73542 -6342 92986 -6106
rect 93222 -6342 93306 -6106
rect 93542 -6342 112986 -6106
rect 113222 -6342 113306 -6106
rect 113542 -6342 132986 -6106
rect 133222 -6342 133306 -6106
rect 133542 -6342 152986 -6106
rect 153222 -6342 153306 -6106
rect 153542 -6342 172986 -6106
rect 173222 -6342 173306 -6106
rect 173542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 212986 -6106
rect 213222 -6342 213306 -6106
rect 213542 -6342 232986 -6106
rect 233222 -6342 233306 -6106
rect 233542 -6342 252986 -6106
rect 253222 -6342 253306 -6106
rect 253542 -6342 272986 -6106
rect 273222 -6342 273306 -6106
rect 273542 -6342 292986 -6106
rect 293222 -6342 293306 -6106
rect 293542 -6342 312986 -6106
rect 313222 -6342 313306 -6106
rect 313542 -6342 332986 -6106
rect 333222 -6342 333306 -6106
rect 333542 -6342 352986 -6106
rect 353222 -6342 353306 -6106
rect 353542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 392986 -6106
rect 393222 -6342 393306 -6106
rect 393542 -6342 412986 -6106
rect 413222 -6342 413306 -6106
rect 413542 -6342 432986 -6106
rect 433222 -6342 433306 -6106
rect 433542 -6342 452986 -6106
rect 453222 -6342 453306 -6106
rect 453542 -6342 472986 -6106
rect 473222 -6342 473306 -6106
rect 473542 -6342 492986 -6106
rect 493222 -6342 493306 -6106
rect 493542 -6342 512986 -6106
rect 513222 -6342 513306 -6106
rect 513542 -6342 532986 -6106
rect 533222 -6342 533306 -6106
rect 533542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 572986 -6106
rect 573222 -6342 573306 -6106
rect 573542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 32986 -6426
rect 33222 -6662 33306 -6426
rect 33542 -6662 52986 -6426
rect 53222 -6662 53306 -6426
rect 53542 -6662 72986 -6426
rect 73222 -6662 73306 -6426
rect 73542 -6662 92986 -6426
rect 93222 -6662 93306 -6426
rect 93542 -6662 112986 -6426
rect 113222 -6662 113306 -6426
rect 113542 -6662 132986 -6426
rect 133222 -6662 133306 -6426
rect 133542 -6662 152986 -6426
rect 153222 -6662 153306 -6426
rect 153542 -6662 172986 -6426
rect 173222 -6662 173306 -6426
rect 173542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 212986 -6426
rect 213222 -6662 213306 -6426
rect 213542 -6662 232986 -6426
rect 233222 -6662 233306 -6426
rect 233542 -6662 252986 -6426
rect 253222 -6662 253306 -6426
rect 253542 -6662 272986 -6426
rect 273222 -6662 273306 -6426
rect 273542 -6662 292986 -6426
rect 293222 -6662 293306 -6426
rect 293542 -6662 312986 -6426
rect 313222 -6662 313306 -6426
rect 313542 -6662 332986 -6426
rect 333222 -6662 333306 -6426
rect 333542 -6662 352986 -6426
rect 353222 -6662 353306 -6426
rect 353542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 392986 -6426
rect 393222 -6662 393306 -6426
rect 393542 -6662 412986 -6426
rect 413222 -6662 413306 -6426
rect 413542 -6662 432986 -6426
rect 433222 -6662 433306 -6426
rect 433542 -6662 452986 -6426
rect 453222 -6662 453306 -6426
rect 453542 -6662 472986 -6426
rect 473222 -6662 473306 -6426
rect 473542 -6662 492986 -6426
rect 493222 -6662 493306 -6426
rect 493542 -6662 512986 -6426
rect 513222 -6662 513306 -6426
rect 513542 -6662 532986 -6426
rect 533222 -6662 533306 -6426
rect 533542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 572986 -6426
rect 573222 -6662 573306 -6426
rect 573542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 22986 -7066
rect 23222 -7302 23306 -7066
rect 23542 -7302 42986 -7066
rect 43222 -7302 43306 -7066
rect 43542 -7302 62986 -7066
rect 63222 -7302 63306 -7066
rect 63542 -7302 82986 -7066
rect 83222 -7302 83306 -7066
rect 83542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 122986 -7066
rect 123222 -7302 123306 -7066
rect 123542 -7302 142986 -7066
rect 143222 -7302 143306 -7066
rect 143542 -7302 162986 -7066
rect 163222 -7302 163306 -7066
rect 163542 -7302 182986 -7066
rect 183222 -7302 183306 -7066
rect 183542 -7302 202986 -7066
rect 203222 -7302 203306 -7066
rect 203542 -7302 222986 -7066
rect 223222 -7302 223306 -7066
rect 223542 -7302 242986 -7066
rect 243222 -7302 243306 -7066
rect 243542 -7302 262986 -7066
rect 263222 -7302 263306 -7066
rect 263542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 302986 -7066
rect 303222 -7302 303306 -7066
rect 303542 -7302 322986 -7066
rect 323222 -7302 323306 -7066
rect 323542 -7302 342986 -7066
rect 343222 -7302 343306 -7066
rect 343542 -7302 362986 -7066
rect 363222 -7302 363306 -7066
rect 363542 -7302 382986 -7066
rect 383222 -7302 383306 -7066
rect 383542 -7302 402986 -7066
rect 403222 -7302 403306 -7066
rect 403542 -7302 422986 -7066
rect 423222 -7302 423306 -7066
rect 423542 -7302 442986 -7066
rect 443222 -7302 443306 -7066
rect 443542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 482986 -7066
rect 483222 -7302 483306 -7066
rect 483542 -7302 502986 -7066
rect 503222 -7302 503306 -7066
rect 503542 -7302 522986 -7066
rect 523222 -7302 523306 -7066
rect 523542 -7302 542986 -7066
rect 543222 -7302 543306 -7066
rect 543542 -7302 562986 -7066
rect 563222 -7302 563306 -7066
rect 563542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 22986 -7386
rect 23222 -7622 23306 -7386
rect 23542 -7622 42986 -7386
rect 43222 -7622 43306 -7386
rect 43542 -7622 62986 -7386
rect 63222 -7622 63306 -7386
rect 63542 -7622 82986 -7386
rect 83222 -7622 83306 -7386
rect 83542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 122986 -7386
rect 123222 -7622 123306 -7386
rect 123542 -7622 142986 -7386
rect 143222 -7622 143306 -7386
rect 143542 -7622 162986 -7386
rect 163222 -7622 163306 -7386
rect 163542 -7622 182986 -7386
rect 183222 -7622 183306 -7386
rect 183542 -7622 202986 -7386
rect 203222 -7622 203306 -7386
rect 203542 -7622 222986 -7386
rect 223222 -7622 223306 -7386
rect 223542 -7622 242986 -7386
rect 243222 -7622 243306 -7386
rect 243542 -7622 262986 -7386
rect 263222 -7622 263306 -7386
rect 263542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 302986 -7386
rect 303222 -7622 303306 -7386
rect 303542 -7622 322986 -7386
rect 323222 -7622 323306 -7386
rect 323542 -7622 342986 -7386
rect 343222 -7622 343306 -7386
rect 343542 -7622 362986 -7386
rect 363222 -7622 363306 -7386
rect 363542 -7622 382986 -7386
rect 383222 -7622 383306 -7386
rect 383542 -7622 402986 -7386
rect 403222 -7622 403306 -7386
rect 403542 -7622 422986 -7386
rect 423222 -7622 423306 -7386
rect 423542 -7622 442986 -7386
rect 443222 -7622 443306 -7386
rect 443542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 482986 -7386
rect 483222 -7622 483306 -7386
rect 483542 -7622 502986 -7386
rect 503222 -7622 503306 -7386
rect 503542 -7622 522986 -7386
rect 523222 -7622 523306 -7386
rect 523542 -7622 542986 -7386
rect 543222 -7622 543306 -7386
rect 543542 -7622 562986 -7386
rect 563222 -7622 563306 -7386
rect 563542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use Marmot  Marmot
timestamp 0
transform 1 0 200000 0 1 60000
box 0 0 357018 359162
use sky130_sram_2kbyte_1rw1r_32x512_8  data_arrays_0_0_ext_ram0h
timestamp 0
transform -1 0 166620 0 1 142000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  data_arrays_0_0_ext_ram0l
timestamp 0
transform -1 0 166620 0 1 30000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  data_arrays_0_0_ext_ram1h
timestamp 0
transform -1 0 166620 0 1 366000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  data_arrays_0_0_ext_ram1l
timestamp 0
transform -1 0 166620 0 1 254000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  data_arrays_0_0_ext_ram2h
timestamp 0
transform -1 0 166620 0 1 590000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  data_arrays_0_0_ext_ram2l
timestamp 0
transform -1 0 166620 0 1 478000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  data_arrays_0_0_ext_ram3h
timestamp 0
transform 1 0 410000 0 1 454000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  data_arrays_0_0_ext_ram3l
timestamp 0
transform -1 0 336620 0 1 454000
box 0 0 136620 83308
use sky130_sram_1kbyte_1rw1r_32x256_8  tag_array_ext_ram0h
timestamp 0
transform 1 0 410000 0 1 578000
box 0 0 95956 79500
use sky130_sram_1kbyte_1rw1r_32x256_8  tag_array_ext_ram0l
timestamp 0
transform -1 0 335956 0 1 578000
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2896 586890 3456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 22896 586890 23456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 42896 586890 43456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 62896 586890 63456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 82896 586890 83456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 102896 586890 103456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 122896 586890 123456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 142896 586890 143456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 162896 586890 163456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182896 586890 183456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 202896 586890 203456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 222896 586890 223456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 242896 586890 243456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 262896 586890 263456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 282896 586890 283456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 302896 586890 303456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 322896 586890 323456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 342896 586890 343456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362896 586890 363456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 382896 586890 383456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 402896 586890 403456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 422896 586890 423456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 442896 586890 443456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 462896 586890 463456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 482896 586890 483456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 502896 586890 503456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 522896 586890 523456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542896 586890 543456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 562896 586890 563456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 582896 586890 583456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 602896 586890 603456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 622896 586890 623456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 642896 586890 643456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 662896 586890 663456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 682896 586890 683456 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 41794 -1894 42414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 61794 -1894 62414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 81794 -1894 82414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 101794 -1894 102414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 121794 -1894 122414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 141794 -1894 142414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 161794 -1894 162414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 201794 -1894 202414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 221794 -1894 222414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 241794 -1894 242414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 261794 -1894 262414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 281794 -1894 282414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 301794 -1894 302414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 321794 -1894 322414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 341794 -1894 342414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 381794 -1894 382414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 401794 -1894 402414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 421794 -1894 422414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 441794 -1894 442414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 461794 -1894 462414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 481794 -1894 482414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 501794 -1894 502414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 521794 -1894 522414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 41794 115308 42414 140000 6 vccd1
port 531 nsew power input
rlabel metal4 s 61794 115308 62414 140000 6 vccd1
port 531 nsew power input
rlabel metal4 s 81794 115308 82414 140000 6 vccd1
port 531 nsew power input
rlabel metal4 s 101794 115308 102414 140000 6 vccd1
port 531 nsew power input
rlabel metal4 s 121794 115308 122414 140000 6 vccd1
port 531 nsew power input
rlabel metal4 s 141794 115308 142414 140000 6 vccd1
port 531 nsew power input
rlabel metal4 s 161794 115308 162414 140000 6 vccd1
port 531 nsew power input
rlabel metal4 s 41794 227308 42414 252000 6 vccd1
port 531 nsew power input
rlabel metal4 s 61794 227308 62414 252000 6 vccd1
port 531 nsew power input
rlabel metal4 s 81794 227308 82414 252000 6 vccd1
port 531 nsew power input
rlabel metal4 s 101794 227308 102414 252000 6 vccd1
port 531 nsew power input
rlabel metal4 s 121794 227308 122414 252000 6 vccd1
port 531 nsew power input
rlabel metal4 s 141794 227308 142414 252000 6 vccd1
port 531 nsew power input
rlabel metal4 s 161794 227308 162414 252000 6 vccd1
port 531 nsew power input
rlabel metal4 s 41794 339308 42414 364000 6 vccd1
port 531 nsew power input
rlabel metal4 s 61794 339308 62414 364000 6 vccd1
port 531 nsew power input
rlabel metal4 s 81794 339308 82414 364000 6 vccd1
port 531 nsew power input
rlabel metal4 s 101794 339308 102414 364000 6 vccd1
port 531 nsew power input
rlabel metal4 s 121794 339308 122414 364000 6 vccd1
port 531 nsew power input
rlabel metal4 s 141794 339308 142414 364000 6 vccd1
port 531 nsew power input
rlabel metal4 s 161794 339308 162414 364000 6 vccd1
port 531 nsew power input
rlabel metal4 s 201794 421162 202414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 221794 421162 222414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 241794 421162 242414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 261794 421162 262414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 281794 421162 282414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 301794 421162 302414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 321794 421162 322414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 421794 421162 422414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 441794 421162 442414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 461794 421162 462414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 481794 421162 482414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 501794 421162 502414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 521794 421162 522414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 421162 542414 452000 6 vccd1
port 531 nsew power input
rlabel metal4 s 41794 451308 42414 476000 6 vccd1
port 531 nsew power input
rlabel metal4 s 61794 451308 62414 476000 6 vccd1
port 531 nsew power input
rlabel metal4 s 81794 451308 82414 476000 6 vccd1
port 531 nsew power input
rlabel metal4 s 101794 451308 102414 476000 6 vccd1
port 531 nsew power input
rlabel metal4 s 121794 451308 122414 476000 6 vccd1
port 531 nsew power input
rlabel metal4 s 141794 451308 142414 476000 6 vccd1
port 531 nsew power input
rlabel metal4 s 161794 451308 162414 476000 6 vccd1
port 531 nsew power input
rlabel metal4 s 241794 539308 242414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 261794 539308 262414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 281794 539308 282414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 301794 539308 302414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 321794 539308 322414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 421794 539308 422414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 441794 539308 442414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 461794 539308 462414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 481794 539308 482414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 501794 539308 502414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 41794 563308 42414 588000 6 vccd1
port 531 nsew power input
rlabel metal4 s 61794 563308 62414 588000 6 vccd1
port 531 nsew power input
rlabel metal4 s 81794 563308 82414 588000 6 vccd1
port 531 nsew power input
rlabel metal4 s 101794 563308 102414 588000 6 vccd1
port 531 nsew power input
rlabel metal4 s 121794 563308 122414 588000 6 vccd1
port 531 nsew power input
rlabel metal4 s 141794 563308 142414 588000 6 vccd1
port 531 nsew power input
rlabel metal4 s 161794 563308 162414 588000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 21794 -1894 22414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 41794 675308 42414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 61794 675308 62414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 81794 675308 82414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 101794 675308 102414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 121794 675308 122414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 141794 675308 142414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 161794 675308 162414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 201794 539308 202414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 221794 539308 222414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 241794 659500 242414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 261794 659500 262414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 281794 659500 282414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 301794 659500 302414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 321794 659500 322414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 341794 421162 342414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 421162 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 381794 421162 382414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 401794 421162 402414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 421794 659500 422414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 441794 659500 442414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 461794 659500 462414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 481794 659500 482414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 501794 659500 502414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 521794 539308 522414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 539308 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 561794 -1894 562414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 581794 -1894 582414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6556 588810 7116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 26556 588810 27116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 46556 588810 47116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 66556 588810 67116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 86556 588810 87116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 106556 588810 107116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 126556 588810 127116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 146556 588810 147116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 166556 588810 167116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186556 588810 187116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 206556 588810 207116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 226556 588810 227116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 246556 588810 247116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 266556 588810 267116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 286556 588810 287116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 306556 588810 307116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 326556 588810 327116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 346556 588810 347116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366556 588810 367116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 386556 588810 387116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 406556 588810 407116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 426556 588810 427116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 446556 588810 447116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 466556 588810 467116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 486556 588810 487116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 506556 588810 507116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 526556 588810 527116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546556 588810 547116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 566556 588810 567116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 586556 588810 587116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 606556 588810 607116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 626556 588810 627116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 646556 588810 647116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 666556 588810 667116 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 686556 588810 687116 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 45514 -3814 46134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 65514 -3814 66134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 85514 -3814 86134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 105514 -3814 106134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 125514 -3814 126134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 145514 -3814 146134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 165514 -3814 166134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 205514 -3814 206134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 225514 -3814 226134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 245514 -3814 246134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 265514 -3814 266134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 285514 -3814 286134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 305514 -3814 306134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 325514 -3814 326134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 345514 -3814 346134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 385514 -3814 386134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 405514 -3814 406134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 425514 -3814 426134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 445514 -3814 446134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 465514 -3814 466134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 485514 -3814 486134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 505514 -3814 506134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 525514 -3814 526134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 45514 115308 46134 140000 6 vccd2
port 532 nsew power input
rlabel metal4 s 65514 115308 66134 140000 6 vccd2
port 532 nsew power input
rlabel metal4 s 85514 115308 86134 140000 6 vccd2
port 532 nsew power input
rlabel metal4 s 105514 115308 106134 140000 6 vccd2
port 532 nsew power input
rlabel metal4 s 125514 115308 126134 140000 6 vccd2
port 532 nsew power input
rlabel metal4 s 145514 115308 146134 140000 6 vccd2
port 532 nsew power input
rlabel metal4 s 165514 115308 166134 140000 6 vccd2
port 532 nsew power input
rlabel metal4 s 45514 227308 46134 252000 6 vccd2
port 532 nsew power input
rlabel metal4 s 65514 227308 66134 252000 6 vccd2
port 532 nsew power input
rlabel metal4 s 85514 227308 86134 252000 6 vccd2
port 532 nsew power input
rlabel metal4 s 105514 227308 106134 252000 6 vccd2
port 532 nsew power input
rlabel metal4 s 125514 227308 126134 252000 6 vccd2
port 532 nsew power input
rlabel metal4 s 145514 227308 146134 252000 6 vccd2
port 532 nsew power input
rlabel metal4 s 165514 227308 166134 252000 6 vccd2
port 532 nsew power input
rlabel metal4 s 45514 339308 46134 364000 6 vccd2
port 532 nsew power input
rlabel metal4 s 65514 339308 66134 364000 6 vccd2
port 532 nsew power input
rlabel metal4 s 85514 339308 86134 364000 6 vccd2
port 532 nsew power input
rlabel metal4 s 105514 339308 106134 364000 6 vccd2
port 532 nsew power input
rlabel metal4 s 125514 339308 126134 364000 6 vccd2
port 532 nsew power input
rlabel metal4 s 145514 339308 146134 364000 6 vccd2
port 532 nsew power input
rlabel metal4 s 165514 339308 166134 364000 6 vccd2
port 532 nsew power input
rlabel metal4 s 205514 421162 206134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 225514 421162 226134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 245514 421162 246134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 265514 421162 266134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 285514 421162 286134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 305514 421162 306134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 325514 421162 326134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 425514 421162 426134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 445514 421162 446134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 465514 421162 466134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 485514 421162 486134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 505514 421162 506134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 525514 421162 526134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 421162 546134 452000 6 vccd2
port 532 nsew power input
rlabel metal4 s 45514 451308 46134 476000 6 vccd2
port 532 nsew power input
rlabel metal4 s 65514 451308 66134 476000 6 vccd2
port 532 nsew power input
rlabel metal4 s 85514 451308 86134 476000 6 vccd2
port 532 nsew power input
rlabel metal4 s 105514 451308 106134 476000 6 vccd2
port 532 nsew power input
rlabel metal4 s 125514 451308 126134 476000 6 vccd2
port 532 nsew power input
rlabel metal4 s 145514 451308 146134 476000 6 vccd2
port 532 nsew power input
rlabel metal4 s 165514 451308 166134 476000 6 vccd2
port 532 nsew power input
rlabel metal4 s 245514 539308 246134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 265514 539308 266134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 285514 539308 286134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 305514 539308 306134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 325514 539308 326134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 425514 539308 426134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 445514 539308 446134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 465514 539308 466134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 485514 539308 486134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 505514 539308 506134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 45514 563308 46134 588000 6 vccd2
port 532 nsew power input
rlabel metal4 s 65514 563308 66134 588000 6 vccd2
port 532 nsew power input
rlabel metal4 s 85514 563308 86134 588000 6 vccd2
port 532 nsew power input
rlabel metal4 s 105514 563308 106134 588000 6 vccd2
port 532 nsew power input
rlabel metal4 s 125514 563308 126134 588000 6 vccd2
port 532 nsew power input
rlabel metal4 s 145514 563308 146134 588000 6 vccd2
port 532 nsew power input
rlabel metal4 s 165514 563308 166134 588000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 25514 -3814 26134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 45514 675308 46134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 65514 675308 66134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 85514 675308 86134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 105514 675308 106134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 125514 675308 126134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 145514 675308 146134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 165514 675308 166134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 205514 539308 206134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 225514 539308 226134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 245514 659500 246134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 265514 659500 266134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 285514 659500 286134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 305514 659500 306134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 325514 659500 326134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 345514 421162 346134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 421162 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 385514 421162 386134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 405514 421162 406134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 425514 659500 426134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 445514 659500 446134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 465514 659500 466134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 485514 659500 486134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 505514 659500 506134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 525514 539308 526134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 539308 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 565514 -3814 566134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10216 590730 10776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 30216 590730 30776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 50216 590730 50776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 70216 590730 70776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 90216 590730 90776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 110216 590730 110776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 130216 590730 130776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 150216 590730 150776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 170216 590730 170776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190216 590730 190776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 210216 590730 210776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 230216 590730 230776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 250216 590730 250776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 270216 590730 270776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 290216 590730 290776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 310216 590730 310776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 330216 590730 330776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 350216 590730 350776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370216 590730 370776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 390216 590730 390776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 410216 590730 410776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 430216 590730 430776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 450216 590730 450776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 470216 590730 470776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 490216 590730 490776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 510216 590730 510776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 530216 590730 530776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550216 590730 550776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 570216 590730 570776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 590216 590730 590776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 610216 590730 610776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 630216 590730 630776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 650216 590730 650776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 670216 590730 670776 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 690216 590730 690776 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 29234 -5734 29854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 49234 -5734 49854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 69234 -5734 69854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 89234 -5734 89854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 109234 -5734 109854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 129234 -5734 129854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 149234 -5734 149854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 209234 -5734 209854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 229234 -5734 229854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 249234 -5734 249854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 269234 -5734 269854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 289234 -5734 289854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 309234 -5734 309854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 329234 -5734 329854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 349234 -5734 349854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 389234 -5734 389854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 409234 -5734 409854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 429234 -5734 429854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 449234 -5734 449854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 469234 -5734 469854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 489234 -5734 489854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 509234 -5734 509854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 529234 -5734 529854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 29234 115308 29854 140000 6 vdda1
port 533 nsew power input
rlabel metal4 s 49234 115308 49854 140000 6 vdda1
port 533 nsew power input
rlabel metal4 s 69234 115308 69854 140000 6 vdda1
port 533 nsew power input
rlabel metal4 s 89234 115308 89854 140000 6 vdda1
port 533 nsew power input
rlabel metal4 s 109234 115308 109854 140000 6 vdda1
port 533 nsew power input
rlabel metal4 s 129234 115308 129854 140000 6 vdda1
port 533 nsew power input
rlabel metal4 s 149234 115308 149854 140000 6 vdda1
port 533 nsew power input
rlabel metal4 s 29234 227308 29854 252000 6 vdda1
port 533 nsew power input
rlabel metal4 s 49234 227308 49854 252000 6 vdda1
port 533 nsew power input
rlabel metal4 s 69234 227308 69854 252000 6 vdda1
port 533 nsew power input
rlabel metal4 s 89234 227308 89854 252000 6 vdda1
port 533 nsew power input
rlabel metal4 s 109234 227308 109854 252000 6 vdda1
port 533 nsew power input
rlabel metal4 s 129234 227308 129854 252000 6 vdda1
port 533 nsew power input
rlabel metal4 s 149234 227308 149854 252000 6 vdda1
port 533 nsew power input
rlabel metal4 s 29234 339308 29854 364000 6 vdda1
port 533 nsew power input
rlabel metal4 s 49234 339308 49854 364000 6 vdda1
port 533 nsew power input
rlabel metal4 s 69234 339308 69854 364000 6 vdda1
port 533 nsew power input
rlabel metal4 s 89234 339308 89854 364000 6 vdda1
port 533 nsew power input
rlabel metal4 s 109234 339308 109854 364000 6 vdda1
port 533 nsew power input
rlabel metal4 s 129234 339308 129854 364000 6 vdda1
port 533 nsew power input
rlabel metal4 s 149234 339308 149854 364000 6 vdda1
port 533 nsew power input
rlabel metal4 s 209234 421162 209854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 229234 421162 229854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 249234 421162 249854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 269234 421162 269854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 289234 421162 289854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 309234 421162 309854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 329234 421162 329854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 409234 421162 409854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 429234 421162 429854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 449234 421162 449854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 469234 421162 469854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 489234 421162 489854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 509234 421162 509854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 529234 421162 529854 452000 6 vdda1
port 533 nsew power input
rlabel metal4 s 29234 451308 29854 476000 6 vdda1
port 533 nsew power input
rlabel metal4 s 49234 451308 49854 476000 6 vdda1
port 533 nsew power input
rlabel metal4 s 69234 451308 69854 476000 6 vdda1
port 533 nsew power input
rlabel metal4 s 89234 451308 89854 476000 6 vdda1
port 533 nsew power input
rlabel metal4 s 109234 451308 109854 476000 6 vdda1
port 533 nsew power input
rlabel metal4 s 129234 451308 129854 476000 6 vdda1
port 533 nsew power input
rlabel metal4 s 149234 451308 149854 476000 6 vdda1
port 533 nsew power input
rlabel metal4 s 249234 539308 249854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 269234 539308 269854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 289234 539308 289854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 309234 539308 309854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 329234 539308 329854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 409234 539308 409854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 429234 539308 429854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 449234 539308 449854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 469234 539308 469854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 489234 539308 489854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s 29234 563308 29854 588000 6 vdda1
port 533 nsew power input
rlabel metal4 s 49234 563308 49854 588000 6 vdda1
port 533 nsew power input
rlabel metal4 s 69234 563308 69854 588000 6 vdda1
port 533 nsew power input
rlabel metal4 s 89234 563308 89854 588000 6 vdda1
port 533 nsew power input
rlabel metal4 s 109234 563308 109854 588000 6 vdda1
port 533 nsew power input
rlabel metal4 s 129234 563308 129854 588000 6 vdda1
port 533 nsew power input
rlabel metal4 s 149234 563308 149854 588000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 29234 675308 29854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 49234 675308 49854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 69234 675308 69854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 89234 675308 89854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 109234 675308 109854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 129234 675308 129854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 149234 675308 149854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 169234 -5734 169854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 209234 539308 209854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 229234 539308 229854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 249234 659500 249854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 269234 659500 269854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 289234 659500 289854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 309234 659500 309854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 329234 659500 329854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 349234 421162 349854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 421162 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 389234 421162 389854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 409234 659500 409854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 429234 659500 429854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 449234 659500 449854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 469234 659500 469854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 489234 659500 489854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 509234 539308 509854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 529234 539308 529854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 421162 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 569234 -5734 569854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 13876 592650 14436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 33876 592650 34436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 53876 592650 54436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 73876 592650 74436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 93876 592650 94436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 113876 592650 114436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 133876 592650 134436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 153876 592650 154436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 173876 592650 174436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 193876 592650 194436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 213876 592650 214436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 233876 592650 234436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 253876 592650 254436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 273876 592650 274436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 293876 592650 294436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 313876 592650 314436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 333876 592650 334436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 353876 592650 354436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 373876 592650 374436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 393876 592650 394436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 413876 592650 414436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 433876 592650 434436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 453876 592650 454436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 473876 592650 474436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 493876 592650 494436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 513876 592650 514436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 533876 592650 534436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 553876 592650 554436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 573876 592650 574436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 593876 592650 594436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 613876 592650 614436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 633876 592650 634436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 653876 592650 654436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 673876 592650 674436 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 693876 592650 694436 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 32954 -7654 33574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 52954 -7654 53574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 72954 -7654 73574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 92954 -7654 93574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 112954 -7654 113574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 132954 -7654 133574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 152954 -7654 153574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 212954 -7654 213574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 232954 -7654 233574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 252954 -7654 253574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 272954 -7654 273574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 292954 -7654 293574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 312954 -7654 313574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 332954 -7654 333574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 352954 -7654 353574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 392954 -7654 393574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 412954 -7654 413574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 432954 -7654 433574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 452954 -7654 453574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 472954 -7654 473574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 492954 -7654 493574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 512954 -7654 513574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 532954 -7654 533574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 32954 115308 33574 140000 6 vdda2
port 534 nsew power input
rlabel metal4 s 52954 115308 53574 140000 6 vdda2
port 534 nsew power input
rlabel metal4 s 72954 115308 73574 140000 6 vdda2
port 534 nsew power input
rlabel metal4 s 92954 115308 93574 140000 6 vdda2
port 534 nsew power input
rlabel metal4 s 112954 115308 113574 140000 6 vdda2
port 534 nsew power input
rlabel metal4 s 132954 115308 133574 140000 6 vdda2
port 534 nsew power input
rlabel metal4 s 152954 115308 153574 140000 6 vdda2
port 534 nsew power input
rlabel metal4 s 32954 227308 33574 252000 6 vdda2
port 534 nsew power input
rlabel metal4 s 52954 227308 53574 252000 6 vdda2
port 534 nsew power input
rlabel metal4 s 72954 227308 73574 252000 6 vdda2
port 534 nsew power input
rlabel metal4 s 92954 227308 93574 252000 6 vdda2
port 534 nsew power input
rlabel metal4 s 112954 227308 113574 252000 6 vdda2
port 534 nsew power input
rlabel metal4 s 132954 227308 133574 252000 6 vdda2
port 534 nsew power input
rlabel metal4 s 152954 227308 153574 252000 6 vdda2
port 534 nsew power input
rlabel metal4 s 32954 339308 33574 364000 6 vdda2
port 534 nsew power input
rlabel metal4 s 52954 339308 53574 364000 6 vdda2
port 534 nsew power input
rlabel metal4 s 72954 339308 73574 364000 6 vdda2
port 534 nsew power input
rlabel metal4 s 92954 339308 93574 364000 6 vdda2
port 534 nsew power input
rlabel metal4 s 112954 339308 113574 364000 6 vdda2
port 534 nsew power input
rlabel metal4 s 132954 339308 133574 364000 6 vdda2
port 534 nsew power input
rlabel metal4 s 152954 339308 153574 364000 6 vdda2
port 534 nsew power input
rlabel metal4 s 212954 421162 213574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 232954 421162 233574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 252954 421162 253574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 272954 421162 273574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 292954 421162 293574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 312954 421162 313574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 332954 421162 333574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 412954 421162 413574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 432954 421162 433574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 452954 421162 453574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 472954 421162 473574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 492954 421162 493574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 512954 421162 513574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 532954 421162 533574 452000 6 vdda2
port 534 nsew power input
rlabel metal4 s 32954 451308 33574 476000 6 vdda2
port 534 nsew power input
rlabel metal4 s 52954 451308 53574 476000 6 vdda2
port 534 nsew power input
rlabel metal4 s 72954 451308 73574 476000 6 vdda2
port 534 nsew power input
rlabel metal4 s 92954 451308 93574 476000 6 vdda2
port 534 nsew power input
rlabel metal4 s 112954 451308 113574 476000 6 vdda2
port 534 nsew power input
rlabel metal4 s 132954 451308 133574 476000 6 vdda2
port 534 nsew power input
rlabel metal4 s 152954 451308 153574 476000 6 vdda2
port 534 nsew power input
rlabel metal4 s 252954 539308 253574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 272954 539308 273574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 292954 539308 293574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 312954 539308 313574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 332954 539308 333574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 412954 539308 413574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 432954 539308 433574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 452954 539308 453574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 472954 539308 473574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 492954 539308 493574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s 32954 563308 33574 588000 6 vdda2
port 534 nsew power input
rlabel metal4 s 52954 563308 53574 588000 6 vdda2
port 534 nsew power input
rlabel metal4 s 72954 563308 73574 588000 6 vdda2
port 534 nsew power input
rlabel metal4 s 92954 563308 93574 588000 6 vdda2
port 534 nsew power input
rlabel metal4 s 112954 563308 113574 588000 6 vdda2
port 534 nsew power input
rlabel metal4 s 132954 563308 133574 588000 6 vdda2
port 534 nsew power input
rlabel metal4 s 152954 563308 153574 588000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 32954 675308 33574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 52954 675308 53574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 72954 675308 73574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 92954 675308 93574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 112954 675308 113574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 132954 675308 133574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 152954 675308 153574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 172954 -7654 173574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 212954 539308 213574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 232954 539308 233574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 252954 659500 253574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 272954 659500 273574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 292954 659500 293574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 312954 659500 313574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 332954 659500 333574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 352954 421162 353574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 421162 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 392954 421162 393574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 412954 659500 413574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 432954 659500 433574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 452954 659500 453574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 472954 659500 473574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 492954 659500 493574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 512954 539308 513574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 532954 539308 533574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 421162 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 572954 -7654 573574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 20216 590730 20776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 40216 590730 40776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 60216 590730 60776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 80216 590730 80776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100216 590730 100776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 120216 590730 120776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 140216 590730 140776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 160216 590730 160776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 180216 590730 180776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 200216 590730 200776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 220216 590730 220776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 240216 590730 240776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 260216 590730 260776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280216 590730 280776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 300216 590730 300776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 320216 590730 320776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 340216 590730 340776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 360216 590730 360776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 380216 590730 380776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 400216 590730 400776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 420216 590730 420776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 440216 590730 440776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460216 590730 460776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 480216 590730 480776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 500216 590730 500776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 520216 590730 520776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 540216 590730 540776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 560216 590730 560776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 580216 590730 580776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 600216 590730 600776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 620216 590730 620776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640216 590730 640776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 660216 590730 660776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 680216 590730 680776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 700216 590730 700776 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 39234 -5734 39854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 59234 -5734 59854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 79234 -5734 79854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 119234 -5734 119854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 139234 -5734 139854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 159234 -5734 159854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 199234 -5734 199854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 219234 -5734 219854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 239234 -5734 239854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 259234 -5734 259854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 299234 -5734 299854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 319234 -5734 319854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 339234 -5734 339854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 359234 -5734 359854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 379234 -5734 379854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 399234 -5734 399854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 419234 -5734 419854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 439234 -5734 439854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 479234 -5734 479854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 499234 -5734 499854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 519234 -5734 519854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 539234 -5734 539854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 39234 115308 39854 140000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 59234 115308 59854 140000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 79234 115308 79854 140000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 115308 99854 140000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 119234 115308 119854 140000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 139234 115308 139854 140000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 159234 115308 159854 140000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 39234 227308 39854 252000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 59234 227308 59854 252000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 79234 227308 79854 252000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 227308 99854 252000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 119234 227308 119854 252000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 139234 227308 139854 252000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 159234 227308 159854 252000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 39234 339308 39854 364000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 59234 339308 59854 364000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 79234 339308 79854 364000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 339308 99854 364000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 119234 339308 119854 364000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 139234 339308 139854 364000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 159234 339308 159854 364000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 199234 421162 199854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 219234 421162 219854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 239234 421162 239854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 259234 421162 259854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 421162 279854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 299234 421162 299854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 319234 421162 319854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 419234 421162 419854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 439234 421162 439854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 421162 459854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 479234 421162 479854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 499234 421162 499854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 519234 421162 519854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 539234 421162 539854 452000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 39234 451308 39854 476000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 59234 451308 59854 476000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 79234 451308 79854 476000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 451308 99854 476000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 119234 451308 119854 476000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 139234 451308 139854 476000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 159234 451308 159854 476000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 239234 539308 239854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 259234 539308 259854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 539308 279854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 299234 539308 299854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 319234 539308 319854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 419234 539308 419854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 439234 539308 439854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 539308 459854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 479234 539308 479854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 499234 539308 499854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 39234 563308 39854 588000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 59234 563308 59854 588000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 79234 563308 79854 588000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 563308 99854 588000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 119234 563308 119854 588000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 139234 563308 139854 588000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 159234 563308 159854 588000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 19234 -5734 19854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 39234 675308 39854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 59234 675308 59854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 79234 675308 79854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 675308 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 119234 675308 119854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 139234 675308 139854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 159234 675308 159854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 179234 -5734 179854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 199234 539308 199854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 219234 539308 219854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 239234 659500 239854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 259234 659500 259854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 659500 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 299234 659500 299854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 319234 659500 319854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 339234 421162 339854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 359234 421162 359854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 379234 421162 379854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 399234 421162 399854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 419234 659500 419854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 439234 659500 439854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 659500 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 479234 659500 479854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 499234 659500 499854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 519234 539308 519854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 539234 539308 539854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 559234 -5734 559854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 579234 -5734 579854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 23876 592650 24436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 43876 592650 44436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 63876 592650 64436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 83876 592650 84436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 103876 592650 104436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 123876 592650 124436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 143876 592650 144436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 163876 592650 164436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 183876 592650 184436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 203876 592650 204436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 223876 592650 224436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 243876 592650 244436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 263876 592650 264436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 283876 592650 284436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 303876 592650 304436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 323876 592650 324436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 343876 592650 344436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 363876 592650 364436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 383876 592650 384436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 403876 592650 404436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 423876 592650 424436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 443876 592650 444436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 463876 592650 464436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 483876 592650 484436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 503876 592650 504436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 523876 592650 524436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 543876 592650 544436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 563876 592650 564436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 583876 592650 584436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 603876 592650 604436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 623876 592650 624436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 643876 592650 644436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 663876 592650 664436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 683876 592650 684436 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 42954 -7654 43574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 62954 -7654 63574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 82954 -7654 83574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 122954 -7654 123574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 142954 -7654 143574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 162954 -7654 163574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 202954 -7654 203574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 222954 -7654 223574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 242954 -7654 243574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 262954 -7654 263574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 302954 -7654 303574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 322954 -7654 323574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 342954 -7654 343574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 362954 -7654 363574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 382954 -7654 383574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 402954 -7654 403574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 422954 -7654 423574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 442954 -7654 443574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 482954 -7654 483574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 502954 -7654 503574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 522954 -7654 523574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 542954 -7654 543574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 42954 115308 43574 140000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 62954 115308 63574 140000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 82954 115308 83574 140000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 115308 103574 140000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 122954 115308 123574 140000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 142954 115308 143574 140000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 162954 115308 163574 140000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 42954 227308 43574 252000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 62954 227308 63574 252000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 82954 227308 83574 252000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 227308 103574 252000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 122954 227308 123574 252000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 142954 227308 143574 252000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 162954 227308 163574 252000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 42954 339308 43574 364000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 62954 339308 63574 364000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 82954 339308 83574 364000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 339308 103574 364000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 122954 339308 123574 364000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 142954 339308 143574 364000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 162954 339308 163574 364000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 202954 421162 203574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 222954 421162 223574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 242954 421162 243574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 262954 421162 263574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 421162 283574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 302954 421162 303574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 322954 421162 323574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 422954 421162 423574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 442954 421162 443574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 421162 463574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 482954 421162 483574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 502954 421162 503574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 522954 421162 523574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 542954 421162 543574 452000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 42954 451308 43574 476000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 62954 451308 63574 476000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 82954 451308 83574 476000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 451308 103574 476000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 122954 451308 123574 476000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 142954 451308 143574 476000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 162954 451308 163574 476000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 242954 539308 243574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 262954 539308 263574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 539308 283574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 302954 539308 303574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 322954 539308 323574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 422954 539308 423574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 442954 539308 443574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 539308 463574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 482954 539308 483574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 502954 539308 503574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 42954 563308 43574 588000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 62954 563308 63574 588000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 82954 563308 83574 588000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 563308 103574 588000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 122954 563308 123574 588000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 142954 563308 143574 588000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 162954 563308 163574 588000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 22954 -7654 23574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 42954 675308 43574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 62954 675308 63574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 82954 675308 83574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 675308 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 122954 675308 123574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 142954 675308 143574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 162954 675308 163574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 182954 -7654 183574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 202954 539308 203574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 222954 539308 223574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 242954 659500 243574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 262954 659500 263574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 659500 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 302954 659500 303574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 322954 659500 323574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 342954 421162 343574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 362954 421162 363574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 382954 421162 383574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 402954 421162 403574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 422954 659500 423574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 442954 659500 443574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 659500 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 482954 659500 483574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 502954 659500 503574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 522954 539308 523574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 542954 539308 543574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 562954 -7654 563574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 12896 586890 13456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 32896 586890 33456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 52896 586890 53456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 72896 586890 73456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92896 586890 93456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 112896 586890 113456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 132896 586890 133456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 152896 586890 153456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 172896 586890 173456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 192896 586890 193456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 212896 586890 213456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 232896 586890 233456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 252896 586890 253456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272896 586890 273456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 292896 586890 293456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 312896 586890 313456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 332896 586890 333456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 352896 586890 353456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 372896 586890 373456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 392896 586890 393456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 412896 586890 413456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 432896 586890 433456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452896 586890 453456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 472896 586890 473456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 492896 586890 493456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 512896 586890 513456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 532896 586890 533456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 552896 586890 553456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 572896 586890 573456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 592896 586890 593456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 612896 586890 613456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632896 586890 633456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 652896 586890 653456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 672896 586890 673456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 692896 586890 693456 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 31794 -1894 32414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 51794 -1894 52414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 71794 -1894 72414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 111794 -1894 112414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 131794 -1894 132414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 151794 -1894 152414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 211794 -1894 212414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 231794 -1894 232414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 251794 -1894 252414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 291794 -1894 292414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 311794 -1894 312414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 331794 -1894 332414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 351794 -1894 352414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 371794 -1894 372414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 391794 -1894 392414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 411794 -1894 412414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 431794 -1894 432414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 471794 -1894 472414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 491794 -1894 492414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 511794 -1894 512414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 531794 -1894 532414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 551794 -1894 552414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 31794 115308 32414 140000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 51794 115308 52414 140000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 71794 115308 72414 140000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 115308 92414 140000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 111794 115308 112414 140000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 131794 115308 132414 140000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 151794 115308 152414 140000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 31794 227308 32414 252000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 51794 227308 52414 252000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 71794 227308 72414 252000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 227308 92414 252000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 111794 227308 112414 252000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 131794 227308 132414 252000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 151794 227308 152414 252000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 31794 339308 32414 364000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 51794 339308 52414 364000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 71794 339308 72414 364000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 339308 92414 364000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 111794 339308 112414 364000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 131794 339308 132414 364000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 151794 339308 152414 364000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 211794 421162 212414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 231794 421162 232414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 251794 421162 252414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 421162 272414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 291794 421162 292414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 311794 421162 312414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 331794 421162 332414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 411794 421162 412414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 431794 421162 432414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 421162 452414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 471794 421162 472414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 491794 421162 492414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 511794 421162 512414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 531794 421162 532414 452000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 31794 451308 32414 476000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 51794 451308 52414 476000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 71794 451308 72414 476000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 451308 92414 476000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 111794 451308 112414 476000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 131794 451308 132414 476000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 151794 451308 152414 476000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 251794 539308 252414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 539308 272414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 291794 539308 292414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 311794 539308 312414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 331794 539308 332414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 411794 539308 412414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 431794 539308 432414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 539308 452414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 471794 539308 472414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 491794 539308 492414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 31794 563308 32414 588000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 51794 563308 52414 588000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 71794 563308 72414 588000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 563308 92414 588000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 111794 563308 112414 588000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 131794 563308 132414 588000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 151794 563308 152414 588000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 11794 -1894 12414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 31794 675308 32414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 51794 675308 52414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 71794 675308 72414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 675308 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 111794 675308 112414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 131794 675308 132414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 151794 675308 152414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 171794 -1894 172414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 191794 -1894 192414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 211794 539308 212414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 231794 539308 232414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 251794 659500 252414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 659500 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 291794 659500 292414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 311794 659500 312414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 331794 659500 332414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 351794 421162 352414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 371794 421162 372414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 391794 421162 392414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 411794 659500 412414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 431794 659500 432414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 659500 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 471794 659500 472414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 491794 659500 492414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 511794 539308 512414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 531794 539308 532414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 551794 421162 552414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 571794 -1894 572414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 16556 588810 17116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 36556 588810 37116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 56556 588810 57116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 76556 588810 77116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96556 588810 97116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 116556 588810 117116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 136556 588810 137116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 156556 588810 157116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 176556 588810 177116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 196556 588810 197116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 216556 588810 217116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 236556 588810 237116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 256556 588810 257116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276556 588810 277116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 296556 588810 297116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 316556 588810 317116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 336556 588810 337116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 356556 588810 357116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 376556 588810 377116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 396556 588810 397116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 416556 588810 417116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 436556 588810 437116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456556 588810 457116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 476556 588810 477116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 496556 588810 497116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 516556 588810 517116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 536556 588810 537116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 556556 588810 557116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 576556 588810 577116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 596556 588810 597116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 616556 588810 617116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636556 588810 637116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 656556 588810 657116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 676556 588810 677116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 696556 588810 697116 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 35514 -3814 36134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 55514 -3814 56134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 75514 -3814 76134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 115514 -3814 116134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 135514 -3814 136134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 155514 -3814 156134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 215514 -3814 216134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 235514 -3814 236134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 255514 -3814 256134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 295514 -3814 296134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 315514 -3814 316134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 335514 -3814 336134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 355514 -3814 356134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 375514 -3814 376134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 395514 -3814 396134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 415514 -3814 416134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 435514 -3814 436134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 475514 -3814 476134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 495514 -3814 496134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 515514 -3814 516134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 535514 -3814 536134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 555514 -3814 556134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 35514 115308 36134 140000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 55514 115308 56134 140000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 75514 115308 76134 140000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 115308 96134 140000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 115514 115308 116134 140000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 135514 115308 136134 140000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 155514 115308 156134 140000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 35514 227308 36134 252000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 55514 227308 56134 252000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 75514 227308 76134 252000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 227308 96134 252000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 115514 227308 116134 252000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 135514 227308 136134 252000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 155514 227308 156134 252000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 35514 339308 36134 364000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 55514 339308 56134 364000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 75514 339308 76134 364000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 339308 96134 364000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 115514 339308 116134 364000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 135514 339308 136134 364000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 155514 339308 156134 364000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 215514 421162 216134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 235514 421162 236134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 255514 421162 256134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 421162 276134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 295514 421162 296134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 315514 421162 316134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 335514 421162 336134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 415514 421162 416134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 435514 421162 436134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 421162 456134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 475514 421162 476134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 495514 421162 496134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 515514 421162 516134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 535514 421162 536134 452000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 35514 451308 36134 476000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 55514 451308 56134 476000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 75514 451308 76134 476000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 451308 96134 476000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 115514 451308 116134 476000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 135514 451308 136134 476000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 155514 451308 156134 476000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 255514 539308 256134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 539308 276134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 295514 539308 296134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 315514 539308 316134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 335514 539308 336134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 415514 539308 416134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 435514 539308 436134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 539308 456134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 475514 539308 476134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 495514 539308 496134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 35514 563308 36134 588000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 55514 563308 56134 588000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 75514 563308 76134 588000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 563308 96134 588000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 115514 563308 116134 588000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 135514 563308 136134 588000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 155514 563308 156134 588000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 15514 -3814 16134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 35514 675308 36134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 55514 675308 56134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 75514 675308 76134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 675308 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 115514 675308 116134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 135514 675308 136134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 155514 675308 156134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 175514 -3814 176134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 195514 -3814 196134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 215514 539308 216134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 235514 539308 236134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 255514 659500 256134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 659500 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 295514 659500 296134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 315514 659500 316134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 335514 659500 336134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 355514 421162 356134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 375514 421162 376134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 395514 421162 396134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 415514 659500 416134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 435514 659500 436134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 659500 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 475514 659500 476134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 495514 659500 496134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 515514 539308 516134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 535514 539308 536134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 555514 421162 556134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 575514 -3814 576134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
