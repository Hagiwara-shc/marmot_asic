magic
tech sky130A
magscale 1 2
timestamp 1647885048
<< obsli1 >>
rect 1104 2159 350060 350897
<< obsm1 >>
rect 290 1980 350874 352844
<< metal2 >>
rect 478 352563 534 353363
rect 1490 352563 1546 353363
rect 2594 352563 2650 353363
rect 3606 352563 3662 353363
rect 4710 352563 4766 353363
rect 5814 352563 5870 353363
rect 6826 352563 6882 353363
rect 7930 352563 7986 353363
rect 8942 352563 8998 353363
rect 10046 352563 10102 353363
rect 11150 352563 11206 353363
rect 12162 352563 12218 353363
rect 13266 352563 13322 353363
rect 14278 352563 14334 353363
rect 15382 352563 15438 353363
rect 16486 352563 16542 353363
rect 17498 352563 17554 353363
rect 18602 352563 18658 353363
rect 19614 352563 19670 353363
rect 20718 352563 20774 353363
rect 21822 352563 21878 353363
rect 22834 352563 22890 353363
rect 23938 352563 23994 353363
rect 24950 352563 25006 353363
rect 26054 352563 26110 353363
rect 27158 352563 27214 353363
rect 28170 352563 28226 353363
rect 29274 352563 29330 353363
rect 30286 352563 30342 353363
rect 31390 352563 31446 353363
rect 32494 352563 32550 353363
rect 33506 352563 33562 353363
rect 34610 352563 34666 353363
rect 35622 352563 35678 353363
rect 36726 352563 36782 353363
rect 37830 352563 37886 353363
rect 38842 352563 38898 353363
rect 39946 352563 40002 353363
rect 40958 352563 41014 353363
rect 42062 352563 42118 353363
rect 43166 352563 43222 353363
rect 44178 352563 44234 353363
rect 45282 352563 45338 353363
rect 46386 352563 46442 353363
rect 47398 352563 47454 353363
rect 48502 352563 48558 353363
rect 49514 352563 49570 353363
rect 50618 352563 50674 353363
rect 51722 352563 51778 353363
rect 52734 352563 52790 353363
rect 53838 352563 53894 353363
rect 54850 352563 54906 353363
rect 55954 352563 56010 353363
rect 57058 352563 57114 353363
rect 58070 352563 58126 353363
rect 59174 352563 59230 353363
rect 60186 352563 60242 353363
rect 61290 352563 61346 353363
rect 62394 352563 62450 353363
rect 63406 352563 63462 353363
rect 64510 352563 64566 353363
rect 65522 352563 65578 353363
rect 66626 352563 66682 353363
rect 67730 352563 67786 353363
rect 68742 352563 68798 353363
rect 69846 352563 69902 353363
rect 70858 352563 70914 353363
rect 71962 352563 72018 353363
rect 73066 352563 73122 353363
rect 74078 352563 74134 353363
rect 75182 352563 75238 353363
rect 76194 352563 76250 353363
rect 77298 352563 77354 353363
rect 78402 352563 78458 353363
rect 79414 352563 79470 353363
rect 80518 352563 80574 353363
rect 81530 352563 81586 353363
rect 82634 352563 82690 353363
rect 83738 352563 83794 353363
rect 84750 352563 84806 353363
rect 85854 352563 85910 353363
rect 86866 352563 86922 353363
rect 87970 352563 88026 353363
rect 89074 352563 89130 353363
rect 90086 352563 90142 353363
rect 91190 352563 91246 353363
rect 92294 352563 92350 353363
rect 93306 352563 93362 353363
rect 94410 352563 94466 353363
rect 95422 352563 95478 353363
rect 96526 352563 96582 353363
rect 97630 352563 97686 353363
rect 98642 352563 98698 353363
rect 99746 352563 99802 353363
rect 100758 352563 100814 353363
rect 101862 352563 101918 353363
rect 102966 352563 103022 353363
rect 103978 352563 104034 353363
rect 105082 352563 105138 353363
rect 106094 352563 106150 353363
rect 107198 352563 107254 353363
rect 108302 352563 108358 353363
rect 109314 352563 109370 353363
rect 110418 352563 110474 353363
rect 111430 352563 111486 353363
rect 112534 352563 112590 353363
rect 113638 352563 113694 353363
rect 114650 352563 114706 353363
rect 115754 352563 115810 353363
rect 116766 352563 116822 353363
rect 117870 352563 117926 353363
rect 118974 352563 119030 353363
rect 119986 352563 120042 353363
rect 121090 352563 121146 353363
rect 122102 352563 122158 353363
rect 123206 352563 123262 353363
rect 124310 352563 124366 353363
rect 125322 352563 125378 353363
rect 126426 352563 126482 353363
rect 127438 352563 127494 353363
rect 128542 352563 128598 353363
rect 129646 352563 129702 353363
rect 130658 352563 130714 353363
rect 131762 352563 131818 353363
rect 132866 352563 132922 353363
rect 133878 352563 133934 353363
rect 134982 352563 135038 353363
rect 135994 352563 136050 353363
rect 137098 352563 137154 353363
rect 138202 352563 138258 353363
rect 139214 352563 139270 353363
rect 140318 352563 140374 353363
rect 141330 352563 141386 353363
rect 142434 352563 142490 353363
rect 143538 352563 143594 353363
rect 144550 352563 144606 353363
rect 145654 352563 145710 353363
rect 146666 352563 146722 353363
rect 147770 352563 147826 353363
rect 148874 352563 148930 353363
rect 149886 352563 149942 353363
rect 150990 352563 151046 353363
rect 152002 352563 152058 353363
rect 153106 352563 153162 353363
rect 154210 352563 154266 353363
rect 155222 352563 155278 353363
rect 156326 352563 156382 353363
rect 157338 352563 157394 353363
rect 158442 352563 158498 353363
rect 159546 352563 159602 353363
rect 160558 352563 160614 353363
rect 161662 352563 161718 353363
rect 162674 352563 162730 353363
rect 163778 352563 163834 353363
rect 164882 352563 164938 353363
rect 165894 352563 165950 353363
rect 166998 352563 167054 353363
rect 168010 352563 168066 353363
rect 169114 352563 169170 353363
rect 170218 352563 170274 353363
rect 171230 352563 171286 353363
rect 172334 352563 172390 353363
rect 173346 352563 173402 353363
rect 174450 352563 174506 353363
rect 175554 352563 175610 353363
rect 176566 352563 176622 353363
rect 177670 352563 177726 353363
rect 178774 352563 178830 353363
rect 179786 352563 179842 353363
rect 180890 352563 180946 353363
rect 181902 352563 181958 353363
rect 183006 352563 183062 353363
rect 184110 352563 184166 353363
rect 185122 352563 185178 353363
rect 186226 352563 186282 353363
rect 187238 352563 187294 353363
rect 188342 352563 188398 353363
rect 189446 352563 189502 353363
rect 190458 352563 190514 353363
rect 191562 352563 191618 353363
rect 192574 352563 192630 353363
rect 193678 352563 193734 353363
rect 194782 352563 194838 353363
rect 195794 352563 195850 353363
rect 196898 352563 196954 353363
rect 197910 352563 197966 353363
rect 199014 352563 199070 353363
rect 200118 352563 200174 353363
rect 201130 352563 201186 353363
rect 202234 352563 202290 353363
rect 203246 352563 203302 353363
rect 204350 352563 204406 353363
rect 205454 352563 205510 353363
rect 206466 352563 206522 353363
rect 207570 352563 207626 353363
rect 208582 352563 208638 353363
rect 209686 352563 209742 353363
rect 210790 352563 210846 353363
rect 211802 352563 211858 353363
rect 212906 352563 212962 353363
rect 213918 352563 213974 353363
rect 215022 352563 215078 353363
rect 216126 352563 216182 353363
rect 217138 352563 217194 353363
rect 218242 352563 218298 353363
rect 219254 352563 219310 353363
rect 220358 352563 220414 353363
rect 221462 352563 221518 353363
rect 222474 352563 222530 353363
rect 223578 352563 223634 353363
rect 224682 352563 224738 353363
rect 225694 352563 225750 353363
rect 226798 352563 226854 353363
rect 227810 352563 227866 353363
rect 228914 352563 228970 353363
rect 230018 352563 230074 353363
rect 231030 352563 231086 353363
rect 232134 352563 232190 353363
rect 233146 352563 233202 353363
rect 234250 352563 234306 353363
rect 235354 352563 235410 353363
rect 236366 352563 236422 353363
rect 237470 352563 237526 353363
rect 238482 352563 238538 353363
rect 239586 352563 239642 353363
rect 240690 352563 240746 353363
rect 241702 352563 241758 353363
rect 242806 352563 242862 353363
rect 243818 352563 243874 353363
rect 244922 352563 244978 353363
rect 246026 352563 246082 353363
rect 247038 352563 247094 353363
rect 248142 352563 248198 353363
rect 249154 352563 249210 353363
rect 250258 352563 250314 353363
rect 251362 352563 251418 353363
rect 252374 352563 252430 353363
rect 253478 352563 253534 353363
rect 254490 352563 254546 353363
rect 255594 352563 255650 353363
rect 256698 352563 256754 353363
rect 257710 352563 257766 353363
rect 258814 352563 258870 353363
rect 259826 352563 259882 353363
rect 260930 352563 260986 353363
rect 262034 352563 262090 353363
rect 263046 352563 263102 353363
rect 264150 352563 264206 353363
rect 265254 352563 265310 353363
rect 266266 352563 266322 353363
rect 267370 352563 267426 353363
rect 268382 352563 268438 353363
rect 269486 352563 269542 353363
rect 270590 352563 270646 353363
rect 271602 352563 271658 353363
rect 272706 352563 272762 353363
rect 273718 352563 273774 353363
rect 274822 352563 274878 353363
rect 275926 352563 275982 353363
rect 276938 352563 276994 353363
rect 278042 352563 278098 353363
rect 279054 352563 279110 353363
rect 280158 352563 280214 353363
rect 281262 352563 281318 353363
rect 282274 352563 282330 353363
rect 283378 352563 283434 353363
rect 284390 352563 284446 353363
rect 285494 352563 285550 353363
rect 286598 352563 286654 353363
rect 287610 352563 287666 353363
rect 288714 352563 288770 353363
rect 289726 352563 289782 353363
rect 290830 352563 290886 353363
rect 291934 352563 291990 353363
rect 292946 352563 293002 353363
rect 294050 352563 294106 353363
rect 295062 352563 295118 353363
rect 296166 352563 296222 353363
rect 297270 352563 297326 353363
rect 298282 352563 298338 353363
rect 299386 352563 299442 353363
rect 300398 352563 300454 353363
rect 301502 352563 301558 353363
rect 302606 352563 302662 353363
rect 303618 352563 303674 353363
rect 304722 352563 304778 353363
rect 305734 352563 305790 353363
rect 306838 352563 306894 353363
rect 307942 352563 307998 353363
rect 308954 352563 309010 353363
rect 310058 352563 310114 353363
rect 311162 352563 311218 353363
rect 312174 352563 312230 353363
rect 313278 352563 313334 353363
rect 314290 352563 314346 353363
rect 315394 352563 315450 353363
rect 316498 352563 316554 353363
rect 317510 352563 317566 353363
rect 318614 352563 318670 353363
rect 319626 352563 319682 353363
rect 320730 352563 320786 353363
rect 321834 352563 321890 353363
rect 322846 352563 322902 353363
rect 323950 352563 324006 353363
rect 324962 352563 325018 353363
rect 326066 352563 326122 353363
rect 327170 352563 327226 353363
rect 328182 352563 328238 353363
rect 329286 352563 329342 353363
rect 330298 352563 330354 353363
rect 331402 352563 331458 353363
rect 332506 352563 332562 353363
rect 333518 352563 333574 353363
rect 334622 352563 334678 353363
rect 335634 352563 335690 353363
rect 336738 352563 336794 353363
rect 337842 352563 337898 353363
rect 338854 352563 338910 353363
rect 339958 352563 340014 353363
rect 340970 352563 341026 353363
rect 342074 352563 342130 353363
rect 343178 352563 343234 353363
rect 344190 352563 344246 353363
rect 345294 352563 345350 353363
rect 346306 352563 346362 353363
rect 347410 352563 347466 353363
rect 348514 352563 348570 353363
rect 349526 352563 349582 353363
rect 350630 352563 350686 353363
rect 294 0 350 800
rect 938 0 994 800
rect 1674 0 1730 800
rect 2410 0 2466 800
rect 3054 0 3110 800
rect 3790 0 3846 800
rect 4526 0 4582 800
rect 5262 0 5318 800
rect 5906 0 5962 800
rect 6642 0 6698 800
rect 7378 0 7434 800
rect 8114 0 8170 800
rect 8758 0 8814 800
rect 9494 0 9550 800
rect 10230 0 10286 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12346 0 12402 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 14462 0 14518 800
rect 15198 0 15254 800
rect 15934 0 15990 800
rect 16670 0 16726 800
rect 17314 0 17370 800
rect 18050 0 18106 800
rect 18786 0 18842 800
rect 19522 0 19578 800
rect 20166 0 20222 800
rect 20902 0 20958 800
rect 21638 0 21694 800
rect 22374 0 22430 800
rect 23018 0 23074 800
rect 23754 0 23810 800
rect 24490 0 24546 800
rect 25226 0 25282 800
rect 25870 0 25926 800
rect 26606 0 26662 800
rect 27342 0 27398 800
rect 28078 0 28134 800
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30194 0 30250 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32310 0 32366 800
rect 33046 0 33102 800
rect 33690 0 33746 800
rect 34426 0 34482 800
rect 35162 0 35218 800
rect 35898 0 35954 800
rect 36542 0 36598 800
rect 37278 0 37334 800
rect 38014 0 38070 800
rect 38750 0 38806 800
rect 39394 0 39450 800
rect 40130 0 40186 800
rect 40866 0 40922 800
rect 41602 0 41658 800
rect 42246 0 42302 800
rect 42982 0 43038 800
rect 43718 0 43774 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45834 0 45890 800
rect 46570 0 46626 800
rect 47306 0 47362 800
rect 47950 0 48006 800
rect 48686 0 48742 800
rect 49422 0 49478 800
rect 50158 0 50214 800
rect 50802 0 50858 800
rect 51538 0 51594 800
rect 52274 0 52330 800
rect 53010 0 53066 800
rect 53654 0 53710 800
rect 54390 0 54446 800
rect 55126 0 55182 800
rect 55862 0 55918 800
rect 56506 0 56562 800
rect 57242 0 57298 800
rect 57978 0 58034 800
rect 58714 0 58770 800
rect 59358 0 59414 800
rect 60094 0 60150 800
rect 60830 0 60886 800
rect 61566 0 61622 800
rect 62210 0 62266 800
rect 62946 0 63002 800
rect 63682 0 63738 800
rect 64326 0 64382 800
rect 65062 0 65118 800
rect 65798 0 65854 800
rect 66534 0 66590 800
rect 67178 0 67234 800
rect 67914 0 67970 800
rect 68650 0 68706 800
rect 69386 0 69442 800
rect 70030 0 70086 800
rect 70766 0 70822 800
rect 71502 0 71558 800
rect 72238 0 72294 800
rect 72882 0 72938 800
rect 73618 0 73674 800
rect 74354 0 74410 800
rect 75090 0 75146 800
rect 75734 0 75790 800
rect 76470 0 76526 800
rect 77206 0 77262 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79322 0 79378 800
rect 80058 0 80114 800
rect 80794 0 80850 800
rect 81438 0 81494 800
rect 82174 0 82230 800
rect 82910 0 82966 800
rect 83646 0 83702 800
rect 84290 0 84346 800
rect 85026 0 85082 800
rect 85762 0 85818 800
rect 86498 0 86554 800
rect 87142 0 87198 800
rect 87878 0 87934 800
rect 88614 0 88670 800
rect 89350 0 89406 800
rect 89994 0 90050 800
rect 90730 0 90786 800
rect 91466 0 91522 800
rect 92202 0 92258 800
rect 92846 0 92902 800
rect 93582 0 93638 800
rect 94318 0 94374 800
rect 95054 0 95110 800
rect 95698 0 95754 800
rect 96434 0 96490 800
rect 97170 0 97226 800
rect 97814 0 97870 800
rect 98550 0 98606 800
rect 99286 0 99342 800
rect 100022 0 100078 800
rect 100666 0 100722 800
rect 101402 0 101458 800
rect 102138 0 102194 800
rect 102874 0 102930 800
rect 103518 0 103574 800
rect 104254 0 104310 800
rect 104990 0 105046 800
rect 105726 0 105782 800
rect 106370 0 106426 800
rect 107106 0 107162 800
rect 107842 0 107898 800
rect 108578 0 108634 800
rect 109222 0 109278 800
rect 109958 0 110014 800
rect 110694 0 110750 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 112810 0 112866 800
rect 113546 0 113602 800
rect 114282 0 114338 800
rect 114926 0 114982 800
rect 115662 0 115718 800
rect 116398 0 116454 800
rect 117134 0 117190 800
rect 117778 0 117834 800
rect 118514 0 118570 800
rect 119250 0 119306 800
rect 119986 0 120042 800
rect 120630 0 120686 800
rect 121366 0 121422 800
rect 122102 0 122158 800
rect 122838 0 122894 800
rect 123482 0 123538 800
rect 124218 0 124274 800
rect 124954 0 125010 800
rect 125690 0 125746 800
rect 126334 0 126390 800
rect 127070 0 127126 800
rect 127806 0 127862 800
rect 128450 0 128506 800
rect 129186 0 129242 800
rect 129922 0 129978 800
rect 130658 0 130714 800
rect 131302 0 131358 800
rect 132038 0 132094 800
rect 132774 0 132830 800
rect 133510 0 133566 800
rect 134154 0 134210 800
rect 134890 0 134946 800
rect 135626 0 135682 800
rect 136362 0 136418 800
rect 137006 0 137062 800
rect 137742 0 137798 800
rect 138478 0 138534 800
rect 139214 0 139270 800
rect 139858 0 139914 800
rect 140594 0 140650 800
rect 141330 0 141386 800
rect 142066 0 142122 800
rect 142710 0 142766 800
rect 143446 0 143502 800
rect 144182 0 144238 800
rect 144918 0 144974 800
rect 145562 0 145618 800
rect 146298 0 146354 800
rect 147034 0 147090 800
rect 147770 0 147826 800
rect 148414 0 148470 800
rect 149150 0 149206 800
rect 149886 0 149942 800
rect 150622 0 150678 800
rect 151266 0 151322 800
rect 152002 0 152058 800
rect 152738 0 152794 800
rect 153474 0 153530 800
rect 154118 0 154174 800
rect 154854 0 154910 800
rect 155590 0 155646 800
rect 156326 0 156382 800
rect 156970 0 157026 800
rect 157706 0 157762 800
rect 158442 0 158498 800
rect 159178 0 159234 800
rect 159822 0 159878 800
rect 160558 0 160614 800
rect 161294 0 161350 800
rect 161938 0 161994 800
rect 162674 0 162730 800
rect 163410 0 163466 800
rect 164146 0 164202 800
rect 164790 0 164846 800
rect 165526 0 165582 800
rect 166262 0 166318 800
rect 166998 0 167054 800
rect 167642 0 167698 800
rect 168378 0 168434 800
rect 169114 0 169170 800
rect 169850 0 169906 800
rect 170494 0 170550 800
rect 171230 0 171286 800
rect 171966 0 172022 800
rect 172702 0 172758 800
rect 173346 0 173402 800
rect 174082 0 174138 800
rect 174818 0 174874 800
rect 175554 0 175610 800
rect 176198 0 176254 800
rect 176934 0 176990 800
rect 177670 0 177726 800
rect 178406 0 178462 800
rect 179050 0 179106 800
rect 179786 0 179842 800
rect 180522 0 180578 800
rect 181258 0 181314 800
rect 181902 0 181958 800
rect 182638 0 182694 800
rect 183374 0 183430 800
rect 184110 0 184166 800
rect 184754 0 184810 800
rect 185490 0 185546 800
rect 186226 0 186282 800
rect 186962 0 187018 800
rect 187606 0 187662 800
rect 188342 0 188398 800
rect 189078 0 189134 800
rect 189814 0 189870 800
rect 190458 0 190514 800
rect 191194 0 191250 800
rect 191930 0 191986 800
rect 192574 0 192630 800
rect 193310 0 193366 800
rect 194046 0 194102 800
rect 194782 0 194838 800
rect 195426 0 195482 800
rect 196162 0 196218 800
rect 196898 0 196954 800
rect 197634 0 197690 800
rect 198278 0 198334 800
rect 199014 0 199070 800
rect 199750 0 199806 800
rect 200486 0 200542 800
rect 201130 0 201186 800
rect 201866 0 201922 800
rect 202602 0 202658 800
rect 203338 0 203394 800
rect 203982 0 204038 800
rect 204718 0 204774 800
rect 205454 0 205510 800
rect 206190 0 206246 800
rect 206834 0 206890 800
rect 207570 0 207626 800
rect 208306 0 208362 800
rect 209042 0 209098 800
rect 209686 0 209742 800
rect 210422 0 210478 800
rect 211158 0 211214 800
rect 211894 0 211950 800
rect 212538 0 212594 800
rect 213274 0 213330 800
rect 214010 0 214066 800
rect 214746 0 214802 800
rect 215390 0 215446 800
rect 216126 0 216182 800
rect 216862 0 216918 800
rect 217598 0 217654 800
rect 218242 0 218298 800
rect 218978 0 219034 800
rect 219714 0 219770 800
rect 220450 0 220506 800
rect 221094 0 221150 800
rect 221830 0 221886 800
rect 222566 0 222622 800
rect 223302 0 223358 800
rect 223946 0 224002 800
rect 224682 0 224738 800
rect 225418 0 225474 800
rect 226062 0 226118 800
rect 226798 0 226854 800
rect 227534 0 227590 800
rect 228270 0 228326 800
rect 228914 0 228970 800
rect 229650 0 229706 800
rect 230386 0 230442 800
rect 231122 0 231178 800
rect 231766 0 231822 800
rect 232502 0 232558 800
rect 233238 0 233294 800
rect 233974 0 234030 800
rect 234618 0 234674 800
rect 235354 0 235410 800
rect 236090 0 236146 800
rect 236826 0 236882 800
rect 237470 0 237526 800
rect 238206 0 238262 800
rect 238942 0 238998 800
rect 239678 0 239734 800
rect 240322 0 240378 800
rect 241058 0 241114 800
rect 241794 0 241850 800
rect 242530 0 242586 800
rect 243174 0 243230 800
rect 243910 0 243966 800
rect 244646 0 244702 800
rect 245382 0 245438 800
rect 246026 0 246082 800
rect 246762 0 246818 800
rect 247498 0 247554 800
rect 248234 0 248290 800
rect 248878 0 248934 800
rect 249614 0 249670 800
rect 250350 0 250406 800
rect 251086 0 251142 800
rect 251730 0 251786 800
rect 252466 0 252522 800
rect 253202 0 253258 800
rect 253938 0 253994 800
rect 254582 0 254638 800
rect 255318 0 255374 800
rect 256054 0 256110 800
rect 256698 0 256754 800
rect 257434 0 257490 800
rect 258170 0 258226 800
rect 258906 0 258962 800
rect 259550 0 259606 800
rect 260286 0 260342 800
rect 261022 0 261078 800
rect 261758 0 261814 800
rect 262402 0 262458 800
rect 263138 0 263194 800
rect 263874 0 263930 800
rect 264610 0 264666 800
rect 265254 0 265310 800
rect 265990 0 266046 800
rect 266726 0 266782 800
rect 267462 0 267518 800
rect 268106 0 268162 800
rect 268842 0 268898 800
rect 269578 0 269634 800
rect 270314 0 270370 800
rect 270958 0 271014 800
rect 271694 0 271750 800
rect 272430 0 272486 800
rect 273166 0 273222 800
rect 273810 0 273866 800
rect 274546 0 274602 800
rect 275282 0 275338 800
rect 276018 0 276074 800
rect 276662 0 276718 800
rect 277398 0 277454 800
rect 278134 0 278190 800
rect 278870 0 278926 800
rect 279514 0 279570 800
rect 280250 0 280306 800
rect 280986 0 281042 800
rect 281722 0 281778 800
rect 282366 0 282422 800
rect 283102 0 283158 800
rect 283838 0 283894 800
rect 284574 0 284630 800
rect 285218 0 285274 800
rect 285954 0 286010 800
rect 286690 0 286746 800
rect 287426 0 287482 800
rect 288070 0 288126 800
rect 288806 0 288862 800
rect 289542 0 289598 800
rect 290186 0 290242 800
rect 290922 0 290978 800
rect 291658 0 291714 800
rect 292394 0 292450 800
rect 293038 0 293094 800
rect 293774 0 293830 800
rect 294510 0 294566 800
rect 295246 0 295302 800
rect 295890 0 295946 800
rect 296626 0 296682 800
rect 297362 0 297418 800
rect 298098 0 298154 800
rect 298742 0 298798 800
rect 299478 0 299534 800
rect 300214 0 300270 800
rect 300950 0 301006 800
rect 301594 0 301650 800
rect 302330 0 302386 800
rect 303066 0 303122 800
rect 303802 0 303858 800
rect 304446 0 304502 800
rect 305182 0 305238 800
rect 305918 0 305974 800
rect 306654 0 306710 800
rect 307298 0 307354 800
rect 308034 0 308090 800
rect 308770 0 308826 800
rect 309506 0 309562 800
rect 310150 0 310206 800
rect 310886 0 310942 800
rect 311622 0 311678 800
rect 312358 0 312414 800
rect 313002 0 313058 800
rect 313738 0 313794 800
rect 314474 0 314530 800
rect 315210 0 315266 800
rect 315854 0 315910 800
rect 316590 0 316646 800
rect 317326 0 317382 800
rect 318062 0 318118 800
rect 318706 0 318762 800
rect 319442 0 319498 800
rect 320178 0 320234 800
rect 320822 0 320878 800
rect 321558 0 321614 800
rect 322294 0 322350 800
rect 323030 0 323086 800
rect 323674 0 323730 800
rect 324410 0 324466 800
rect 325146 0 325202 800
rect 325882 0 325938 800
rect 326526 0 326582 800
rect 327262 0 327318 800
rect 327998 0 328054 800
rect 328734 0 328790 800
rect 329378 0 329434 800
rect 330114 0 330170 800
rect 330850 0 330906 800
rect 331586 0 331642 800
rect 332230 0 332286 800
rect 332966 0 333022 800
rect 333702 0 333758 800
rect 334438 0 334494 800
rect 335082 0 335138 800
rect 335818 0 335874 800
rect 336554 0 336610 800
rect 337290 0 337346 800
rect 337934 0 337990 800
rect 338670 0 338726 800
rect 339406 0 339462 800
rect 340142 0 340198 800
rect 340786 0 340842 800
rect 341522 0 341578 800
rect 342258 0 342314 800
rect 342994 0 343050 800
rect 343638 0 343694 800
rect 344374 0 344430 800
rect 345110 0 345166 800
rect 345846 0 345902 800
rect 346490 0 346546 800
rect 347226 0 347282 800
rect 347962 0 348018 800
rect 348698 0 348754 800
rect 349342 0 349398 800
rect 350078 0 350134 800
rect 350814 0 350870 800
<< obsm2 >>
rect 296 352507 422 353161
rect 590 352507 1434 353161
rect 1602 352507 2538 353161
rect 2706 352507 3550 353161
rect 3718 352507 4654 353161
rect 4822 352507 5758 353161
rect 5926 352507 6770 353161
rect 6938 352507 7874 353161
rect 8042 352507 8886 353161
rect 9054 352507 9990 353161
rect 10158 352507 11094 353161
rect 11262 352507 12106 353161
rect 12274 352507 13210 353161
rect 13378 352507 14222 353161
rect 14390 352507 15326 353161
rect 15494 352507 16430 353161
rect 16598 352507 17442 353161
rect 17610 352507 18546 353161
rect 18714 352507 19558 353161
rect 19726 352507 20662 353161
rect 20830 352507 21766 353161
rect 21934 352507 22778 353161
rect 22946 352507 23882 353161
rect 24050 352507 24894 353161
rect 25062 352507 25998 353161
rect 26166 352507 27102 353161
rect 27270 352507 28114 353161
rect 28282 352507 29218 353161
rect 29386 352507 30230 353161
rect 30398 352507 31334 353161
rect 31502 352507 32438 353161
rect 32606 352507 33450 353161
rect 33618 352507 34554 353161
rect 34722 352507 35566 353161
rect 35734 352507 36670 353161
rect 36838 352507 37774 353161
rect 37942 352507 38786 353161
rect 38954 352507 39890 353161
rect 40058 352507 40902 353161
rect 41070 352507 42006 353161
rect 42174 352507 43110 353161
rect 43278 352507 44122 353161
rect 44290 352507 45226 353161
rect 45394 352507 46330 353161
rect 46498 352507 47342 353161
rect 47510 352507 48446 353161
rect 48614 352507 49458 353161
rect 49626 352507 50562 353161
rect 50730 352507 51666 353161
rect 51834 352507 52678 353161
rect 52846 352507 53782 353161
rect 53950 352507 54794 353161
rect 54962 352507 55898 353161
rect 56066 352507 57002 353161
rect 57170 352507 58014 353161
rect 58182 352507 59118 353161
rect 59286 352507 60130 353161
rect 60298 352507 61234 353161
rect 61402 352507 62338 353161
rect 62506 352507 63350 353161
rect 63518 352507 64454 353161
rect 64622 352507 65466 353161
rect 65634 352507 66570 353161
rect 66738 352507 67674 353161
rect 67842 352507 68686 353161
rect 68854 352507 69790 353161
rect 69958 352507 70802 353161
rect 70970 352507 71906 353161
rect 72074 352507 73010 353161
rect 73178 352507 74022 353161
rect 74190 352507 75126 353161
rect 75294 352507 76138 353161
rect 76306 352507 77242 353161
rect 77410 352507 78346 353161
rect 78514 352507 79358 353161
rect 79526 352507 80462 353161
rect 80630 352507 81474 353161
rect 81642 352507 82578 353161
rect 82746 352507 83682 353161
rect 83850 352507 84694 353161
rect 84862 352507 85798 353161
rect 85966 352507 86810 353161
rect 86978 352507 87914 353161
rect 88082 352507 89018 353161
rect 89186 352507 90030 353161
rect 90198 352507 91134 353161
rect 91302 352507 92238 353161
rect 92406 352507 93250 353161
rect 93418 352507 94354 353161
rect 94522 352507 95366 353161
rect 95534 352507 96470 353161
rect 96638 352507 97574 353161
rect 97742 352507 98586 353161
rect 98754 352507 99690 353161
rect 99858 352507 100702 353161
rect 100870 352507 101806 353161
rect 101974 352507 102910 353161
rect 103078 352507 103922 353161
rect 104090 352507 105026 353161
rect 105194 352507 106038 353161
rect 106206 352507 107142 353161
rect 107310 352507 108246 353161
rect 108414 352507 109258 353161
rect 109426 352507 110362 353161
rect 110530 352507 111374 353161
rect 111542 352507 112478 353161
rect 112646 352507 113582 353161
rect 113750 352507 114594 353161
rect 114762 352507 115698 353161
rect 115866 352507 116710 353161
rect 116878 352507 117814 353161
rect 117982 352507 118918 353161
rect 119086 352507 119930 353161
rect 120098 352507 121034 353161
rect 121202 352507 122046 353161
rect 122214 352507 123150 353161
rect 123318 352507 124254 353161
rect 124422 352507 125266 353161
rect 125434 352507 126370 353161
rect 126538 352507 127382 353161
rect 127550 352507 128486 353161
rect 128654 352507 129590 353161
rect 129758 352507 130602 353161
rect 130770 352507 131706 353161
rect 131874 352507 132810 353161
rect 132978 352507 133822 353161
rect 133990 352507 134926 353161
rect 135094 352507 135938 353161
rect 136106 352507 137042 353161
rect 137210 352507 138146 353161
rect 138314 352507 139158 353161
rect 139326 352507 140262 353161
rect 140430 352507 141274 353161
rect 141442 352507 142378 353161
rect 142546 352507 143482 353161
rect 143650 352507 144494 353161
rect 144662 352507 145598 353161
rect 145766 352507 146610 353161
rect 146778 352507 147714 353161
rect 147882 352507 148818 353161
rect 148986 352507 149830 353161
rect 149998 352507 150934 353161
rect 151102 352507 151946 353161
rect 152114 352507 153050 353161
rect 153218 352507 154154 353161
rect 154322 352507 155166 353161
rect 155334 352507 156270 353161
rect 156438 352507 157282 353161
rect 157450 352507 158386 353161
rect 158554 352507 159490 353161
rect 159658 352507 160502 353161
rect 160670 352507 161606 353161
rect 161774 352507 162618 353161
rect 162786 352507 163722 353161
rect 163890 352507 164826 353161
rect 164994 352507 165838 353161
rect 166006 352507 166942 353161
rect 167110 352507 167954 353161
rect 168122 352507 169058 353161
rect 169226 352507 170162 353161
rect 170330 352507 171174 353161
rect 171342 352507 172278 353161
rect 172446 352507 173290 353161
rect 173458 352507 174394 353161
rect 174562 352507 175498 353161
rect 175666 352507 176510 353161
rect 176678 352507 177614 353161
rect 177782 352507 178718 353161
rect 178886 352507 179730 353161
rect 179898 352507 180834 353161
rect 181002 352507 181846 353161
rect 182014 352507 182950 353161
rect 183118 352507 184054 353161
rect 184222 352507 185066 353161
rect 185234 352507 186170 353161
rect 186338 352507 187182 353161
rect 187350 352507 188286 353161
rect 188454 352507 189390 353161
rect 189558 352507 190402 353161
rect 190570 352507 191506 353161
rect 191674 352507 192518 353161
rect 192686 352507 193622 353161
rect 193790 352507 194726 353161
rect 194894 352507 195738 353161
rect 195906 352507 196842 353161
rect 197010 352507 197854 353161
rect 198022 352507 198958 353161
rect 199126 352507 200062 353161
rect 200230 352507 201074 353161
rect 201242 352507 202178 353161
rect 202346 352507 203190 353161
rect 203358 352507 204294 353161
rect 204462 352507 205398 353161
rect 205566 352507 206410 353161
rect 206578 352507 207514 353161
rect 207682 352507 208526 353161
rect 208694 352507 209630 353161
rect 209798 352507 210734 353161
rect 210902 352507 211746 353161
rect 211914 352507 212850 353161
rect 213018 352507 213862 353161
rect 214030 352507 214966 353161
rect 215134 352507 216070 353161
rect 216238 352507 217082 353161
rect 217250 352507 218186 353161
rect 218354 352507 219198 353161
rect 219366 352507 220302 353161
rect 220470 352507 221406 353161
rect 221574 352507 222418 353161
rect 222586 352507 223522 353161
rect 223690 352507 224626 353161
rect 224794 352507 225638 353161
rect 225806 352507 226742 353161
rect 226910 352507 227754 353161
rect 227922 352507 228858 353161
rect 229026 352507 229962 353161
rect 230130 352507 230974 353161
rect 231142 352507 232078 353161
rect 232246 352507 233090 353161
rect 233258 352507 234194 353161
rect 234362 352507 235298 353161
rect 235466 352507 236310 353161
rect 236478 352507 237414 353161
rect 237582 352507 238426 353161
rect 238594 352507 239530 353161
rect 239698 352507 240634 353161
rect 240802 352507 241646 353161
rect 241814 352507 242750 353161
rect 242918 352507 243762 353161
rect 243930 352507 244866 353161
rect 245034 352507 245970 353161
rect 246138 352507 246982 353161
rect 247150 352507 248086 353161
rect 248254 352507 249098 353161
rect 249266 352507 250202 353161
rect 250370 352507 251306 353161
rect 251474 352507 252318 353161
rect 252486 352507 253422 353161
rect 253590 352507 254434 353161
rect 254602 352507 255538 353161
rect 255706 352507 256642 353161
rect 256810 352507 257654 353161
rect 257822 352507 258758 353161
rect 258926 352507 259770 353161
rect 259938 352507 260874 353161
rect 261042 352507 261978 353161
rect 262146 352507 262990 353161
rect 263158 352507 264094 353161
rect 264262 352507 265198 353161
rect 265366 352507 266210 353161
rect 266378 352507 267314 353161
rect 267482 352507 268326 353161
rect 268494 352507 269430 353161
rect 269598 352507 270534 353161
rect 270702 352507 271546 353161
rect 271714 352507 272650 353161
rect 272818 352507 273662 353161
rect 273830 352507 274766 353161
rect 274934 352507 275870 353161
rect 276038 352507 276882 353161
rect 277050 352507 277986 353161
rect 278154 352507 278998 353161
rect 279166 352507 280102 353161
rect 280270 352507 281206 353161
rect 281374 352507 282218 353161
rect 282386 352507 283322 353161
rect 283490 352507 284334 353161
rect 284502 352507 285438 353161
rect 285606 352507 286542 353161
rect 286710 352507 287554 353161
rect 287722 352507 288658 353161
rect 288826 352507 289670 353161
rect 289838 352507 290774 353161
rect 290942 352507 291878 353161
rect 292046 352507 292890 353161
rect 293058 352507 293994 353161
rect 294162 352507 295006 353161
rect 295174 352507 296110 353161
rect 296278 352507 297214 353161
rect 297382 352507 298226 353161
rect 298394 352507 299330 353161
rect 299498 352507 300342 353161
rect 300510 352507 301446 353161
rect 301614 352507 302550 353161
rect 302718 352507 303562 353161
rect 303730 352507 304666 353161
rect 304834 352507 305678 353161
rect 305846 352507 306782 353161
rect 306950 352507 307886 353161
rect 308054 352507 308898 353161
rect 309066 352507 310002 353161
rect 310170 352507 311106 353161
rect 311274 352507 312118 353161
rect 312286 352507 313222 353161
rect 313390 352507 314234 353161
rect 314402 352507 315338 353161
rect 315506 352507 316442 353161
rect 316610 352507 317454 353161
rect 317622 352507 318558 353161
rect 318726 352507 319570 353161
rect 319738 352507 320674 353161
rect 320842 352507 321778 353161
rect 321946 352507 322790 353161
rect 322958 352507 323894 353161
rect 324062 352507 324906 353161
rect 325074 352507 326010 353161
rect 326178 352507 327114 353161
rect 327282 352507 328126 353161
rect 328294 352507 329230 353161
rect 329398 352507 330242 353161
rect 330410 352507 331346 353161
rect 331514 352507 332450 353161
rect 332618 352507 333462 353161
rect 333630 352507 334566 353161
rect 334734 352507 335578 353161
rect 335746 352507 336682 353161
rect 336850 352507 337786 353161
rect 337954 352507 338798 353161
rect 338966 352507 339902 353161
rect 340070 352507 340914 353161
rect 341082 352507 342018 353161
rect 342186 352507 343122 353161
rect 343290 352507 344134 353161
rect 344302 352507 345238 353161
rect 345406 352507 346250 353161
rect 346418 352507 347354 353161
rect 347522 352507 348458 353161
rect 348626 352507 349470 353161
rect 349638 352507 350574 353161
rect 350742 352507 350868 353161
rect 296 856 350868 352507
rect 406 800 882 856
rect 1050 800 1618 856
rect 1786 800 2354 856
rect 2522 800 2998 856
rect 3166 800 3734 856
rect 3902 800 4470 856
rect 4638 800 5206 856
rect 5374 800 5850 856
rect 6018 800 6586 856
rect 6754 800 7322 856
rect 7490 800 8058 856
rect 8226 800 8702 856
rect 8870 800 9438 856
rect 9606 800 10174 856
rect 10342 800 10910 856
rect 11078 800 11554 856
rect 11722 800 12290 856
rect 12458 800 13026 856
rect 13194 800 13762 856
rect 13930 800 14406 856
rect 14574 800 15142 856
rect 15310 800 15878 856
rect 16046 800 16614 856
rect 16782 800 17258 856
rect 17426 800 17994 856
rect 18162 800 18730 856
rect 18898 800 19466 856
rect 19634 800 20110 856
rect 20278 800 20846 856
rect 21014 800 21582 856
rect 21750 800 22318 856
rect 22486 800 22962 856
rect 23130 800 23698 856
rect 23866 800 24434 856
rect 24602 800 25170 856
rect 25338 800 25814 856
rect 25982 800 26550 856
rect 26718 800 27286 856
rect 27454 800 28022 856
rect 28190 800 28666 856
rect 28834 800 29402 856
rect 29570 800 30138 856
rect 30306 800 30874 856
rect 31042 800 31518 856
rect 31686 800 32254 856
rect 32422 800 32990 856
rect 33158 800 33634 856
rect 33802 800 34370 856
rect 34538 800 35106 856
rect 35274 800 35842 856
rect 36010 800 36486 856
rect 36654 800 37222 856
rect 37390 800 37958 856
rect 38126 800 38694 856
rect 38862 800 39338 856
rect 39506 800 40074 856
rect 40242 800 40810 856
rect 40978 800 41546 856
rect 41714 800 42190 856
rect 42358 800 42926 856
rect 43094 800 43662 856
rect 43830 800 44398 856
rect 44566 800 45042 856
rect 45210 800 45778 856
rect 45946 800 46514 856
rect 46682 800 47250 856
rect 47418 800 47894 856
rect 48062 800 48630 856
rect 48798 800 49366 856
rect 49534 800 50102 856
rect 50270 800 50746 856
rect 50914 800 51482 856
rect 51650 800 52218 856
rect 52386 800 52954 856
rect 53122 800 53598 856
rect 53766 800 54334 856
rect 54502 800 55070 856
rect 55238 800 55806 856
rect 55974 800 56450 856
rect 56618 800 57186 856
rect 57354 800 57922 856
rect 58090 800 58658 856
rect 58826 800 59302 856
rect 59470 800 60038 856
rect 60206 800 60774 856
rect 60942 800 61510 856
rect 61678 800 62154 856
rect 62322 800 62890 856
rect 63058 800 63626 856
rect 63794 800 64270 856
rect 64438 800 65006 856
rect 65174 800 65742 856
rect 65910 800 66478 856
rect 66646 800 67122 856
rect 67290 800 67858 856
rect 68026 800 68594 856
rect 68762 800 69330 856
rect 69498 800 69974 856
rect 70142 800 70710 856
rect 70878 800 71446 856
rect 71614 800 72182 856
rect 72350 800 72826 856
rect 72994 800 73562 856
rect 73730 800 74298 856
rect 74466 800 75034 856
rect 75202 800 75678 856
rect 75846 800 76414 856
rect 76582 800 77150 856
rect 77318 800 77886 856
rect 78054 800 78530 856
rect 78698 800 79266 856
rect 79434 800 80002 856
rect 80170 800 80738 856
rect 80906 800 81382 856
rect 81550 800 82118 856
rect 82286 800 82854 856
rect 83022 800 83590 856
rect 83758 800 84234 856
rect 84402 800 84970 856
rect 85138 800 85706 856
rect 85874 800 86442 856
rect 86610 800 87086 856
rect 87254 800 87822 856
rect 87990 800 88558 856
rect 88726 800 89294 856
rect 89462 800 89938 856
rect 90106 800 90674 856
rect 90842 800 91410 856
rect 91578 800 92146 856
rect 92314 800 92790 856
rect 92958 800 93526 856
rect 93694 800 94262 856
rect 94430 800 94998 856
rect 95166 800 95642 856
rect 95810 800 96378 856
rect 96546 800 97114 856
rect 97282 800 97758 856
rect 97926 800 98494 856
rect 98662 800 99230 856
rect 99398 800 99966 856
rect 100134 800 100610 856
rect 100778 800 101346 856
rect 101514 800 102082 856
rect 102250 800 102818 856
rect 102986 800 103462 856
rect 103630 800 104198 856
rect 104366 800 104934 856
rect 105102 800 105670 856
rect 105838 800 106314 856
rect 106482 800 107050 856
rect 107218 800 107786 856
rect 107954 800 108522 856
rect 108690 800 109166 856
rect 109334 800 109902 856
rect 110070 800 110638 856
rect 110806 800 111374 856
rect 111542 800 112018 856
rect 112186 800 112754 856
rect 112922 800 113490 856
rect 113658 800 114226 856
rect 114394 800 114870 856
rect 115038 800 115606 856
rect 115774 800 116342 856
rect 116510 800 117078 856
rect 117246 800 117722 856
rect 117890 800 118458 856
rect 118626 800 119194 856
rect 119362 800 119930 856
rect 120098 800 120574 856
rect 120742 800 121310 856
rect 121478 800 122046 856
rect 122214 800 122782 856
rect 122950 800 123426 856
rect 123594 800 124162 856
rect 124330 800 124898 856
rect 125066 800 125634 856
rect 125802 800 126278 856
rect 126446 800 127014 856
rect 127182 800 127750 856
rect 127918 800 128394 856
rect 128562 800 129130 856
rect 129298 800 129866 856
rect 130034 800 130602 856
rect 130770 800 131246 856
rect 131414 800 131982 856
rect 132150 800 132718 856
rect 132886 800 133454 856
rect 133622 800 134098 856
rect 134266 800 134834 856
rect 135002 800 135570 856
rect 135738 800 136306 856
rect 136474 800 136950 856
rect 137118 800 137686 856
rect 137854 800 138422 856
rect 138590 800 139158 856
rect 139326 800 139802 856
rect 139970 800 140538 856
rect 140706 800 141274 856
rect 141442 800 142010 856
rect 142178 800 142654 856
rect 142822 800 143390 856
rect 143558 800 144126 856
rect 144294 800 144862 856
rect 145030 800 145506 856
rect 145674 800 146242 856
rect 146410 800 146978 856
rect 147146 800 147714 856
rect 147882 800 148358 856
rect 148526 800 149094 856
rect 149262 800 149830 856
rect 149998 800 150566 856
rect 150734 800 151210 856
rect 151378 800 151946 856
rect 152114 800 152682 856
rect 152850 800 153418 856
rect 153586 800 154062 856
rect 154230 800 154798 856
rect 154966 800 155534 856
rect 155702 800 156270 856
rect 156438 800 156914 856
rect 157082 800 157650 856
rect 157818 800 158386 856
rect 158554 800 159122 856
rect 159290 800 159766 856
rect 159934 800 160502 856
rect 160670 800 161238 856
rect 161406 800 161882 856
rect 162050 800 162618 856
rect 162786 800 163354 856
rect 163522 800 164090 856
rect 164258 800 164734 856
rect 164902 800 165470 856
rect 165638 800 166206 856
rect 166374 800 166942 856
rect 167110 800 167586 856
rect 167754 800 168322 856
rect 168490 800 169058 856
rect 169226 800 169794 856
rect 169962 800 170438 856
rect 170606 800 171174 856
rect 171342 800 171910 856
rect 172078 800 172646 856
rect 172814 800 173290 856
rect 173458 800 174026 856
rect 174194 800 174762 856
rect 174930 800 175498 856
rect 175666 800 176142 856
rect 176310 800 176878 856
rect 177046 800 177614 856
rect 177782 800 178350 856
rect 178518 800 178994 856
rect 179162 800 179730 856
rect 179898 800 180466 856
rect 180634 800 181202 856
rect 181370 800 181846 856
rect 182014 800 182582 856
rect 182750 800 183318 856
rect 183486 800 184054 856
rect 184222 800 184698 856
rect 184866 800 185434 856
rect 185602 800 186170 856
rect 186338 800 186906 856
rect 187074 800 187550 856
rect 187718 800 188286 856
rect 188454 800 189022 856
rect 189190 800 189758 856
rect 189926 800 190402 856
rect 190570 800 191138 856
rect 191306 800 191874 856
rect 192042 800 192518 856
rect 192686 800 193254 856
rect 193422 800 193990 856
rect 194158 800 194726 856
rect 194894 800 195370 856
rect 195538 800 196106 856
rect 196274 800 196842 856
rect 197010 800 197578 856
rect 197746 800 198222 856
rect 198390 800 198958 856
rect 199126 800 199694 856
rect 199862 800 200430 856
rect 200598 800 201074 856
rect 201242 800 201810 856
rect 201978 800 202546 856
rect 202714 800 203282 856
rect 203450 800 203926 856
rect 204094 800 204662 856
rect 204830 800 205398 856
rect 205566 800 206134 856
rect 206302 800 206778 856
rect 206946 800 207514 856
rect 207682 800 208250 856
rect 208418 800 208986 856
rect 209154 800 209630 856
rect 209798 800 210366 856
rect 210534 800 211102 856
rect 211270 800 211838 856
rect 212006 800 212482 856
rect 212650 800 213218 856
rect 213386 800 213954 856
rect 214122 800 214690 856
rect 214858 800 215334 856
rect 215502 800 216070 856
rect 216238 800 216806 856
rect 216974 800 217542 856
rect 217710 800 218186 856
rect 218354 800 218922 856
rect 219090 800 219658 856
rect 219826 800 220394 856
rect 220562 800 221038 856
rect 221206 800 221774 856
rect 221942 800 222510 856
rect 222678 800 223246 856
rect 223414 800 223890 856
rect 224058 800 224626 856
rect 224794 800 225362 856
rect 225530 800 226006 856
rect 226174 800 226742 856
rect 226910 800 227478 856
rect 227646 800 228214 856
rect 228382 800 228858 856
rect 229026 800 229594 856
rect 229762 800 230330 856
rect 230498 800 231066 856
rect 231234 800 231710 856
rect 231878 800 232446 856
rect 232614 800 233182 856
rect 233350 800 233918 856
rect 234086 800 234562 856
rect 234730 800 235298 856
rect 235466 800 236034 856
rect 236202 800 236770 856
rect 236938 800 237414 856
rect 237582 800 238150 856
rect 238318 800 238886 856
rect 239054 800 239622 856
rect 239790 800 240266 856
rect 240434 800 241002 856
rect 241170 800 241738 856
rect 241906 800 242474 856
rect 242642 800 243118 856
rect 243286 800 243854 856
rect 244022 800 244590 856
rect 244758 800 245326 856
rect 245494 800 245970 856
rect 246138 800 246706 856
rect 246874 800 247442 856
rect 247610 800 248178 856
rect 248346 800 248822 856
rect 248990 800 249558 856
rect 249726 800 250294 856
rect 250462 800 251030 856
rect 251198 800 251674 856
rect 251842 800 252410 856
rect 252578 800 253146 856
rect 253314 800 253882 856
rect 254050 800 254526 856
rect 254694 800 255262 856
rect 255430 800 255998 856
rect 256166 800 256642 856
rect 256810 800 257378 856
rect 257546 800 258114 856
rect 258282 800 258850 856
rect 259018 800 259494 856
rect 259662 800 260230 856
rect 260398 800 260966 856
rect 261134 800 261702 856
rect 261870 800 262346 856
rect 262514 800 263082 856
rect 263250 800 263818 856
rect 263986 800 264554 856
rect 264722 800 265198 856
rect 265366 800 265934 856
rect 266102 800 266670 856
rect 266838 800 267406 856
rect 267574 800 268050 856
rect 268218 800 268786 856
rect 268954 800 269522 856
rect 269690 800 270258 856
rect 270426 800 270902 856
rect 271070 800 271638 856
rect 271806 800 272374 856
rect 272542 800 273110 856
rect 273278 800 273754 856
rect 273922 800 274490 856
rect 274658 800 275226 856
rect 275394 800 275962 856
rect 276130 800 276606 856
rect 276774 800 277342 856
rect 277510 800 278078 856
rect 278246 800 278814 856
rect 278982 800 279458 856
rect 279626 800 280194 856
rect 280362 800 280930 856
rect 281098 800 281666 856
rect 281834 800 282310 856
rect 282478 800 283046 856
rect 283214 800 283782 856
rect 283950 800 284518 856
rect 284686 800 285162 856
rect 285330 800 285898 856
rect 286066 800 286634 856
rect 286802 800 287370 856
rect 287538 800 288014 856
rect 288182 800 288750 856
rect 288918 800 289486 856
rect 289654 800 290130 856
rect 290298 800 290866 856
rect 291034 800 291602 856
rect 291770 800 292338 856
rect 292506 800 292982 856
rect 293150 800 293718 856
rect 293886 800 294454 856
rect 294622 800 295190 856
rect 295358 800 295834 856
rect 296002 800 296570 856
rect 296738 800 297306 856
rect 297474 800 298042 856
rect 298210 800 298686 856
rect 298854 800 299422 856
rect 299590 800 300158 856
rect 300326 800 300894 856
rect 301062 800 301538 856
rect 301706 800 302274 856
rect 302442 800 303010 856
rect 303178 800 303746 856
rect 303914 800 304390 856
rect 304558 800 305126 856
rect 305294 800 305862 856
rect 306030 800 306598 856
rect 306766 800 307242 856
rect 307410 800 307978 856
rect 308146 800 308714 856
rect 308882 800 309450 856
rect 309618 800 310094 856
rect 310262 800 310830 856
rect 310998 800 311566 856
rect 311734 800 312302 856
rect 312470 800 312946 856
rect 313114 800 313682 856
rect 313850 800 314418 856
rect 314586 800 315154 856
rect 315322 800 315798 856
rect 315966 800 316534 856
rect 316702 800 317270 856
rect 317438 800 318006 856
rect 318174 800 318650 856
rect 318818 800 319386 856
rect 319554 800 320122 856
rect 320290 800 320766 856
rect 320934 800 321502 856
rect 321670 800 322238 856
rect 322406 800 322974 856
rect 323142 800 323618 856
rect 323786 800 324354 856
rect 324522 800 325090 856
rect 325258 800 325826 856
rect 325994 800 326470 856
rect 326638 800 327206 856
rect 327374 800 327942 856
rect 328110 800 328678 856
rect 328846 800 329322 856
rect 329490 800 330058 856
rect 330226 800 330794 856
rect 330962 800 331530 856
rect 331698 800 332174 856
rect 332342 800 332910 856
rect 333078 800 333646 856
rect 333814 800 334382 856
rect 334550 800 335026 856
rect 335194 800 335762 856
rect 335930 800 336498 856
rect 336666 800 337234 856
rect 337402 800 337878 856
rect 338046 800 338614 856
rect 338782 800 339350 856
rect 339518 800 340086 856
rect 340254 800 340730 856
rect 340898 800 341466 856
rect 341634 800 342202 856
rect 342370 800 342938 856
rect 343106 800 343582 856
rect 343750 800 344318 856
rect 344486 800 345054 856
rect 345222 800 345790 856
rect 345958 800 346434 856
rect 346602 800 347170 856
rect 347338 800 347906 856
rect 348074 800 348642 856
rect 348810 800 349286 856
rect 349454 800 350022 856
rect 350190 800 350758 856
<< metal3 >>
rect 0 352384 800 352504
rect 0 350888 800 351008
rect 0 349256 800 349376
rect 0 347760 800 347880
rect 0 346128 800 346248
rect 0 344632 800 344752
rect 0 343000 800 343120
rect 0 341504 800 341624
rect 0 339872 800 339992
rect 0 338376 800 338496
rect 0 336744 800 336864
rect 0 335248 800 335368
rect 0 333616 800 333736
rect 0 332120 800 332240
rect 0 330488 800 330608
rect 0 328992 800 329112
rect 0 327360 800 327480
rect 0 325864 800 325984
rect 0 324232 800 324352
rect 0 322736 800 322856
rect 0 321104 800 321224
rect 0 319608 800 319728
rect 0 317976 800 318096
rect 0 316480 800 316600
rect 0 314848 800 314968
rect 0 313352 800 313472
rect 0 311720 800 311840
rect 0 310224 800 310344
rect 0 308592 800 308712
rect 0 307096 800 307216
rect 0 305464 800 305584
rect 0 303968 800 304088
rect 0 302336 800 302456
rect 0 300840 800 300960
rect 0 299208 800 299328
rect 0 297712 800 297832
rect 0 296080 800 296200
rect 0 294584 800 294704
rect 0 292952 800 293072
rect 0 291456 800 291576
rect 0 289824 800 289944
rect 0 288328 800 288448
rect 0 286696 800 286816
rect 0 285200 800 285320
rect 0 283568 800 283688
rect 0 282072 800 282192
rect 0 280440 800 280560
rect 0 278944 800 279064
rect 0 277312 800 277432
rect 0 275816 800 275936
rect 0 274184 800 274304
rect 0 272688 800 272808
rect 0 271056 800 271176
rect 0 269560 800 269680
rect 0 267928 800 268048
rect 0 266432 800 266552
rect 0 264800 800 264920
rect 0 263304 800 263424
rect 0 261672 800 261792
rect 0 260176 800 260296
rect 0 258544 800 258664
rect 0 257048 800 257168
rect 0 255416 800 255536
rect 0 253920 800 254040
rect 0 252288 800 252408
rect 0 250792 800 250912
rect 0 249160 800 249280
rect 0 247664 800 247784
rect 0 246032 800 246152
rect 0 244536 800 244656
rect 0 242904 800 243024
rect 0 241408 800 241528
rect 0 239776 800 239896
rect 0 238280 800 238400
rect 0 236648 800 236768
rect 0 235152 800 235272
rect 0 233520 800 233640
rect 0 232024 800 232144
rect 0 230392 800 230512
rect 0 228896 800 229016
rect 0 227264 800 227384
rect 0 225768 800 225888
rect 0 224136 800 224256
rect 0 222640 800 222760
rect 0 221008 800 221128
rect 0 219512 800 219632
rect 0 217880 800 218000
rect 0 216384 800 216504
rect 0 214752 800 214872
rect 0 213256 800 213376
rect 0 211624 800 211744
rect 0 210128 800 210248
rect 0 208496 800 208616
rect 0 207000 800 207120
rect 0 205368 800 205488
rect 0 203872 800 203992
rect 0 202240 800 202360
rect 0 200744 800 200864
rect 0 199112 800 199232
rect 0 197616 800 197736
rect 0 195984 800 196104
rect 0 194488 800 194608
rect 0 192856 800 192976
rect 0 191360 800 191480
rect 0 189728 800 189848
rect 0 188232 800 188352
rect 0 186600 800 186720
rect 0 185104 800 185224
rect 0 183472 800 183592
rect 0 181976 800 182096
rect 0 180344 800 180464
rect 0 178848 800 178968
rect 0 177352 800 177472
rect 0 175720 800 175840
rect 0 174224 800 174344
rect 0 172592 800 172712
rect 0 171096 800 171216
rect 0 169464 800 169584
rect 0 167968 800 168088
rect 0 166336 800 166456
rect 0 164840 800 164960
rect 0 163208 800 163328
rect 0 161712 800 161832
rect 0 160080 800 160200
rect 0 158584 800 158704
rect 0 156952 800 157072
rect 0 155456 800 155576
rect 0 153824 800 153944
rect 0 152328 800 152448
rect 0 150696 800 150816
rect 0 149200 800 149320
rect 0 147568 800 147688
rect 0 146072 800 146192
rect 0 144440 800 144560
rect 0 142944 800 143064
rect 0 141312 800 141432
rect 0 139816 800 139936
rect 0 138184 800 138304
rect 0 136688 800 136808
rect 0 135056 800 135176
rect 0 133560 800 133680
rect 0 131928 800 132048
rect 0 130432 800 130552
rect 0 128800 800 128920
rect 0 127304 800 127424
rect 0 125672 800 125792
rect 0 124176 800 124296
rect 0 122544 800 122664
rect 0 121048 800 121168
rect 0 119416 800 119536
rect 0 117920 800 118040
rect 0 116288 800 116408
rect 0 114792 800 114912
rect 0 113160 800 113280
rect 0 111664 800 111784
rect 0 110032 800 110152
rect 0 108536 800 108656
rect 0 106904 800 107024
rect 0 105408 800 105528
rect 0 103776 800 103896
rect 0 102280 800 102400
rect 0 100648 800 100768
rect 0 99152 800 99272
rect 0 97520 800 97640
rect 0 96024 800 96144
rect 0 94392 800 94512
rect 0 92896 800 93016
rect 0 91264 800 91384
rect 0 89768 800 89888
rect 0 88136 800 88256
rect 0 86640 800 86760
rect 0 85008 800 85128
rect 0 83512 800 83632
rect 0 81880 800 82000
rect 0 80384 800 80504
rect 0 78752 800 78872
rect 0 77256 800 77376
rect 0 75624 800 75744
rect 0 74128 800 74248
rect 0 72496 800 72616
rect 0 71000 800 71120
rect 0 69368 800 69488
rect 0 67872 800 67992
rect 0 66240 800 66360
rect 0 64744 800 64864
rect 0 63112 800 63232
rect 0 61616 800 61736
rect 0 59984 800 60104
rect 0 58488 800 58608
rect 0 56856 800 56976
rect 0 55360 800 55480
rect 0 53728 800 53848
rect 0 52232 800 52352
rect 0 50600 800 50720
rect 0 49104 800 49224
rect 0 47472 800 47592
rect 0 45976 800 46096
rect 0 44344 800 44464
rect 0 42848 800 42968
rect 0 41216 800 41336
rect 0 39720 800 39840
rect 0 38088 800 38208
rect 0 36592 800 36712
rect 0 34960 800 35080
rect 0 33464 800 33584
rect 0 31832 800 31952
rect 0 30336 800 30456
rect 0 28704 800 28824
rect 0 27208 800 27328
rect 0 25576 800 25696
rect 0 24080 800 24200
rect 0 22448 800 22568
rect 0 20952 800 21072
rect 0 19320 800 19440
rect 0 17824 800 17944
rect 0 16192 800 16312
rect 0 14696 800 14816
rect 0 13064 800 13184
rect 0 11568 800 11688
rect 0 9936 800 10056
rect 0 8440 800 8560
rect 0 6808 800 6928
rect 0 5312 800 5432
rect 0 3680 800 3800
rect 0 2184 800 2304
rect 0 688 800 808
<< obsm3 >>
rect 606 352584 348391 353157
rect 880 352304 348391 352584
rect 606 351088 348391 352304
rect 880 350808 348391 351088
rect 606 349456 348391 350808
rect 880 349176 348391 349456
rect 606 347960 348391 349176
rect 880 347680 348391 347960
rect 606 346328 348391 347680
rect 880 346048 348391 346328
rect 606 344832 348391 346048
rect 880 344552 348391 344832
rect 606 343200 348391 344552
rect 880 342920 348391 343200
rect 606 341704 348391 342920
rect 880 341424 348391 341704
rect 606 340072 348391 341424
rect 880 339792 348391 340072
rect 606 338576 348391 339792
rect 880 338296 348391 338576
rect 606 336944 348391 338296
rect 880 336664 348391 336944
rect 606 335448 348391 336664
rect 880 335168 348391 335448
rect 606 333816 348391 335168
rect 880 333536 348391 333816
rect 606 332320 348391 333536
rect 880 332040 348391 332320
rect 606 330688 348391 332040
rect 880 330408 348391 330688
rect 606 329192 348391 330408
rect 880 328912 348391 329192
rect 606 327560 348391 328912
rect 880 327280 348391 327560
rect 606 326064 348391 327280
rect 880 325784 348391 326064
rect 606 324432 348391 325784
rect 880 324152 348391 324432
rect 606 322936 348391 324152
rect 880 322656 348391 322936
rect 606 321304 348391 322656
rect 880 321024 348391 321304
rect 606 319808 348391 321024
rect 880 319528 348391 319808
rect 606 318176 348391 319528
rect 880 317896 348391 318176
rect 606 316680 348391 317896
rect 880 316400 348391 316680
rect 606 315048 348391 316400
rect 880 314768 348391 315048
rect 606 313552 348391 314768
rect 880 313272 348391 313552
rect 606 311920 348391 313272
rect 880 311640 348391 311920
rect 606 310424 348391 311640
rect 880 310144 348391 310424
rect 606 308792 348391 310144
rect 880 308512 348391 308792
rect 606 307296 348391 308512
rect 880 307016 348391 307296
rect 606 305664 348391 307016
rect 880 305384 348391 305664
rect 606 304168 348391 305384
rect 880 303888 348391 304168
rect 606 302536 348391 303888
rect 880 302256 348391 302536
rect 606 301040 348391 302256
rect 880 300760 348391 301040
rect 606 299408 348391 300760
rect 880 299128 348391 299408
rect 606 297912 348391 299128
rect 880 297632 348391 297912
rect 606 296280 348391 297632
rect 880 296000 348391 296280
rect 606 294784 348391 296000
rect 880 294504 348391 294784
rect 606 293152 348391 294504
rect 880 292872 348391 293152
rect 606 291656 348391 292872
rect 880 291376 348391 291656
rect 606 290024 348391 291376
rect 880 289744 348391 290024
rect 606 288528 348391 289744
rect 880 288248 348391 288528
rect 606 286896 348391 288248
rect 880 286616 348391 286896
rect 606 285400 348391 286616
rect 880 285120 348391 285400
rect 606 283768 348391 285120
rect 880 283488 348391 283768
rect 606 282272 348391 283488
rect 880 281992 348391 282272
rect 606 280640 348391 281992
rect 880 280360 348391 280640
rect 606 279144 348391 280360
rect 880 278864 348391 279144
rect 606 277512 348391 278864
rect 880 277232 348391 277512
rect 606 276016 348391 277232
rect 880 275736 348391 276016
rect 606 274384 348391 275736
rect 880 274104 348391 274384
rect 606 272888 348391 274104
rect 880 272608 348391 272888
rect 606 271256 348391 272608
rect 880 270976 348391 271256
rect 606 269760 348391 270976
rect 880 269480 348391 269760
rect 606 268128 348391 269480
rect 880 267848 348391 268128
rect 606 266632 348391 267848
rect 880 266352 348391 266632
rect 606 265000 348391 266352
rect 880 264720 348391 265000
rect 606 263504 348391 264720
rect 880 263224 348391 263504
rect 606 261872 348391 263224
rect 880 261592 348391 261872
rect 606 260376 348391 261592
rect 880 260096 348391 260376
rect 606 258744 348391 260096
rect 880 258464 348391 258744
rect 606 257248 348391 258464
rect 880 256968 348391 257248
rect 606 255616 348391 256968
rect 880 255336 348391 255616
rect 606 254120 348391 255336
rect 880 253840 348391 254120
rect 606 252488 348391 253840
rect 880 252208 348391 252488
rect 606 250992 348391 252208
rect 880 250712 348391 250992
rect 606 249360 348391 250712
rect 880 249080 348391 249360
rect 606 247864 348391 249080
rect 880 247584 348391 247864
rect 606 246232 348391 247584
rect 880 245952 348391 246232
rect 606 244736 348391 245952
rect 880 244456 348391 244736
rect 606 243104 348391 244456
rect 880 242824 348391 243104
rect 606 241608 348391 242824
rect 880 241328 348391 241608
rect 606 239976 348391 241328
rect 880 239696 348391 239976
rect 606 238480 348391 239696
rect 880 238200 348391 238480
rect 606 236848 348391 238200
rect 880 236568 348391 236848
rect 606 235352 348391 236568
rect 880 235072 348391 235352
rect 606 233720 348391 235072
rect 880 233440 348391 233720
rect 606 232224 348391 233440
rect 880 231944 348391 232224
rect 606 230592 348391 231944
rect 880 230312 348391 230592
rect 606 229096 348391 230312
rect 880 228816 348391 229096
rect 606 227464 348391 228816
rect 880 227184 348391 227464
rect 606 225968 348391 227184
rect 880 225688 348391 225968
rect 606 224336 348391 225688
rect 880 224056 348391 224336
rect 606 222840 348391 224056
rect 880 222560 348391 222840
rect 606 221208 348391 222560
rect 880 220928 348391 221208
rect 606 219712 348391 220928
rect 880 219432 348391 219712
rect 606 218080 348391 219432
rect 880 217800 348391 218080
rect 606 216584 348391 217800
rect 880 216304 348391 216584
rect 606 214952 348391 216304
rect 880 214672 348391 214952
rect 606 213456 348391 214672
rect 880 213176 348391 213456
rect 606 211824 348391 213176
rect 880 211544 348391 211824
rect 606 210328 348391 211544
rect 880 210048 348391 210328
rect 606 208696 348391 210048
rect 880 208416 348391 208696
rect 606 207200 348391 208416
rect 880 206920 348391 207200
rect 606 205568 348391 206920
rect 880 205288 348391 205568
rect 606 204072 348391 205288
rect 880 203792 348391 204072
rect 606 202440 348391 203792
rect 880 202160 348391 202440
rect 606 200944 348391 202160
rect 880 200664 348391 200944
rect 606 199312 348391 200664
rect 880 199032 348391 199312
rect 606 197816 348391 199032
rect 880 197536 348391 197816
rect 606 196184 348391 197536
rect 880 195904 348391 196184
rect 606 194688 348391 195904
rect 880 194408 348391 194688
rect 606 193056 348391 194408
rect 880 192776 348391 193056
rect 606 191560 348391 192776
rect 880 191280 348391 191560
rect 606 189928 348391 191280
rect 880 189648 348391 189928
rect 606 188432 348391 189648
rect 880 188152 348391 188432
rect 606 186800 348391 188152
rect 880 186520 348391 186800
rect 606 185304 348391 186520
rect 880 185024 348391 185304
rect 606 183672 348391 185024
rect 880 183392 348391 183672
rect 606 182176 348391 183392
rect 880 181896 348391 182176
rect 606 180544 348391 181896
rect 880 180264 348391 180544
rect 606 179048 348391 180264
rect 880 178768 348391 179048
rect 606 177552 348391 178768
rect 880 177272 348391 177552
rect 606 175920 348391 177272
rect 880 175640 348391 175920
rect 606 174424 348391 175640
rect 880 174144 348391 174424
rect 606 172792 348391 174144
rect 880 172512 348391 172792
rect 606 171296 348391 172512
rect 880 171016 348391 171296
rect 606 169664 348391 171016
rect 880 169384 348391 169664
rect 606 168168 348391 169384
rect 880 167888 348391 168168
rect 606 166536 348391 167888
rect 880 166256 348391 166536
rect 606 165040 348391 166256
rect 880 164760 348391 165040
rect 606 163408 348391 164760
rect 880 163128 348391 163408
rect 606 161912 348391 163128
rect 880 161632 348391 161912
rect 606 160280 348391 161632
rect 880 160000 348391 160280
rect 606 158784 348391 160000
rect 880 158504 348391 158784
rect 606 157152 348391 158504
rect 880 156872 348391 157152
rect 606 155656 348391 156872
rect 880 155376 348391 155656
rect 606 154024 348391 155376
rect 880 153744 348391 154024
rect 606 152528 348391 153744
rect 880 152248 348391 152528
rect 606 150896 348391 152248
rect 880 150616 348391 150896
rect 606 149400 348391 150616
rect 880 149120 348391 149400
rect 606 147768 348391 149120
rect 880 147488 348391 147768
rect 606 146272 348391 147488
rect 880 145992 348391 146272
rect 606 144640 348391 145992
rect 880 144360 348391 144640
rect 606 143144 348391 144360
rect 880 142864 348391 143144
rect 606 141512 348391 142864
rect 880 141232 348391 141512
rect 606 140016 348391 141232
rect 880 139736 348391 140016
rect 606 138384 348391 139736
rect 880 138104 348391 138384
rect 606 136888 348391 138104
rect 880 136608 348391 136888
rect 606 135256 348391 136608
rect 880 134976 348391 135256
rect 606 133760 348391 134976
rect 880 133480 348391 133760
rect 606 132128 348391 133480
rect 880 131848 348391 132128
rect 606 130632 348391 131848
rect 880 130352 348391 130632
rect 606 129000 348391 130352
rect 880 128720 348391 129000
rect 606 127504 348391 128720
rect 880 127224 348391 127504
rect 606 125872 348391 127224
rect 880 125592 348391 125872
rect 606 124376 348391 125592
rect 880 124096 348391 124376
rect 606 122744 348391 124096
rect 880 122464 348391 122744
rect 606 121248 348391 122464
rect 880 120968 348391 121248
rect 606 119616 348391 120968
rect 880 119336 348391 119616
rect 606 118120 348391 119336
rect 880 117840 348391 118120
rect 606 116488 348391 117840
rect 880 116208 348391 116488
rect 606 114992 348391 116208
rect 880 114712 348391 114992
rect 606 113360 348391 114712
rect 880 113080 348391 113360
rect 606 111864 348391 113080
rect 880 111584 348391 111864
rect 606 110232 348391 111584
rect 880 109952 348391 110232
rect 606 108736 348391 109952
rect 880 108456 348391 108736
rect 606 107104 348391 108456
rect 880 106824 348391 107104
rect 606 105608 348391 106824
rect 880 105328 348391 105608
rect 606 103976 348391 105328
rect 880 103696 348391 103976
rect 606 102480 348391 103696
rect 880 102200 348391 102480
rect 606 100848 348391 102200
rect 880 100568 348391 100848
rect 606 99352 348391 100568
rect 880 99072 348391 99352
rect 606 97720 348391 99072
rect 880 97440 348391 97720
rect 606 96224 348391 97440
rect 880 95944 348391 96224
rect 606 94592 348391 95944
rect 880 94312 348391 94592
rect 606 93096 348391 94312
rect 880 92816 348391 93096
rect 606 91464 348391 92816
rect 880 91184 348391 91464
rect 606 89968 348391 91184
rect 880 89688 348391 89968
rect 606 88336 348391 89688
rect 880 88056 348391 88336
rect 606 86840 348391 88056
rect 880 86560 348391 86840
rect 606 85208 348391 86560
rect 880 84928 348391 85208
rect 606 83712 348391 84928
rect 880 83432 348391 83712
rect 606 82080 348391 83432
rect 880 81800 348391 82080
rect 606 80584 348391 81800
rect 880 80304 348391 80584
rect 606 78952 348391 80304
rect 880 78672 348391 78952
rect 606 77456 348391 78672
rect 880 77176 348391 77456
rect 606 75824 348391 77176
rect 880 75544 348391 75824
rect 606 74328 348391 75544
rect 880 74048 348391 74328
rect 606 72696 348391 74048
rect 880 72416 348391 72696
rect 606 71200 348391 72416
rect 880 70920 348391 71200
rect 606 69568 348391 70920
rect 880 69288 348391 69568
rect 606 68072 348391 69288
rect 880 67792 348391 68072
rect 606 66440 348391 67792
rect 880 66160 348391 66440
rect 606 64944 348391 66160
rect 880 64664 348391 64944
rect 606 63312 348391 64664
rect 880 63032 348391 63312
rect 606 61816 348391 63032
rect 880 61536 348391 61816
rect 606 60184 348391 61536
rect 880 59904 348391 60184
rect 606 58688 348391 59904
rect 880 58408 348391 58688
rect 606 57056 348391 58408
rect 880 56776 348391 57056
rect 606 55560 348391 56776
rect 880 55280 348391 55560
rect 606 53928 348391 55280
rect 880 53648 348391 53928
rect 606 52432 348391 53648
rect 880 52152 348391 52432
rect 606 50800 348391 52152
rect 880 50520 348391 50800
rect 606 49304 348391 50520
rect 880 49024 348391 49304
rect 606 47672 348391 49024
rect 880 47392 348391 47672
rect 606 46176 348391 47392
rect 880 45896 348391 46176
rect 606 44544 348391 45896
rect 880 44264 348391 44544
rect 606 43048 348391 44264
rect 880 42768 348391 43048
rect 606 41416 348391 42768
rect 880 41136 348391 41416
rect 606 39920 348391 41136
rect 880 39640 348391 39920
rect 606 38288 348391 39640
rect 880 38008 348391 38288
rect 606 36792 348391 38008
rect 880 36512 348391 36792
rect 606 35160 348391 36512
rect 880 34880 348391 35160
rect 606 33664 348391 34880
rect 880 33384 348391 33664
rect 606 32032 348391 33384
rect 880 31752 348391 32032
rect 606 30536 348391 31752
rect 880 30256 348391 30536
rect 606 28904 348391 30256
rect 880 28624 348391 28904
rect 606 27408 348391 28624
rect 880 27128 348391 27408
rect 606 25776 348391 27128
rect 880 25496 348391 25776
rect 606 24280 348391 25496
rect 880 24000 348391 24280
rect 606 22648 348391 24000
rect 880 22368 348391 22648
rect 606 21152 348391 22368
rect 880 20872 348391 21152
rect 606 19520 348391 20872
rect 880 19240 348391 19520
rect 606 18024 348391 19240
rect 880 17744 348391 18024
rect 606 16392 348391 17744
rect 880 16112 348391 16392
rect 606 14896 348391 16112
rect 880 14616 348391 14896
rect 606 13264 348391 14616
rect 880 12984 348391 13264
rect 606 11768 348391 12984
rect 880 11488 348391 11768
rect 606 10136 348391 11488
rect 880 9856 348391 10136
rect 606 8640 348391 9856
rect 880 8360 348391 8640
rect 606 7008 348391 8360
rect 880 6728 348391 7008
rect 606 5512 348391 6728
rect 880 5232 348391 5512
rect 606 3880 348391 5232
rect 880 3600 348391 3880
rect 606 2384 348391 3600
rect 880 2104 348391 2384
rect 606 888 348391 2104
rect 880 718 348391 888
<< metal4 >>
rect 4208 2128 4528 350928
rect 19568 2128 19888 350928
rect 34928 2128 35248 350928
rect 50288 2128 50608 350928
rect 65648 2128 65968 350928
rect 81008 2128 81328 350928
rect 96368 2128 96688 350928
rect 111728 2128 112048 350928
rect 127088 2128 127408 350928
rect 142448 2128 142768 350928
rect 157808 2128 158128 350928
rect 173168 2128 173488 350928
rect 188528 2128 188848 350928
rect 203888 2128 204208 350928
rect 219248 2128 219568 350928
rect 234608 2128 234928 350928
rect 249968 2128 250288 350928
rect 265328 2128 265648 350928
rect 280688 2128 281008 350928
rect 296048 2128 296368 350928
rect 311408 2128 311728 350928
rect 326768 2128 327088 350928
rect 342128 2128 342448 350928
<< obsm4 >>
rect 611 351008 344573 353157
rect 611 2048 4128 351008
rect 4608 2048 19488 351008
rect 19968 2048 34848 351008
rect 35328 2048 50208 351008
rect 50688 2048 65568 351008
rect 66048 2048 80928 351008
rect 81408 2048 96288 351008
rect 96768 2048 111648 351008
rect 112128 2048 127008 351008
rect 127488 2048 142368 351008
rect 142848 2048 157728 351008
rect 158208 2048 173088 351008
rect 173568 2048 188448 351008
rect 188928 2048 203808 351008
rect 204288 2048 219168 351008
rect 219648 2048 234528 351008
rect 235008 2048 249888 351008
rect 250368 2048 265248 351008
rect 265728 2048 280608 351008
rect 281088 2048 295968 351008
rect 296448 2048 311328 351008
rect 311808 2048 326688 351008
rect 327168 2048 342048 351008
rect 342528 2048 344573 351008
rect 611 1667 344573 2048
<< labels >>
rlabel metal3 s 0 239776 800 239896 6 data_arrays_0_0_ext_ram_addr1[0]
port 1 nsew signal output
rlabel metal3 s 0 241408 800 241528 6 data_arrays_0_0_ext_ram_addr1[1]
port 2 nsew signal output
rlabel metal3 s 0 242904 800 243024 6 data_arrays_0_0_ext_ram_addr1[2]
port 3 nsew signal output
rlabel metal3 s 0 244536 800 244656 6 data_arrays_0_0_ext_ram_addr1[3]
port 4 nsew signal output
rlabel metal3 s 0 246032 800 246152 6 data_arrays_0_0_ext_ram_addr1[4]
port 5 nsew signal output
rlabel metal3 s 0 247664 800 247784 6 data_arrays_0_0_ext_ram_addr1[5]
port 6 nsew signal output
rlabel metal3 s 0 249160 800 249280 6 data_arrays_0_0_ext_ram_addr1[6]
port 7 nsew signal output
rlabel metal3 s 0 250792 800 250912 6 data_arrays_0_0_ext_ram_addr1[7]
port 8 nsew signal output
rlabel metal3 s 0 252288 800 252408 6 data_arrays_0_0_ext_ram_addr1[8]
port 9 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 data_arrays_0_0_ext_ram_addr[0]
port 10 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 data_arrays_0_0_ext_ram_addr[1]
port 11 nsew signal output
rlabel metal3 s 0 103776 800 103896 6 data_arrays_0_0_ext_ram_addr[2]
port 12 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 data_arrays_0_0_ext_ram_addr[3]
port 13 nsew signal output
rlabel metal3 s 0 106904 800 107024 6 data_arrays_0_0_ext_ram_addr[4]
port 14 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 data_arrays_0_0_ext_ram_addr[5]
port 15 nsew signal output
rlabel metal3 s 0 110032 800 110152 6 data_arrays_0_0_ext_ram_addr[6]
port 16 nsew signal output
rlabel metal3 s 0 111664 800 111784 6 data_arrays_0_0_ext_ram_addr[7]
port 17 nsew signal output
rlabel metal3 s 0 113160 800 113280 6 data_arrays_0_0_ext_ram_addr[8]
port 18 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 data_arrays_0_0_ext_ram_clk
port 19 nsew signal output
rlabel metal3 s 0 227264 800 227384 6 data_arrays_0_0_ext_ram_csb1[0]
port 20 nsew signal output
rlabel metal3 s 0 228896 800 229016 6 data_arrays_0_0_ext_ram_csb1[1]
port 21 nsew signal output
rlabel metal3 s 0 230392 800 230512 6 data_arrays_0_0_ext_ram_csb1[2]
port 22 nsew signal output
rlabel metal3 s 0 232024 800 232144 6 data_arrays_0_0_ext_ram_csb1[3]
port 23 nsew signal output
rlabel metal3 s 0 233520 800 233640 6 data_arrays_0_0_ext_ram_csb1[4]
port 24 nsew signal output
rlabel metal3 s 0 235152 800 235272 6 data_arrays_0_0_ext_ram_csb1[5]
port 25 nsew signal output
rlabel metal3 s 0 236648 800 236768 6 data_arrays_0_0_ext_ram_csb1[6]
port 26 nsew signal output
rlabel metal3 s 0 238280 800 238400 6 data_arrays_0_0_ext_ram_csb1[7]
port 27 nsew signal output
rlabel metal3 s 0 219512 800 219632 6 data_arrays_0_0_ext_ram_csb[0]
port 28 nsew signal output
rlabel metal3 s 0 221008 800 221128 6 data_arrays_0_0_ext_ram_csb[1]
port 29 nsew signal output
rlabel metal3 s 0 222640 800 222760 6 data_arrays_0_0_ext_ram_csb[2]
port 30 nsew signal output
rlabel metal3 s 0 224136 800 224256 6 data_arrays_0_0_ext_ram_csb[3]
port 31 nsew signal output
rlabel metal3 s 0 688 800 808 6 data_arrays_0_0_ext_ram_rdata0[0]
port 32 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 data_arrays_0_0_ext_ram_rdata0[10]
port 33 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 data_arrays_0_0_ext_ram_rdata0[11]
port 34 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 data_arrays_0_0_ext_ram_rdata0[12]
port 35 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 data_arrays_0_0_ext_ram_rdata0[13]
port 36 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 data_arrays_0_0_ext_ram_rdata0[14]
port 37 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 data_arrays_0_0_ext_ram_rdata0[15]
port 38 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 data_arrays_0_0_ext_ram_rdata0[16]
port 39 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 data_arrays_0_0_ext_ram_rdata0[17]
port 40 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 data_arrays_0_0_ext_ram_rdata0[18]
port 41 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 data_arrays_0_0_ext_ram_rdata0[19]
port 42 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 data_arrays_0_0_ext_ram_rdata0[1]
port 43 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 data_arrays_0_0_ext_ram_rdata0[20]
port 44 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 data_arrays_0_0_ext_ram_rdata0[21]
port 45 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 data_arrays_0_0_ext_ram_rdata0[22]
port 46 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 data_arrays_0_0_ext_ram_rdata0[23]
port 47 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 data_arrays_0_0_ext_ram_rdata0[24]
port 48 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 data_arrays_0_0_ext_ram_rdata0[25]
port 49 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 data_arrays_0_0_ext_ram_rdata0[26]
port 50 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 data_arrays_0_0_ext_ram_rdata0[27]
port 51 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 data_arrays_0_0_ext_ram_rdata0[28]
port 52 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 data_arrays_0_0_ext_ram_rdata0[29]
port 53 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 data_arrays_0_0_ext_ram_rdata0[2]
port 54 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 data_arrays_0_0_ext_ram_rdata0[30]
port 55 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 data_arrays_0_0_ext_ram_rdata0[31]
port 56 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 data_arrays_0_0_ext_ram_rdata0[32]
port 57 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 data_arrays_0_0_ext_ram_rdata0[33]
port 58 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 data_arrays_0_0_ext_ram_rdata0[34]
port 59 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 data_arrays_0_0_ext_ram_rdata0[35]
port 60 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 data_arrays_0_0_ext_ram_rdata0[36]
port 61 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 data_arrays_0_0_ext_ram_rdata0[37]
port 62 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 data_arrays_0_0_ext_ram_rdata0[38]
port 63 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 data_arrays_0_0_ext_ram_rdata0[39]
port 64 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 data_arrays_0_0_ext_ram_rdata0[3]
port 65 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 data_arrays_0_0_ext_ram_rdata0[40]
port 66 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 data_arrays_0_0_ext_ram_rdata0[41]
port 67 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 data_arrays_0_0_ext_ram_rdata0[42]
port 68 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 data_arrays_0_0_ext_ram_rdata0[43]
port 69 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 data_arrays_0_0_ext_ram_rdata0[44]
port 70 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 data_arrays_0_0_ext_ram_rdata0[45]
port 71 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 data_arrays_0_0_ext_ram_rdata0[46]
port 72 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 data_arrays_0_0_ext_ram_rdata0[47]
port 73 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 data_arrays_0_0_ext_ram_rdata0[48]
port 74 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 data_arrays_0_0_ext_ram_rdata0[49]
port 75 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 data_arrays_0_0_ext_ram_rdata0[4]
port 76 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 data_arrays_0_0_ext_ram_rdata0[50]
port 77 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 data_arrays_0_0_ext_ram_rdata0[51]
port 78 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 data_arrays_0_0_ext_ram_rdata0[52]
port 79 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 data_arrays_0_0_ext_ram_rdata0[53]
port 80 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 data_arrays_0_0_ext_ram_rdata0[54]
port 81 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 data_arrays_0_0_ext_ram_rdata0[55]
port 82 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 data_arrays_0_0_ext_ram_rdata0[56]
port 83 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 data_arrays_0_0_ext_ram_rdata0[57]
port 84 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 data_arrays_0_0_ext_ram_rdata0[58]
port 85 nsew signal input
rlabel metal3 s 0 92896 800 93016 6 data_arrays_0_0_ext_ram_rdata0[59]
port 86 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 data_arrays_0_0_ext_ram_rdata0[5]
port 87 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 data_arrays_0_0_ext_ram_rdata0[60]
port 88 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 data_arrays_0_0_ext_ram_rdata0[61]
port 89 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 data_arrays_0_0_ext_ram_rdata0[62]
port 90 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 data_arrays_0_0_ext_ram_rdata0[63]
port 91 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 data_arrays_0_0_ext_ram_rdata0[6]
port 92 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 data_arrays_0_0_ext_ram_rdata0[7]
port 93 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 data_arrays_0_0_ext_ram_rdata0[8]
port 94 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 data_arrays_0_0_ext_ram_rdata0[9]
port 95 nsew signal input
rlabel metal3 s 0 253920 800 254040 6 data_arrays_0_0_ext_ram_rdata1[0]
port 96 nsew signal input
rlabel metal3 s 0 269560 800 269680 6 data_arrays_0_0_ext_ram_rdata1[10]
port 97 nsew signal input
rlabel metal3 s 0 271056 800 271176 6 data_arrays_0_0_ext_ram_rdata1[11]
port 98 nsew signal input
rlabel metal3 s 0 272688 800 272808 6 data_arrays_0_0_ext_ram_rdata1[12]
port 99 nsew signal input
rlabel metal3 s 0 274184 800 274304 6 data_arrays_0_0_ext_ram_rdata1[13]
port 100 nsew signal input
rlabel metal3 s 0 275816 800 275936 6 data_arrays_0_0_ext_ram_rdata1[14]
port 101 nsew signal input
rlabel metal3 s 0 277312 800 277432 6 data_arrays_0_0_ext_ram_rdata1[15]
port 102 nsew signal input
rlabel metal3 s 0 278944 800 279064 6 data_arrays_0_0_ext_ram_rdata1[16]
port 103 nsew signal input
rlabel metal3 s 0 280440 800 280560 6 data_arrays_0_0_ext_ram_rdata1[17]
port 104 nsew signal input
rlabel metal3 s 0 282072 800 282192 6 data_arrays_0_0_ext_ram_rdata1[18]
port 105 nsew signal input
rlabel metal3 s 0 283568 800 283688 6 data_arrays_0_0_ext_ram_rdata1[19]
port 106 nsew signal input
rlabel metal3 s 0 255416 800 255536 6 data_arrays_0_0_ext_ram_rdata1[1]
port 107 nsew signal input
rlabel metal3 s 0 285200 800 285320 6 data_arrays_0_0_ext_ram_rdata1[20]
port 108 nsew signal input
rlabel metal3 s 0 286696 800 286816 6 data_arrays_0_0_ext_ram_rdata1[21]
port 109 nsew signal input
rlabel metal3 s 0 288328 800 288448 6 data_arrays_0_0_ext_ram_rdata1[22]
port 110 nsew signal input
rlabel metal3 s 0 289824 800 289944 6 data_arrays_0_0_ext_ram_rdata1[23]
port 111 nsew signal input
rlabel metal3 s 0 291456 800 291576 6 data_arrays_0_0_ext_ram_rdata1[24]
port 112 nsew signal input
rlabel metal3 s 0 292952 800 293072 6 data_arrays_0_0_ext_ram_rdata1[25]
port 113 nsew signal input
rlabel metal3 s 0 294584 800 294704 6 data_arrays_0_0_ext_ram_rdata1[26]
port 114 nsew signal input
rlabel metal3 s 0 296080 800 296200 6 data_arrays_0_0_ext_ram_rdata1[27]
port 115 nsew signal input
rlabel metal3 s 0 297712 800 297832 6 data_arrays_0_0_ext_ram_rdata1[28]
port 116 nsew signal input
rlabel metal3 s 0 299208 800 299328 6 data_arrays_0_0_ext_ram_rdata1[29]
port 117 nsew signal input
rlabel metal3 s 0 257048 800 257168 6 data_arrays_0_0_ext_ram_rdata1[2]
port 118 nsew signal input
rlabel metal3 s 0 300840 800 300960 6 data_arrays_0_0_ext_ram_rdata1[30]
port 119 nsew signal input
rlabel metal3 s 0 302336 800 302456 6 data_arrays_0_0_ext_ram_rdata1[31]
port 120 nsew signal input
rlabel metal3 s 0 303968 800 304088 6 data_arrays_0_0_ext_ram_rdata1[32]
port 121 nsew signal input
rlabel metal3 s 0 305464 800 305584 6 data_arrays_0_0_ext_ram_rdata1[33]
port 122 nsew signal input
rlabel metal3 s 0 307096 800 307216 6 data_arrays_0_0_ext_ram_rdata1[34]
port 123 nsew signal input
rlabel metal3 s 0 308592 800 308712 6 data_arrays_0_0_ext_ram_rdata1[35]
port 124 nsew signal input
rlabel metal3 s 0 310224 800 310344 6 data_arrays_0_0_ext_ram_rdata1[36]
port 125 nsew signal input
rlabel metal3 s 0 311720 800 311840 6 data_arrays_0_0_ext_ram_rdata1[37]
port 126 nsew signal input
rlabel metal3 s 0 313352 800 313472 6 data_arrays_0_0_ext_ram_rdata1[38]
port 127 nsew signal input
rlabel metal3 s 0 314848 800 314968 6 data_arrays_0_0_ext_ram_rdata1[39]
port 128 nsew signal input
rlabel metal3 s 0 258544 800 258664 6 data_arrays_0_0_ext_ram_rdata1[3]
port 129 nsew signal input
rlabel metal3 s 0 316480 800 316600 6 data_arrays_0_0_ext_ram_rdata1[40]
port 130 nsew signal input
rlabel metal3 s 0 317976 800 318096 6 data_arrays_0_0_ext_ram_rdata1[41]
port 131 nsew signal input
rlabel metal3 s 0 319608 800 319728 6 data_arrays_0_0_ext_ram_rdata1[42]
port 132 nsew signal input
rlabel metal3 s 0 321104 800 321224 6 data_arrays_0_0_ext_ram_rdata1[43]
port 133 nsew signal input
rlabel metal3 s 0 322736 800 322856 6 data_arrays_0_0_ext_ram_rdata1[44]
port 134 nsew signal input
rlabel metal3 s 0 324232 800 324352 6 data_arrays_0_0_ext_ram_rdata1[45]
port 135 nsew signal input
rlabel metal3 s 0 325864 800 325984 6 data_arrays_0_0_ext_ram_rdata1[46]
port 136 nsew signal input
rlabel metal3 s 0 327360 800 327480 6 data_arrays_0_0_ext_ram_rdata1[47]
port 137 nsew signal input
rlabel metal3 s 0 328992 800 329112 6 data_arrays_0_0_ext_ram_rdata1[48]
port 138 nsew signal input
rlabel metal3 s 0 330488 800 330608 6 data_arrays_0_0_ext_ram_rdata1[49]
port 139 nsew signal input
rlabel metal3 s 0 260176 800 260296 6 data_arrays_0_0_ext_ram_rdata1[4]
port 140 nsew signal input
rlabel metal3 s 0 332120 800 332240 6 data_arrays_0_0_ext_ram_rdata1[50]
port 141 nsew signal input
rlabel metal3 s 0 333616 800 333736 6 data_arrays_0_0_ext_ram_rdata1[51]
port 142 nsew signal input
rlabel metal3 s 0 335248 800 335368 6 data_arrays_0_0_ext_ram_rdata1[52]
port 143 nsew signal input
rlabel metal3 s 0 336744 800 336864 6 data_arrays_0_0_ext_ram_rdata1[53]
port 144 nsew signal input
rlabel metal3 s 0 338376 800 338496 6 data_arrays_0_0_ext_ram_rdata1[54]
port 145 nsew signal input
rlabel metal3 s 0 339872 800 339992 6 data_arrays_0_0_ext_ram_rdata1[55]
port 146 nsew signal input
rlabel metal3 s 0 341504 800 341624 6 data_arrays_0_0_ext_ram_rdata1[56]
port 147 nsew signal input
rlabel metal3 s 0 343000 800 343120 6 data_arrays_0_0_ext_ram_rdata1[57]
port 148 nsew signal input
rlabel metal3 s 0 344632 800 344752 6 data_arrays_0_0_ext_ram_rdata1[58]
port 149 nsew signal input
rlabel metal3 s 0 346128 800 346248 6 data_arrays_0_0_ext_ram_rdata1[59]
port 150 nsew signal input
rlabel metal3 s 0 261672 800 261792 6 data_arrays_0_0_ext_ram_rdata1[5]
port 151 nsew signal input
rlabel metal3 s 0 347760 800 347880 6 data_arrays_0_0_ext_ram_rdata1[60]
port 152 nsew signal input
rlabel metal3 s 0 349256 800 349376 6 data_arrays_0_0_ext_ram_rdata1[61]
port 153 nsew signal input
rlabel metal3 s 0 350888 800 351008 6 data_arrays_0_0_ext_ram_rdata1[62]
port 154 nsew signal input
rlabel metal3 s 0 352384 800 352504 6 data_arrays_0_0_ext_ram_rdata1[63]
port 155 nsew signal input
rlabel metal3 s 0 263304 800 263424 6 data_arrays_0_0_ext_ram_rdata1[6]
port 156 nsew signal input
rlabel metal3 s 0 264800 800 264920 6 data_arrays_0_0_ext_ram_rdata1[7]
port 157 nsew signal input
rlabel metal3 s 0 266432 800 266552 6 data_arrays_0_0_ext_ram_rdata1[8]
port 158 nsew signal input
rlabel metal3 s 0 267928 800 268048 6 data_arrays_0_0_ext_ram_rdata1[9]
port 159 nsew signal input
rlabel metal2 s 283378 352563 283434 353363 6 data_arrays_0_0_ext_ram_rdata2[0]
port 160 nsew signal input
rlabel metal2 s 294050 352563 294106 353363 6 data_arrays_0_0_ext_ram_rdata2[10]
port 161 nsew signal input
rlabel metal2 s 295062 352563 295118 353363 6 data_arrays_0_0_ext_ram_rdata2[11]
port 162 nsew signal input
rlabel metal2 s 296166 352563 296222 353363 6 data_arrays_0_0_ext_ram_rdata2[12]
port 163 nsew signal input
rlabel metal2 s 297270 352563 297326 353363 6 data_arrays_0_0_ext_ram_rdata2[13]
port 164 nsew signal input
rlabel metal2 s 298282 352563 298338 353363 6 data_arrays_0_0_ext_ram_rdata2[14]
port 165 nsew signal input
rlabel metal2 s 299386 352563 299442 353363 6 data_arrays_0_0_ext_ram_rdata2[15]
port 166 nsew signal input
rlabel metal2 s 300398 352563 300454 353363 6 data_arrays_0_0_ext_ram_rdata2[16]
port 167 nsew signal input
rlabel metal2 s 301502 352563 301558 353363 6 data_arrays_0_0_ext_ram_rdata2[17]
port 168 nsew signal input
rlabel metal2 s 302606 352563 302662 353363 6 data_arrays_0_0_ext_ram_rdata2[18]
port 169 nsew signal input
rlabel metal2 s 303618 352563 303674 353363 6 data_arrays_0_0_ext_ram_rdata2[19]
port 170 nsew signal input
rlabel metal2 s 284390 352563 284446 353363 6 data_arrays_0_0_ext_ram_rdata2[1]
port 171 nsew signal input
rlabel metal2 s 304722 352563 304778 353363 6 data_arrays_0_0_ext_ram_rdata2[20]
port 172 nsew signal input
rlabel metal2 s 305734 352563 305790 353363 6 data_arrays_0_0_ext_ram_rdata2[21]
port 173 nsew signal input
rlabel metal2 s 306838 352563 306894 353363 6 data_arrays_0_0_ext_ram_rdata2[22]
port 174 nsew signal input
rlabel metal2 s 307942 352563 307998 353363 6 data_arrays_0_0_ext_ram_rdata2[23]
port 175 nsew signal input
rlabel metal2 s 308954 352563 309010 353363 6 data_arrays_0_0_ext_ram_rdata2[24]
port 176 nsew signal input
rlabel metal2 s 310058 352563 310114 353363 6 data_arrays_0_0_ext_ram_rdata2[25]
port 177 nsew signal input
rlabel metal2 s 311162 352563 311218 353363 6 data_arrays_0_0_ext_ram_rdata2[26]
port 178 nsew signal input
rlabel metal2 s 312174 352563 312230 353363 6 data_arrays_0_0_ext_ram_rdata2[27]
port 179 nsew signal input
rlabel metal2 s 313278 352563 313334 353363 6 data_arrays_0_0_ext_ram_rdata2[28]
port 180 nsew signal input
rlabel metal2 s 314290 352563 314346 353363 6 data_arrays_0_0_ext_ram_rdata2[29]
port 181 nsew signal input
rlabel metal2 s 285494 352563 285550 353363 6 data_arrays_0_0_ext_ram_rdata2[2]
port 182 nsew signal input
rlabel metal2 s 315394 352563 315450 353363 6 data_arrays_0_0_ext_ram_rdata2[30]
port 183 nsew signal input
rlabel metal2 s 316498 352563 316554 353363 6 data_arrays_0_0_ext_ram_rdata2[31]
port 184 nsew signal input
rlabel metal2 s 317510 352563 317566 353363 6 data_arrays_0_0_ext_ram_rdata2[32]
port 185 nsew signal input
rlabel metal2 s 318614 352563 318670 353363 6 data_arrays_0_0_ext_ram_rdata2[33]
port 186 nsew signal input
rlabel metal2 s 319626 352563 319682 353363 6 data_arrays_0_0_ext_ram_rdata2[34]
port 187 nsew signal input
rlabel metal2 s 320730 352563 320786 353363 6 data_arrays_0_0_ext_ram_rdata2[35]
port 188 nsew signal input
rlabel metal2 s 321834 352563 321890 353363 6 data_arrays_0_0_ext_ram_rdata2[36]
port 189 nsew signal input
rlabel metal2 s 322846 352563 322902 353363 6 data_arrays_0_0_ext_ram_rdata2[37]
port 190 nsew signal input
rlabel metal2 s 323950 352563 324006 353363 6 data_arrays_0_0_ext_ram_rdata2[38]
port 191 nsew signal input
rlabel metal2 s 324962 352563 325018 353363 6 data_arrays_0_0_ext_ram_rdata2[39]
port 192 nsew signal input
rlabel metal2 s 286598 352563 286654 353363 6 data_arrays_0_0_ext_ram_rdata2[3]
port 193 nsew signal input
rlabel metal2 s 326066 352563 326122 353363 6 data_arrays_0_0_ext_ram_rdata2[40]
port 194 nsew signal input
rlabel metal2 s 327170 352563 327226 353363 6 data_arrays_0_0_ext_ram_rdata2[41]
port 195 nsew signal input
rlabel metal2 s 328182 352563 328238 353363 6 data_arrays_0_0_ext_ram_rdata2[42]
port 196 nsew signal input
rlabel metal2 s 329286 352563 329342 353363 6 data_arrays_0_0_ext_ram_rdata2[43]
port 197 nsew signal input
rlabel metal2 s 330298 352563 330354 353363 6 data_arrays_0_0_ext_ram_rdata2[44]
port 198 nsew signal input
rlabel metal2 s 331402 352563 331458 353363 6 data_arrays_0_0_ext_ram_rdata2[45]
port 199 nsew signal input
rlabel metal2 s 332506 352563 332562 353363 6 data_arrays_0_0_ext_ram_rdata2[46]
port 200 nsew signal input
rlabel metal2 s 333518 352563 333574 353363 6 data_arrays_0_0_ext_ram_rdata2[47]
port 201 nsew signal input
rlabel metal2 s 334622 352563 334678 353363 6 data_arrays_0_0_ext_ram_rdata2[48]
port 202 nsew signal input
rlabel metal2 s 335634 352563 335690 353363 6 data_arrays_0_0_ext_ram_rdata2[49]
port 203 nsew signal input
rlabel metal2 s 287610 352563 287666 353363 6 data_arrays_0_0_ext_ram_rdata2[4]
port 204 nsew signal input
rlabel metal2 s 336738 352563 336794 353363 6 data_arrays_0_0_ext_ram_rdata2[50]
port 205 nsew signal input
rlabel metal2 s 337842 352563 337898 353363 6 data_arrays_0_0_ext_ram_rdata2[51]
port 206 nsew signal input
rlabel metal2 s 338854 352563 338910 353363 6 data_arrays_0_0_ext_ram_rdata2[52]
port 207 nsew signal input
rlabel metal2 s 339958 352563 340014 353363 6 data_arrays_0_0_ext_ram_rdata2[53]
port 208 nsew signal input
rlabel metal2 s 340970 352563 341026 353363 6 data_arrays_0_0_ext_ram_rdata2[54]
port 209 nsew signal input
rlabel metal2 s 342074 352563 342130 353363 6 data_arrays_0_0_ext_ram_rdata2[55]
port 210 nsew signal input
rlabel metal2 s 343178 352563 343234 353363 6 data_arrays_0_0_ext_ram_rdata2[56]
port 211 nsew signal input
rlabel metal2 s 344190 352563 344246 353363 6 data_arrays_0_0_ext_ram_rdata2[57]
port 212 nsew signal input
rlabel metal2 s 345294 352563 345350 353363 6 data_arrays_0_0_ext_ram_rdata2[58]
port 213 nsew signal input
rlabel metal2 s 346306 352563 346362 353363 6 data_arrays_0_0_ext_ram_rdata2[59]
port 214 nsew signal input
rlabel metal2 s 288714 352563 288770 353363 6 data_arrays_0_0_ext_ram_rdata2[5]
port 215 nsew signal input
rlabel metal2 s 347410 352563 347466 353363 6 data_arrays_0_0_ext_ram_rdata2[60]
port 216 nsew signal input
rlabel metal2 s 348514 352563 348570 353363 6 data_arrays_0_0_ext_ram_rdata2[61]
port 217 nsew signal input
rlabel metal2 s 349526 352563 349582 353363 6 data_arrays_0_0_ext_ram_rdata2[62]
port 218 nsew signal input
rlabel metal2 s 350630 352563 350686 353363 6 data_arrays_0_0_ext_ram_rdata2[63]
port 219 nsew signal input
rlabel metal2 s 289726 352563 289782 353363 6 data_arrays_0_0_ext_ram_rdata2[6]
port 220 nsew signal input
rlabel metal2 s 290830 352563 290886 353363 6 data_arrays_0_0_ext_ram_rdata2[7]
port 221 nsew signal input
rlabel metal2 s 291934 352563 291990 353363 6 data_arrays_0_0_ext_ram_rdata2[8]
port 222 nsew signal input
rlabel metal2 s 292946 352563 293002 353363 6 data_arrays_0_0_ext_ram_rdata2[9]
port 223 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 data_arrays_0_0_ext_ram_wdata[0]
port 224 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 data_arrays_0_0_ext_ram_wdata[10]
port 225 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 data_arrays_0_0_ext_ram_wdata[11]
port 226 nsew signal output
rlabel metal3 s 0 135056 800 135176 6 data_arrays_0_0_ext_ram_wdata[12]
port 227 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 data_arrays_0_0_ext_ram_wdata[13]
port 228 nsew signal output
rlabel metal3 s 0 138184 800 138304 6 data_arrays_0_0_ext_ram_wdata[14]
port 229 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 data_arrays_0_0_ext_ram_wdata[15]
port 230 nsew signal output
rlabel metal3 s 0 141312 800 141432 6 data_arrays_0_0_ext_ram_wdata[16]
port 231 nsew signal output
rlabel metal3 s 0 142944 800 143064 6 data_arrays_0_0_ext_ram_wdata[17]
port 232 nsew signal output
rlabel metal3 s 0 144440 800 144560 6 data_arrays_0_0_ext_ram_wdata[18]
port 233 nsew signal output
rlabel metal3 s 0 146072 800 146192 6 data_arrays_0_0_ext_ram_wdata[19]
port 234 nsew signal output
rlabel metal3 s 0 117920 800 118040 6 data_arrays_0_0_ext_ram_wdata[1]
port 235 nsew signal output
rlabel metal3 s 0 147568 800 147688 6 data_arrays_0_0_ext_ram_wdata[20]
port 236 nsew signal output
rlabel metal3 s 0 149200 800 149320 6 data_arrays_0_0_ext_ram_wdata[21]
port 237 nsew signal output
rlabel metal3 s 0 150696 800 150816 6 data_arrays_0_0_ext_ram_wdata[22]
port 238 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 data_arrays_0_0_ext_ram_wdata[23]
port 239 nsew signal output
rlabel metal3 s 0 153824 800 153944 6 data_arrays_0_0_ext_ram_wdata[24]
port 240 nsew signal output
rlabel metal3 s 0 155456 800 155576 6 data_arrays_0_0_ext_ram_wdata[25]
port 241 nsew signal output
rlabel metal3 s 0 156952 800 157072 6 data_arrays_0_0_ext_ram_wdata[26]
port 242 nsew signal output
rlabel metal3 s 0 158584 800 158704 6 data_arrays_0_0_ext_ram_wdata[27]
port 243 nsew signal output
rlabel metal3 s 0 160080 800 160200 6 data_arrays_0_0_ext_ram_wdata[28]
port 244 nsew signal output
rlabel metal3 s 0 161712 800 161832 6 data_arrays_0_0_ext_ram_wdata[29]
port 245 nsew signal output
rlabel metal3 s 0 119416 800 119536 6 data_arrays_0_0_ext_ram_wdata[2]
port 246 nsew signal output
rlabel metal3 s 0 163208 800 163328 6 data_arrays_0_0_ext_ram_wdata[30]
port 247 nsew signal output
rlabel metal3 s 0 164840 800 164960 6 data_arrays_0_0_ext_ram_wdata[31]
port 248 nsew signal output
rlabel metal3 s 0 166336 800 166456 6 data_arrays_0_0_ext_ram_wdata[32]
port 249 nsew signal output
rlabel metal3 s 0 167968 800 168088 6 data_arrays_0_0_ext_ram_wdata[33]
port 250 nsew signal output
rlabel metal3 s 0 169464 800 169584 6 data_arrays_0_0_ext_ram_wdata[34]
port 251 nsew signal output
rlabel metal3 s 0 171096 800 171216 6 data_arrays_0_0_ext_ram_wdata[35]
port 252 nsew signal output
rlabel metal3 s 0 172592 800 172712 6 data_arrays_0_0_ext_ram_wdata[36]
port 253 nsew signal output
rlabel metal3 s 0 174224 800 174344 6 data_arrays_0_0_ext_ram_wdata[37]
port 254 nsew signal output
rlabel metal3 s 0 175720 800 175840 6 data_arrays_0_0_ext_ram_wdata[38]
port 255 nsew signal output
rlabel metal3 s 0 177352 800 177472 6 data_arrays_0_0_ext_ram_wdata[39]
port 256 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 data_arrays_0_0_ext_ram_wdata[3]
port 257 nsew signal output
rlabel metal3 s 0 178848 800 178968 6 data_arrays_0_0_ext_ram_wdata[40]
port 258 nsew signal output
rlabel metal3 s 0 180344 800 180464 6 data_arrays_0_0_ext_ram_wdata[41]
port 259 nsew signal output
rlabel metal3 s 0 181976 800 182096 6 data_arrays_0_0_ext_ram_wdata[42]
port 260 nsew signal output
rlabel metal3 s 0 183472 800 183592 6 data_arrays_0_0_ext_ram_wdata[43]
port 261 nsew signal output
rlabel metal3 s 0 185104 800 185224 6 data_arrays_0_0_ext_ram_wdata[44]
port 262 nsew signal output
rlabel metal3 s 0 186600 800 186720 6 data_arrays_0_0_ext_ram_wdata[45]
port 263 nsew signal output
rlabel metal3 s 0 188232 800 188352 6 data_arrays_0_0_ext_ram_wdata[46]
port 264 nsew signal output
rlabel metal3 s 0 189728 800 189848 6 data_arrays_0_0_ext_ram_wdata[47]
port 265 nsew signal output
rlabel metal3 s 0 191360 800 191480 6 data_arrays_0_0_ext_ram_wdata[48]
port 266 nsew signal output
rlabel metal3 s 0 192856 800 192976 6 data_arrays_0_0_ext_ram_wdata[49]
port 267 nsew signal output
rlabel metal3 s 0 122544 800 122664 6 data_arrays_0_0_ext_ram_wdata[4]
port 268 nsew signal output
rlabel metal3 s 0 194488 800 194608 6 data_arrays_0_0_ext_ram_wdata[50]
port 269 nsew signal output
rlabel metal3 s 0 195984 800 196104 6 data_arrays_0_0_ext_ram_wdata[51]
port 270 nsew signal output
rlabel metal3 s 0 197616 800 197736 6 data_arrays_0_0_ext_ram_wdata[52]
port 271 nsew signal output
rlabel metal3 s 0 199112 800 199232 6 data_arrays_0_0_ext_ram_wdata[53]
port 272 nsew signal output
rlabel metal3 s 0 200744 800 200864 6 data_arrays_0_0_ext_ram_wdata[54]
port 273 nsew signal output
rlabel metal3 s 0 202240 800 202360 6 data_arrays_0_0_ext_ram_wdata[55]
port 274 nsew signal output
rlabel metal3 s 0 203872 800 203992 6 data_arrays_0_0_ext_ram_wdata[56]
port 275 nsew signal output
rlabel metal3 s 0 205368 800 205488 6 data_arrays_0_0_ext_ram_wdata[57]
port 276 nsew signal output
rlabel metal3 s 0 207000 800 207120 6 data_arrays_0_0_ext_ram_wdata[58]
port 277 nsew signal output
rlabel metal3 s 0 208496 800 208616 6 data_arrays_0_0_ext_ram_wdata[59]
port 278 nsew signal output
rlabel metal3 s 0 124176 800 124296 6 data_arrays_0_0_ext_ram_wdata[5]
port 279 nsew signal output
rlabel metal3 s 0 210128 800 210248 6 data_arrays_0_0_ext_ram_wdata[60]
port 280 nsew signal output
rlabel metal3 s 0 211624 800 211744 6 data_arrays_0_0_ext_ram_wdata[61]
port 281 nsew signal output
rlabel metal3 s 0 213256 800 213376 6 data_arrays_0_0_ext_ram_wdata[62]
port 282 nsew signal output
rlabel metal3 s 0 214752 800 214872 6 data_arrays_0_0_ext_ram_wdata[63]
port 283 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 data_arrays_0_0_ext_ram_wdata[6]
port 284 nsew signal output
rlabel metal3 s 0 127304 800 127424 6 data_arrays_0_0_ext_ram_wdata[7]
port 285 nsew signal output
rlabel metal3 s 0 128800 800 128920 6 data_arrays_0_0_ext_ram_wdata[8]
port 286 nsew signal output
rlabel metal3 s 0 130432 800 130552 6 data_arrays_0_0_ext_ram_wdata[9]
port 287 nsew signal output
rlabel metal3 s 0 225768 800 225888 6 data_arrays_0_0_ext_ram_web
port 288 nsew signal output
rlabel metal3 s 0 216384 800 216504 6 data_arrays_0_0_ext_ram_wmask[0]
port 289 nsew signal output
rlabel metal3 s 0 217880 800 218000 6 data_arrays_0_0_ext_ram_wmask[1]
port 290 nsew signal output
rlabel metal2 s 161662 352563 161718 353363 6 io_in[0]
port 291 nsew signal input
rlabel metal2 s 193678 352563 193734 353363 6 io_in[10]
port 292 nsew signal input
rlabel metal2 s 196898 352563 196954 353363 6 io_in[11]
port 293 nsew signal input
rlabel metal2 s 200118 352563 200174 353363 6 io_in[12]
port 294 nsew signal input
rlabel metal2 s 203246 352563 203302 353363 6 io_in[13]
port 295 nsew signal input
rlabel metal2 s 206466 352563 206522 353363 6 io_in[14]
port 296 nsew signal input
rlabel metal2 s 209686 352563 209742 353363 6 io_in[15]
port 297 nsew signal input
rlabel metal2 s 212906 352563 212962 353363 6 io_in[16]
port 298 nsew signal input
rlabel metal2 s 216126 352563 216182 353363 6 io_in[17]
port 299 nsew signal input
rlabel metal2 s 219254 352563 219310 353363 6 io_in[18]
port 300 nsew signal input
rlabel metal2 s 222474 352563 222530 353363 6 io_in[19]
port 301 nsew signal input
rlabel metal2 s 164882 352563 164938 353363 6 io_in[1]
port 302 nsew signal input
rlabel metal2 s 225694 352563 225750 353363 6 io_in[20]
port 303 nsew signal input
rlabel metal2 s 228914 352563 228970 353363 6 io_in[21]
port 304 nsew signal input
rlabel metal2 s 232134 352563 232190 353363 6 io_in[22]
port 305 nsew signal input
rlabel metal2 s 235354 352563 235410 353363 6 io_in[23]
port 306 nsew signal input
rlabel metal2 s 238482 352563 238538 353363 6 io_in[24]
port 307 nsew signal input
rlabel metal2 s 241702 352563 241758 353363 6 io_in[25]
port 308 nsew signal input
rlabel metal2 s 244922 352563 244978 353363 6 io_in[26]
port 309 nsew signal input
rlabel metal2 s 248142 352563 248198 353363 6 io_in[27]
port 310 nsew signal input
rlabel metal2 s 251362 352563 251418 353363 6 io_in[28]
port 311 nsew signal input
rlabel metal2 s 254490 352563 254546 353363 6 io_in[29]
port 312 nsew signal input
rlabel metal2 s 168010 352563 168066 353363 6 io_in[2]
port 313 nsew signal input
rlabel metal2 s 257710 352563 257766 353363 6 io_in[30]
port 314 nsew signal input
rlabel metal2 s 260930 352563 260986 353363 6 io_in[31]
port 315 nsew signal input
rlabel metal2 s 264150 352563 264206 353363 6 io_in[32]
port 316 nsew signal input
rlabel metal2 s 267370 352563 267426 353363 6 io_in[33]
port 317 nsew signal input
rlabel metal2 s 270590 352563 270646 353363 6 io_in[34]
port 318 nsew signal input
rlabel metal2 s 273718 352563 273774 353363 6 io_in[35]
port 319 nsew signal input
rlabel metal2 s 276938 352563 276994 353363 6 io_in[36]
port 320 nsew signal input
rlabel metal2 s 280158 352563 280214 353363 6 io_in[37]
port 321 nsew signal input
rlabel metal2 s 171230 352563 171286 353363 6 io_in[3]
port 322 nsew signal input
rlabel metal2 s 174450 352563 174506 353363 6 io_in[4]
port 323 nsew signal input
rlabel metal2 s 177670 352563 177726 353363 6 io_in[5]
port 324 nsew signal input
rlabel metal2 s 180890 352563 180946 353363 6 io_in[6]
port 325 nsew signal input
rlabel metal2 s 184110 352563 184166 353363 6 io_in[7]
port 326 nsew signal input
rlabel metal2 s 187238 352563 187294 353363 6 io_in[8]
port 327 nsew signal input
rlabel metal2 s 190458 352563 190514 353363 6 io_in[9]
port 328 nsew signal input
rlabel metal2 s 162674 352563 162730 353363 6 io_oeb[0]
port 329 nsew signal output
rlabel metal2 s 194782 352563 194838 353363 6 io_oeb[10]
port 330 nsew signal output
rlabel metal2 s 197910 352563 197966 353363 6 io_oeb[11]
port 331 nsew signal output
rlabel metal2 s 201130 352563 201186 353363 6 io_oeb[12]
port 332 nsew signal output
rlabel metal2 s 204350 352563 204406 353363 6 io_oeb[13]
port 333 nsew signal output
rlabel metal2 s 207570 352563 207626 353363 6 io_oeb[14]
port 334 nsew signal output
rlabel metal2 s 210790 352563 210846 353363 6 io_oeb[15]
port 335 nsew signal output
rlabel metal2 s 213918 352563 213974 353363 6 io_oeb[16]
port 336 nsew signal output
rlabel metal2 s 217138 352563 217194 353363 6 io_oeb[17]
port 337 nsew signal output
rlabel metal2 s 220358 352563 220414 353363 6 io_oeb[18]
port 338 nsew signal output
rlabel metal2 s 223578 352563 223634 353363 6 io_oeb[19]
port 339 nsew signal output
rlabel metal2 s 165894 352563 165950 353363 6 io_oeb[1]
port 340 nsew signal output
rlabel metal2 s 226798 352563 226854 353363 6 io_oeb[20]
port 341 nsew signal output
rlabel metal2 s 230018 352563 230074 353363 6 io_oeb[21]
port 342 nsew signal output
rlabel metal2 s 233146 352563 233202 353363 6 io_oeb[22]
port 343 nsew signal output
rlabel metal2 s 236366 352563 236422 353363 6 io_oeb[23]
port 344 nsew signal output
rlabel metal2 s 239586 352563 239642 353363 6 io_oeb[24]
port 345 nsew signal output
rlabel metal2 s 242806 352563 242862 353363 6 io_oeb[25]
port 346 nsew signal output
rlabel metal2 s 246026 352563 246082 353363 6 io_oeb[26]
port 347 nsew signal output
rlabel metal2 s 249154 352563 249210 353363 6 io_oeb[27]
port 348 nsew signal output
rlabel metal2 s 252374 352563 252430 353363 6 io_oeb[28]
port 349 nsew signal output
rlabel metal2 s 255594 352563 255650 353363 6 io_oeb[29]
port 350 nsew signal output
rlabel metal2 s 169114 352563 169170 353363 6 io_oeb[2]
port 351 nsew signal output
rlabel metal2 s 258814 352563 258870 353363 6 io_oeb[30]
port 352 nsew signal output
rlabel metal2 s 262034 352563 262090 353363 6 io_oeb[31]
port 353 nsew signal output
rlabel metal2 s 265254 352563 265310 353363 6 io_oeb[32]
port 354 nsew signal output
rlabel metal2 s 268382 352563 268438 353363 6 io_oeb[33]
port 355 nsew signal output
rlabel metal2 s 271602 352563 271658 353363 6 io_oeb[34]
port 356 nsew signal output
rlabel metal2 s 274822 352563 274878 353363 6 io_oeb[35]
port 357 nsew signal output
rlabel metal2 s 278042 352563 278098 353363 6 io_oeb[36]
port 358 nsew signal output
rlabel metal2 s 281262 352563 281318 353363 6 io_oeb[37]
port 359 nsew signal output
rlabel metal2 s 172334 352563 172390 353363 6 io_oeb[3]
port 360 nsew signal output
rlabel metal2 s 175554 352563 175610 353363 6 io_oeb[4]
port 361 nsew signal output
rlabel metal2 s 178774 352563 178830 353363 6 io_oeb[5]
port 362 nsew signal output
rlabel metal2 s 181902 352563 181958 353363 6 io_oeb[6]
port 363 nsew signal output
rlabel metal2 s 185122 352563 185178 353363 6 io_oeb[7]
port 364 nsew signal output
rlabel metal2 s 188342 352563 188398 353363 6 io_oeb[8]
port 365 nsew signal output
rlabel metal2 s 191562 352563 191618 353363 6 io_oeb[9]
port 366 nsew signal output
rlabel metal2 s 163778 352563 163834 353363 6 io_out[0]
port 367 nsew signal output
rlabel metal2 s 195794 352563 195850 353363 6 io_out[10]
port 368 nsew signal output
rlabel metal2 s 199014 352563 199070 353363 6 io_out[11]
port 369 nsew signal output
rlabel metal2 s 202234 352563 202290 353363 6 io_out[12]
port 370 nsew signal output
rlabel metal2 s 205454 352563 205510 353363 6 io_out[13]
port 371 nsew signal output
rlabel metal2 s 208582 352563 208638 353363 6 io_out[14]
port 372 nsew signal output
rlabel metal2 s 211802 352563 211858 353363 6 io_out[15]
port 373 nsew signal output
rlabel metal2 s 215022 352563 215078 353363 6 io_out[16]
port 374 nsew signal output
rlabel metal2 s 218242 352563 218298 353363 6 io_out[17]
port 375 nsew signal output
rlabel metal2 s 221462 352563 221518 353363 6 io_out[18]
port 376 nsew signal output
rlabel metal2 s 224682 352563 224738 353363 6 io_out[19]
port 377 nsew signal output
rlabel metal2 s 166998 352563 167054 353363 6 io_out[1]
port 378 nsew signal output
rlabel metal2 s 227810 352563 227866 353363 6 io_out[20]
port 379 nsew signal output
rlabel metal2 s 231030 352563 231086 353363 6 io_out[21]
port 380 nsew signal output
rlabel metal2 s 234250 352563 234306 353363 6 io_out[22]
port 381 nsew signal output
rlabel metal2 s 237470 352563 237526 353363 6 io_out[23]
port 382 nsew signal output
rlabel metal2 s 240690 352563 240746 353363 6 io_out[24]
port 383 nsew signal output
rlabel metal2 s 243818 352563 243874 353363 6 io_out[25]
port 384 nsew signal output
rlabel metal2 s 247038 352563 247094 353363 6 io_out[26]
port 385 nsew signal output
rlabel metal2 s 250258 352563 250314 353363 6 io_out[27]
port 386 nsew signal output
rlabel metal2 s 253478 352563 253534 353363 6 io_out[28]
port 387 nsew signal output
rlabel metal2 s 256698 352563 256754 353363 6 io_out[29]
port 388 nsew signal output
rlabel metal2 s 170218 352563 170274 353363 6 io_out[2]
port 389 nsew signal output
rlabel metal2 s 259826 352563 259882 353363 6 io_out[30]
port 390 nsew signal output
rlabel metal2 s 263046 352563 263102 353363 6 io_out[31]
port 391 nsew signal output
rlabel metal2 s 266266 352563 266322 353363 6 io_out[32]
port 392 nsew signal output
rlabel metal2 s 269486 352563 269542 353363 6 io_out[33]
port 393 nsew signal output
rlabel metal2 s 272706 352563 272762 353363 6 io_out[34]
port 394 nsew signal output
rlabel metal2 s 275926 352563 275982 353363 6 io_out[35]
port 395 nsew signal output
rlabel metal2 s 279054 352563 279110 353363 6 io_out[36]
port 396 nsew signal output
rlabel metal2 s 282274 352563 282330 353363 6 io_out[37]
port 397 nsew signal output
rlabel metal2 s 173346 352563 173402 353363 6 io_out[3]
port 398 nsew signal output
rlabel metal2 s 176566 352563 176622 353363 6 io_out[4]
port 399 nsew signal output
rlabel metal2 s 179786 352563 179842 353363 6 io_out[5]
port 400 nsew signal output
rlabel metal2 s 183006 352563 183062 353363 6 io_out[6]
port 401 nsew signal output
rlabel metal2 s 186226 352563 186282 353363 6 io_out[7]
port 402 nsew signal output
rlabel metal2 s 189446 352563 189502 353363 6 io_out[8]
port 403 nsew signal output
rlabel metal2 s 192574 352563 192630 353363 6 io_out[9]
port 404 nsew signal output
rlabel metal2 s 349342 0 349398 800 6 irq[0]
port 405 nsew signal output
rlabel metal2 s 350078 0 350134 800 6 irq[1]
port 406 nsew signal output
rlabel metal2 s 350814 0 350870 800 6 irq[2]
port 407 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_in[0]
port 408 nsew signal input
rlabel metal2 s 289542 0 289598 800 6 la_data_in[100]
port 409 nsew signal input
rlabel metal2 s 291658 0 291714 800 6 la_data_in[101]
port 410 nsew signal input
rlabel metal2 s 293774 0 293830 800 6 la_data_in[102]
port 411 nsew signal input
rlabel metal2 s 295890 0 295946 800 6 la_data_in[103]
port 412 nsew signal input
rlabel metal2 s 298098 0 298154 800 6 la_data_in[104]
port 413 nsew signal input
rlabel metal2 s 300214 0 300270 800 6 la_data_in[105]
port 414 nsew signal input
rlabel metal2 s 302330 0 302386 800 6 la_data_in[106]
port 415 nsew signal input
rlabel metal2 s 304446 0 304502 800 6 la_data_in[107]
port 416 nsew signal input
rlabel metal2 s 306654 0 306710 800 6 la_data_in[108]
port 417 nsew signal input
rlabel metal2 s 308770 0 308826 800 6 la_data_in[109]
port 418 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_data_in[10]
port 419 nsew signal input
rlabel metal2 s 310886 0 310942 800 6 la_data_in[110]
port 420 nsew signal input
rlabel metal2 s 313002 0 313058 800 6 la_data_in[111]
port 421 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_data_in[112]
port 422 nsew signal input
rlabel metal2 s 317326 0 317382 800 6 la_data_in[113]
port 423 nsew signal input
rlabel metal2 s 319442 0 319498 800 6 la_data_in[114]
port 424 nsew signal input
rlabel metal2 s 321558 0 321614 800 6 la_data_in[115]
port 425 nsew signal input
rlabel metal2 s 323674 0 323730 800 6 la_data_in[116]
port 426 nsew signal input
rlabel metal2 s 325882 0 325938 800 6 la_data_in[117]
port 427 nsew signal input
rlabel metal2 s 327998 0 328054 800 6 la_data_in[118]
port 428 nsew signal input
rlabel metal2 s 330114 0 330170 800 6 la_data_in[119]
port 429 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[11]
port 430 nsew signal input
rlabel metal2 s 332230 0 332286 800 6 la_data_in[120]
port 431 nsew signal input
rlabel metal2 s 334438 0 334494 800 6 la_data_in[121]
port 432 nsew signal input
rlabel metal2 s 336554 0 336610 800 6 la_data_in[122]
port 433 nsew signal input
rlabel metal2 s 338670 0 338726 800 6 la_data_in[123]
port 434 nsew signal input
rlabel metal2 s 340786 0 340842 800 6 la_data_in[124]
port 435 nsew signal input
rlabel metal2 s 342994 0 343050 800 6 la_data_in[125]
port 436 nsew signal input
rlabel metal2 s 345110 0 345166 800 6 la_data_in[126]
port 437 nsew signal input
rlabel metal2 s 347226 0 347282 800 6 la_data_in[127]
port 438 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[12]
port 439 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_data_in[13]
port 440 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_data_in[14]
port 441 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[15]
port 442 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[16]
port 443 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_data_in[17]
port 444 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[18]
port 445 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[19]
port 446 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[1]
port 447 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[20]
port 448 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_data_in[21]
port 449 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[22]
port 450 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[23]
port 451 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_data_in[24]
port 452 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_data_in[25]
port 453 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[26]
port 454 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[27]
port 455 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_data_in[28]
port 456 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[29]
port 457 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[2]
port 458 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_data_in[30]
port 459 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_data_in[31]
port 460 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[32]
port 461 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[33]
port 462 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[34]
port 463 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_data_in[35]
port 464 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[36]
port 465 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_data_in[37]
port 466 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[38]
port 467 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_data_in[39]
port 468 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[3]
port 469 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_data_in[40]
port 470 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[41]
port 471 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_data_in[42]
port 472 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[43]
port 473 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_data_in[44]
port 474 nsew signal input
rlabel metal2 s 171966 0 172022 800 6 la_data_in[45]
port 475 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_data_in[46]
port 476 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_data_in[47]
port 477 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_data_in[48]
port 478 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_data_in[49]
port 479 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[4]
port 480 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_data_in[50]
port 481 nsew signal input
rlabel metal2 s 184754 0 184810 800 6 la_data_in[51]
port 482 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_data_in[52]
port 483 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_data_in[53]
port 484 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_data_in[54]
port 485 nsew signal input
rlabel metal2 s 193310 0 193366 800 6 la_data_in[55]
port 486 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_data_in[56]
port 487 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_data_in[57]
port 488 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 la_data_in[58]
port 489 nsew signal input
rlabel metal2 s 201866 0 201922 800 6 la_data_in[59]
port 490 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_data_in[5]
port 491 nsew signal input
rlabel metal2 s 203982 0 204038 800 6 la_data_in[60]
port 492 nsew signal input
rlabel metal2 s 206190 0 206246 800 6 la_data_in[61]
port 493 nsew signal input
rlabel metal2 s 208306 0 208362 800 6 la_data_in[62]
port 494 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_data_in[63]
port 495 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_data_in[64]
port 496 nsew signal input
rlabel metal2 s 214746 0 214802 800 6 la_data_in[65]
port 497 nsew signal input
rlabel metal2 s 216862 0 216918 800 6 la_data_in[66]
port 498 nsew signal input
rlabel metal2 s 218978 0 219034 800 6 la_data_in[67]
port 499 nsew signal input
rlabel metal2 s 221094 0 221150 800 6 la_data_in[68]
port 500 nsew signal input
rlabel metal2 s 223302 0 223358 800 6 la_data_in[69]
port 501 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[6]
port 502 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_data_in[70]
port 503 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 la_data_in[71]
port 504 nsew signal input
rlabel metal2 s 229650 0 229706 800 6 la_data_in[72]
port 505 nsew signal input
rlabel metal2 s 231766 0 231822 800 6 la_data_in[73]
port 506 nsew signal input
rlabel metal2 s 233974 0 234030 800 6 la_data_in[74]
port 507 nsew signal input
rlabel metal2 s 236090 0 236146 800 6 la_data_in[75]
port 508 nsew signal input
rlabel metal2 s 238206 0 238262 800 6 la_data_in[76]
port 509 nsew signal input
rlabel metal2 s 240322 0 240378 800 6 la_data_in[77]
port 510 nsew signal input
rlabel metal2 s 242530 0 242586 800 6 la_data_in[78]
port 511 nsew signal input
rlabel metal2 s 244646 0 244702 800 6 la_data_in[79]
port 512 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[7]
port 513 nsew signal input
rlabel metal2 s 246762 0 246818 800 6 la_data_in[80]
port 514 nsew signal input
rlabel metal2 s 248878 0 248934 800 6 la_data_in[81]
port 515 nsew signal input
rlabel metal2 s 251086 0 251142 800 6 la_data_in[82]
port 516 nsew signal input
rlabel metal2 s 253202 0 253258 800 6 la_data_in[83]
port 517 nsew signal input
rlabel metal2 s 255318 0 255374 800 6 la_data_in[84]
port 518 nsew signal input
rlabel metal2 s 257434 0 257490 800 6 la_data_in[85]
port 519 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_data_in[86]
port 520 nsew signal input
rlabel metal2 s 261758 0 261814 800 6 la_data_in[87]
port 521 nsew signal input
rlabel metal2 s 263874 0 263930 800 6 la_data_in[88]
port 522 nsew signal input
rlabel metal2 s 265990 0 266046 800 6 la_data_in[89]
port 523 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[8]
port 524 nsew signal input
rlabel metal2 s 268106 0 268162 800 6 la_data_in[90]
port 525 nsew signal input
rlabel metal2 s 270314 0 270370 800 6 la_data_in[91]
port 526 nsew signal input
rlabel metal2 s 272430 0 272486 800 6 la_data_in[92]
port 527 nsew signal input
rlabel metal2 s 274546 0 274602 800 6 la_data_in[93]
port 528 nsew signal input
rlabel metal2 s 276662 0 276718 800 6 la_data_in[94]
port 529 nsew signal input
rlabel metal2 s 278870 0 278926 800 6 la_data_in[95]
port 530 nsew signal input
rlabel metal2 s 280986 0 281042 800 6 la_data_in[96]
port 531 nsew signal input
rlabel metal2 s 283102 0 283158 800 6 la_data_in[97]
port 532 nsew signal input
rlabel metal2 s 285218 0 285274 800 6 la_data_in[98]
port 533 nsew signal input
rlabel metal2 s 287426 0 287482 800 6 la_data_in[99]
port 534 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_data_in[9]
port 535 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_out[0]
port 536 nsew signal output
rlabel metal2 s 290186 0 290242 800 6 la_data_out[100]
port 537 nsew signal output
rlabel metal2 s 292394 0 292450 800 6 la_data_out[101]
port 538 nsew signal output
rlabel metal2 s 294510 0 294566 800 6 la_data_out[102]
port 539 nsew signal output
rlabel metal2 s 296626 0 296682 800 6 la_data_out[103]
port 540 nsew signal output
rlabel metal2 s 298742 0 298798 800 6 la_data_out[104]
port 541 nsew signal output
rlabel metal2 s 300950 0 301006 800 6 la_data_out[105]
port 542 nsew signal output
rlabel metal2 s 303066 0 303122 800 6 la_data_out[106]
port 543 nsew signal output
rlabel metal2 s 305182 0 305238 800 6 la_data_out[107]
port 544 nsew signal output
rlabel metal2 s 307298 0 307354 800 6 la_data_out[108]
port 545 nsew signal output
rlabel metal2 s 309506 0 309562 800 6 la_data_out[109]
port 546 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[10]
port 547 nsew signal output
rlabel metal2 s 311622 0 311678 800 6 la_data_out[110]
port 548 nsew signal output
rlabel metal2 s 313738 0 313794 800 6 la_data_out[111]
port 549 nsew signal output
rlabel metal2 s 315854 0 315910 800 6 la_data_out[112]
port 550 nsew signal output
rlabel metal2 s 318062 0 318118 800 6 la_data_out[113]
port 551 nsew signal output
rlabel metal2 s 320178 0 320234 800 6 la_data_out[114]
port 552 nsew signal output
rlabel metal2 s 322294 0 322350 800 6 la_data_out[115]
port 553 nsew signal output
rlabel metal2 s 324410 0 324466 800 6 la_data_out[116]
port 554 nsew signal output
rlabel metal2 s 326526 0 326582 800 6 la_data_out[117]
port 555 nsew signal output
rlabel metal2 s 328734 0 328790 800 6 la_data_out[118]
port 556 nsew signal output
rlabel metal2 s 330850 0 330906 800 6 la_data_out[119]
port 557 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[11]
port 558 nsew signal output
rlabel metal2 s 332966 0 333022 800 6 la_data_out[120]
port 559 nsew signal output
rlabel metal2 s 335082 0 335138 800 6 la_data_out[121]
port 560 nsew signal output
rlabel metal2 s 337290 0 337346 800 6 la_data_out[122]
port 561 nsew signal output
rlabel metal2 s 339406 0 339462 800 6 la_data_out[123]
port 562 nsew signal output
rlabel metal2 s 341522 0 341578 800 6 la_data_out[124]
port 563 nsew signal output
rlabel metal2 s 343638 0 343694 800 6 la_data_out[125]
port 564 nsew signal output
rlabel metal2 s 345846 0 345902 800 6 la_data_out[126]
port 565 nsew signal output
rlabel metal2 s 347962 0 348018 800 6 la_data_out[127]
port 566 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[12]
port 567 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[13]
port 568 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[14]
port 569 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[15]
port 570 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[16]
port 571 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[17]
port 572 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 la_data_out[18]
port 573 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 la_data_out[19]
port 574 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[1]
port 575 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 la_data_out[20]
port 576 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[21]
port 577 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 la_data_out[22]
port 578 nsew signal output
rlabel metal2 s 125690 0 125746 800 6 la_data_out[23]
port 579 nsew signal output
rlabel metal2 s 127806 0 127862 800 6 la_data_out[24]
port 580 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 la_data_out[25]
port 581 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[26]
port 582 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[27]
port 583 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[28]
port 584 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 la_data_out[29]
port 585 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[2]
port 586 nsew signal output
rlabel metal2 s 140594 0 140650 800 6 la_data_out[30]
port 587 nsew signal output
rlabel metal2 s 142710 0 142766 800 6 la_data_out[31]
port 588 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[32]
port 589 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[33]
port 590 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[34]
port 591 nsew signal output
rlabel metal2 s 151266 0 151322 800 6 la_data_out[35]
port 592 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 la_data_out[36]
port 593 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[37]
port 594 nsew signal output
rlabel metal2 s 157706 0 157762 800 6 la_data_out[38]
port 595 nsew signal output
rlabel metal2 s 159822 0 159878 800 6 la_data_out[39]
port 596 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[3]
port 597 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[40]
port 598 nsew signal output
rlabel metal2 s 164146 0 164202 800 6 la_data_out[41]
port 599 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 la_data_out[42]
port 600 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 la_data_out[43]
port 601 nsew signal output
rlabel metal2 s 170494 0 170550 800 6 la_data_out[44]
port 602 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 la_data_out[45]
port 603 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[46]
port 604 nsew signal output
rlabel metal2 s 176934 0 176990 800 6 la_data_out[47]
port 605 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 la_data_out[48]
port 606 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 la_data_out[49]
port 607 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[4]
port 608 nsew signal output
rlabel metal2 s 183374 0 183430 800 6 la_data_out[50]
port 609 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 la_data_out[51]
port 610 nsew signal output
rlabel metal2 s 187606 0 187662 800 6 la_data_out[52]
port 611 nsew signal output
rlabel metal2 s 189814 0 189870 800 6 la_data_out[53]
port 612 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 la_data_out[54]
port 613 nsew signal output
rlabel metal2 s 194046 0 194102 800 6 la_data_out[55]
port 614 nsew signal output
rlabel metal2 s 196162 0 196218 800 6 la_data_out[56]
port 615 nsew signal output
rlabel metal2 s 198278 0 198334 800 6 la_data_out[57]
port 616 nsew signal output
rlabel metal2 s 200486 0 200542 800 6 la_data_out[58]
port 617 nsew signal output
rlabel metal2 s 202602 0 202658 800 6 la_data_out[59]
port 618 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[5]
port 619 nsew signal output
rlabel metal2 s 204718 0 204774 800 6 la_data_out[60]
port 620 nsew signal output
rlabel metal2 s 206834 0 206890 800 6 la_data_out[61]
port 621 nsew signal output
rlabel metal2 s 209042 0 209098 800 6 la_data_out[62]
port 622 nsew signal output
rlabel metal2 s 211158 0 211214 800 6 la_data_out[63]
port 623 nsew signal output
rlabel metal2 s 213274 0 213330 800 6 la_data_out[64]
port 624 nsew signal output
rlabel metal2 s 215390 0 215446 800 6 la_data_out[65]
port 625 nsew signal output
rlabel metal2 s 217598 0 217654 800 6 la_data_out[66]
port 626 nsew signal output
rlabel metal2 s 219714 0 219770 800 6 la_data_out[67]
port 627 nsew signal output
rlabel metal2 s 221830 0 221886 800 6 la_data_out[68]
port 628 nsew signal output
rlabel metal2 s 223946 0 224002 800 6 la_data_out[69]
port 629 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[6]
port 630 nsew signal output
rlabel metal2 s 226062 0 226118 800 6 la_data_out[70]
port 631 nsew signal output
rlabel metal2 s 228270 0 228326 800 6 la_data_out[71]
port 632 nsew signal output
rlabel metal2 s 230386 0 230442 800 6 la_data_out[72]
port 633 nsew signal output
rlabel metal2 s 232502 0 232558 800 6 la_data_out[73]
port 634 nsew signal output
rlabel metal2 s 234618 0 234674 800 6 la_data_out[74]
port 635 nsew signal output
rlabel metal2 s 236826 0 236882 800 6 la_data_out[75]
port 636 nsew signal output
rlabel metal2 s 238942 0 238998 800 6 la_data_out[76]
port 637 nsew signal output
rlabel metal2 s 241058 0 241114 800 6 la_data_out[77]
port 638 nsew signal output
rlabel metal2 s 243174 0 243230 800 6 la_data_out[78]
port 639 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 la_data_out[79]
port 640 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[7]
port 641 nsew signal output
rlabel metal2 s 247498 0 247554 800 6 la_data_out[80]
port 642 nsew signal output
rlabel metal2 s 249614 0 249670 800 6 la_data_out[81]
port 643 nsew signal output
rlabel metal2 s 251730 0 251786 800 6 la_data_out[82]
port 644 nsew signal output
rlabel metal2 s 253938 0 253994 800 6 la_data_out[83]
port 645 nsew signal output
rlabel metal2 s 256054 0 256110 800 6 la_data_out[84]
port 646 nsew signal output
rlabel metal2 s 258170 0 258226 800 6 la_data_out[85]
port 647 nsew signal output
rlabel metal2 s 260286 0 260342 800 6 la_data_out[86]
port 648 nsew signal output
rlabel metal2 s 262402 0 262458 800 6 la_data_out[87]
port 649 nsew signal output
rlabel metal2 s 264610 0 264666 800 6 la_data_out[88]
port 650 nsew signal output
rlabel metal2 s 266726 0 266782 800 6 la_data_out[89]
port 651 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[8]
port 652 nsew signal output
rlabel metal2 s 268842 0 268898 800 6 la_data_out[90]
port 653 nsew signal output
rlabel metal2 s 270958 0 271014 800 6 la_data_out[91]
port 654 nsew signal output
rlabel metal2 s 273166 0 273222 800 6 la_data_out[92]
port 655 nsew signal output
rlabel metal2 s 275282 0 275338 800 6 la_data_out[93]
port 656 nsew signal output
rlabel metal2 s 277398 0 277454 800 6 la_data_out[94]
port 657 nsew signal output
rlabel metal2 s 279514 0 279570 800 6 la_data_out[95]
port 658 nsew signal output
rlabel metal2 s 281722 0 281778 800 6 la_data_out[96]
port 659 nsew signal output
rlabel metal2 s 283838 0 283894 800 6 la_data_out[97]
port 660 nsew signal output
rlabel metal2 s 285954 0 286010 800 6 la_data_out[98]
port 661 nsew signal output
rlabel metal2 s 288070 0 288126 800 6 la_data_out[99]
port 662 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_data_out[9]
port 663 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 la_oenb[0]
port 664 nsew signal input
rlabel metal2 s 290922 0 290978 800 6 la_oenb[100]
port 665 nsew signal input
rlabel metal2 s 293038 0 293094 800 6 la_oenb[101]
port 666 nsew signal input
rlabel metal2 s 295246 0 295302 800 6 la_oenb[102]
port 667 nsew signal input
rlabel metal2 s 297362 0 297418 800 6 la_oenb[103]
port 668 nsew signal input
rlabel metal2 s 299478 0 299534 800 6 la_oenb[104]
port 669 nsew signal input
rlabel metal2 s 301594 0 301650 800 6 la_oenb[105]
port 670 nsew signal input
rlabel metal2 s 303802 0 303858 800 6 la_oenb[106]
port 671 nsew signal input
rlabel metal2 s 305918 0 305974 800 6 la_oenb[107]
port 672 nsew signal input
rlabel metal2 s 308034 0 308090 800 6 la_oenb[108]
port 673 nsew signal input
rlabel metal2 s 310150 0 310206 800 6 la_oenb[109]
port 674 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_oenb[10]
port 675 nsew signal input
rlabel metal2 s 312358 0 312414 800 6 la_oenb[110]
port 676 nsew signal input
rlabel metal2 s 314474 0 314530 800 6 la_oenb[111]
port 677 nsew signal input
rlabel metal2 s 316590 0 316646 800 6 la_oenb[112]
port 678 nsew signal input
rlabel metal2 s 318706 0 318762 800 6 la_oenb[113]
port 679 nsew signal input
rlabel metal2 s 320822 0 320878 800 6 la_oenb[114]
port 680 nsew signal input
rlabel metal2 s 323030 0 323086 800 6 la_oenb[115]
port 681 nsew signal input
rlabel metal2 s 325146 0 325202 800 6 la_oenb[116]
port 682 nsew signal input
rlabel metal2 s 327262 0 327318 800 6 la_oenb[117]
port 683 nsew signal input
rlabel metal2 s 329378 0 329434 800 6 la_oenb[118]
port 684 nsew signal input
rlabel metal2 s 331586 0 331642 800 6 la_oenb[119]
port 685 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_oenb[11]
port 686 nsew signal input
rlabel metal2 s 333702 0 333758 800 6 la_oenb[120]
port 687 nsew signal input
rlabel metal2 s 335818 0 335874 800 6 la_oenb[121]
port 688 nsew signal input
rlabel metal2 s 337934 0 337990 800 6 la_oenb[122]
port 689 nsew signal input
rlabel metal2 s 340142 0 340198 800 6 la_oenb[123]
port 690 nsew signal input
rlabel metal2 s 342258 0 342314 800 6 la_oenb[124]
port 691 nsew signal input
rlabel metal2 s 344374 0 344430 800 6 la_oenb[125]
port 692 nsew signal input
rlabel metal2 s 346490 0 346546 800 6 la_oenb[126]
port 693 nsew signal input
rlabel metal2 s 348698 0 348754 800 6 la_oenb[127]
port 694 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[12]
port 695 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[13]
port 696 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_oenb[14]
port 697 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oenb[15]
port 698 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[16]
port 699 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_oenb[17]
port 700 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[18]
port 701 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[19]
port 702 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[1]
port 703 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_oenb[20]
port 704 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_oenb[21]
port 705 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_oenb[22]
port 706 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_oenb[23]
port 707 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_oenb[24]
port 708 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_oenb[25]
port 709 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_oenb[26]
port 710 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_oenb[27]
port 711 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[28]
port 712 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oenb[29]
port 713 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[2]
port 714 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[30]
port 715 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_oenb[31]
port 716 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[32]
port 717 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oenb[33]
port 718 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_oenb[34]
port 719 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_oenb[35]
port 720 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oenb[36]
port 721 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_oenb[37]
port 722 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oenb[38]
port 723 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oenb[39]
port 724 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[3]
port 725 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_oenb[40]
port 726 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 la_oenb[41]
port 727 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_oenb[42]
port 728 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_oenb[43]
port 729 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_oenb[44]
port 730 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 la_oenb[45]
port 731 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_oenb[46]
port 732 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oenb[47]
port 733 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_oenb[48]
port 734 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_oenb[49]
port 735 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[4]
port 736 nsew signal input
rlabel metal2 s 184110 0 184166 800 6 la_oenb[50]
port 737 nsew signal input
rlabel metal2 s 186226 0 186282 800 6 la_oenb[51]
port 738 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_oenb[52]
port 739 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 la_oenb[53]
port 740 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_oenb[54]
port 741 nsew signal input
rlabel metal2 s 194782 0 194838 800 6 la_oenb[55]
port 742 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_oenb[56]
port 743 nsew signal input
rlabel metal2 s 199014 0 199070 800 6 la_oenb[57]
port 744 nsew signal input
rlabel metal2 s 201130 0 201186 800 6 la_oenb[58]
port 745 nsew signal input
rlabel metal2 s 203338 0 203394 800 6 la_oenb[59]
port 746 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[5]
port 747 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_oenb[60]
port 748 nsew signal input
rlabel metal2 s 207570 0 207626 800 6 la_oenb[61]
port 749 nsew signal input
rlabel metal2 s 209686 0 209742 800 6 la_oenb[62]
port 750 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 la_oenb[63]
port 751 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 la_oenb[64]
port 752 nsew signal input
rlabel metal2 s 216126 0 216182 800 6 la_oenb[65]
port 753 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_oenb[66]
port 754 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_oenb[67]
port 755 nsew signal input
rlabel metal2 s 222566 0 222622 800 6 la_oenb[68]
port 756 nsew signal input
rlabel metal2 s 224682 0 224738 800 6 la_oenb[69]
port 757 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_oenb[6]
port 758 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_oenb[70]
port 759 nsew signal input
rlabel metal2 s 228914 0 228970 800 6 la_oenb[71]
port 760 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_oenb[72]
port 761 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_oenb[73]
port 762 nsew signal input
rlabel metal2 s 235354 0 235410 800 6 la_oenb[74]
port 763 nsew signal input
rlabel metal2 s 237470 0 237526 800 6 la_oenb[75]
port 764 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_oenb[76]
port 765 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_oenb[77]
port 766 nsew signal input
rlabel metal2 s 243910 0 243966 800 6 la_oenb[78]
port 767 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 la_oenb[79]
port 768 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[7]
port 769 nsew signal input
rlabel metal2 s 248234 0 248290 800 6 la_oenb[80]
port 770 nsew signal input
rlabel metal2 s 250350 0 250406 800 6 la_oenb[81]
port 771 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 la_oenb[82]
port 772 nsew signal input
rlabel metal2 s 254582 0 254638 800 6 la_oenb[83]
port 773 nsew signal input
rlabel metal2 s 256698 0 256754 800 6 la_oenb[84]
port 774 nsew signal input
rlabel metal2 s 258906 0 258962 800 6 la_oenb[85]
port 775 nsew signal input
rlabel metal2 s 261022 0 261078 800 6 la_oenb[86]
port 776 nsew signal input
rlabel metal2 s 263138 0 263194 800 6 la_oenb[87]
port 777 nsew signal input
rlabel metal2 s 265254 0 265310 800 6 la_oenb[88]
port 778 nsew signal input
rlabel metal2 s 267462 0 267518 800 6 la_oenb[89]
port 779 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_oenb[8]
port 780 nsew signal input
rlabel metal2 s 269578 0 269634 800 6 la_oenb[90]
port 781 nsew signal input
rlabel metal2 s 271694 0 271750 800 6 la_oenb[91]
port 782 nsew signal input
rlabel metal2 s 273810 0 273866 800 6 la_oenb[92]
port 783 nsew signal input
rlabel metal2 s 276018 0 276074 800 6 la_oenb[93]
port 784 nsew signal input
rlabel metal2 s 278134 0 278190 800 6 la_oenb[94]
port 785 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 la_oenb[95]
port 786 nsew signal input
rlabel metal2 s 282366 0 282422 800 6 la_oenb[96]
port 787 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 la_oenb[97]
port 788 nsew signal input
rlabel metal2 s 286690 0 286746 800 6 la_oenb[98]
port 789 nsew signal input
rlabel metal2 s 288806 0 288862 800 6 la_oenb[99]
port 790 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[9]
port 791 nsew signal input
rlabel metal2 s 118974 352563 119030 353363 6 tag_array_ext_ram_addr1[0]
port 792 nsew signal output
rlabel metal2 s 119986 352563 120042 353363 6 tag_array_ext_ram_addr1[1]
port 793 nsew signal output
rlabel metal2 s 121090 352563 121146 353363 6 tag_array_ext_ram_addr1[2]
port 794 nsew signal output
rlabel metal2 s 122102 352563 122158 353363 6 tag_array_ext_ram_addr1[3]
port 795 nsew signal output
rlabel metal2 s 123206 352563 123262 353363 6 tag_array_ext_ram_addr1[4]
port 796 nsew signal output
rlabel metal2 s 124310 352563 124366 353363 6 tag_array_ext_ram_addr1[5]
port 797 nsew signal output
rlabel metal2 s 125322 352563 125378 353363 6 tag_array_ext_ram_addr1[6]
port 798 nsew signal output
rlabel metal2 s 126426 352563 126482 353363 6 tag_array_ext_ram_addr1[7]
port 799 nsew signal output
rlabel metal2 s 34610 352563 34666 353363 6 tag_array_ext_ram_addr[0]
port 800 nsew signal output
rlabel metal2 s 35622 352563 35678 353363 6 tag_array_ext_ram_addr[1]
port 801 nsew signal output
rlabel metal2 s 36726 352563 36782 353363 6 tag_array_ext_ram_addr[2]
port 802 nsew signal output
rlabel metal2 s 37830 352563 37886 353363 6 tag_array_ext_ram_addr[3]
port 803 nsew signal output
rlabel metal2 s 38842 352563 38898 353363 6 tag_array_ext_ram_addr[4]
port 804 nsew signal output
rlabel metal2 s 39946 352563 40002 353363 6 tag_array_ext_ram_addr[5]
port 805 nsew signal output
rlabel metal2 s 40958 352563 41014 353363 6 tag_array_ext_ram_addr[6]
port 806 nsew signal output
rlabel metal2 s 42062 352563 42118 353363 6 tag_array_ext_ram_addr[7]
port 807 nsew signal output
rlabel metal2 s 43166 352563 43222 353363 6 tag_array_ext_ram_clk
port 808 nsew signal output
rlabel metal2 s 114650 352563 114706 353363 6 tag_array_ext_ram_csb
port 809 nsew signal output
rlabel metal2 s 116766 352563 116822 353363 6 tag_array_ext_ram_csb1[0]
port 810 nsew signal output
rlabel metal2 s 117870 352563 117926 353363 6 tag_array_ext_ram_csb1[1]
port 811 nsew signal output
rlabel metal2 s 478 352563 534 353363 6 tag_array_ext_ram_rdata0[0]
port 812 nsew signal input
rlabel metal2 s 11150 352563 11206 353363 6 tag_array_ext_ram_rdata0[10]
port 813 nsew signal input
rlabel metal2 s 12162 352563 12218 353363 6 tag_array_ext_ram_rdata0[11]
port 814 nsew signal input
rlabel metal2 s 13266 352563 13322 353363 6 tag_array_ext_ram_rdata0[12]
port 815 nsew signal input
rlabel metal2 s 14278 352563 14334 353363 6 tag_array_ext_ram_rdata0[13]
port 816 nsew signal input
rlabel metal2 s 15382 352563 15438 353363 6 tag_array_ext_ram_rdata0[14]
port 817 nsew signal input
rlabel metal2 s 16486 352563 16542 353363 6 tag_array_ext_ram_rdata0[15]
port 818 nsew signal input
rlabel metal2 s 17498 352563 17554 353363 6 tag_array_ext_ram_rdata0[16]
port 819 nsew signal input
rlabel metal2 s 18602 352563 18658 353363 6 tag_array_ext_ram_rdata0[17]
port 820 nsew signal input
rlabel metal2 s 19614 352563 19670 353363 6 tag_array_ext_ram_rdata0[18]
port 821 nsew signal input
rlabel metal2 s 20718 352563 20774 353363 6 tag_array_ext_ram_rdata0[19]
port 822 nsew signal input
rlabel metal2 s 1490 352563 1546 353363 6 tag_array_ext_ram_rdata0[1]
port 823 nsew signal input
rlabel metal2 s 21822 352563 21878 353363 6 tag_array_ext_ram_rdata0[20]
port 824 nsew signal input
rlabel metal2 s 22834 352563 22890 353363 6 tag_array_ext_ram_rdata0[21]
port 825 nsew signal input
rlabel metal2 s 23938 352563 23994 353363 6 tag_array_ext_ram_rdata0[22]
port 826 nsew signal input
rlabel metal2 s 24950 352563 25006 353363 6 tag_array_ext_ram_rdata0[23]
port 827 nsew signal input
rlabel metal2 s 26054 352563 26110 353363 6 tag_array_ext_ram_rdata0[24]
port 828 nsew signal input
rlabel metal2 s 27158 352563 27214 353363 6 tag_array_ext_ram_rdata0[25]
port 829 nsew signal input
rlabel metal2 s 28170 352563 28226 353363 6 tag_array_ext_ram_rdata0[26]
port 830 nsew signal input
rlabel metal2 s 29274 352563 29330 353363 6 tag_array_ext_ram_rdata0[27]
port 831 nsew signal input
rlabel metal2 s 30286 352563 30342 353363 6 tag_array_ext_ram_rdata0[28]
port 832 nsew signal input
rlabel metal2 s 31390 352563 31446 353363 6 tag_array_ext_ram_rdata0[29]
port 833 nsew signal input
rlabel metal2 s 2594 352563 2650 353363 6 tag_array_ext_ram_rdata0[2]
port 834 nsew signal input
rlabel metal2 s 32494 352563 32550 353363 6 tag_array_ext_ram_rdata0[30]
port 835 nsew signal input
rlabel metal2 s 33506 352563 33562 353363 6 tag_array_ext_ram_rdata0[31]
port 836 nsew signal input
rlabel metal2 s 3606 352563 3662 353363 6 tag_array_ext_ram_rdata0[3]
port 837 nsew signal input
rlabel metal2 s 4710 352563 4766 353363 6 tag_array_ext_ram_rdata0[4]
port 838 nsew signal input
rlabel metal2 s 5814 352563 5870 353363 6 tag_array_ext_ram_rdata0[5]
port 839 nsew signal input
rlabel metal2 s 6826 352563 6882 353363 6 tag_array_ext_ram_rdata0[6]
port 840 nsew signal input
rlabel metal2 s 7930 352563 7986 353363 6 tag_array_ext_ram_rdata0[7]
port 841 nsew signal input
rlabel metal2 s 8942 352563 8998 353363 6 tag_array_ext_ram_rdata0[8]
port 842 nsew signal input
rlabel metal2 s 10046 352563 10102 353363 6 tag_array_ext_ram_rdata0[9]
port 843 nsew signal input
rlabel metal2 s 127438 352563 127494 353363 6 tag_array_ext_ram_rdata1[0]
port 844 nsew signal input
rlabel metal2 s 138202 352563 138258 353363 6 tag_array_ext_ram_rdata1[10]
port 845 nsew signal input
rlabel metal2 s 139214 352563 139270 353363 6 tag_array_ext_ram_rdata1[11]
port 846 nsew signal input
rlabel metal2 s 140318 352563 140374 353363 6 tag_array_ext_ram_rdata1[12]
port 847 nsew signal input
rlabel metal2 s 141330 352563 141386 353363 6 tag_array_ext_ram_rdata1[13]
port 848 nsew signal input
rlabel metal2 s 142434 352563 142490 353363 6 tag_array_ext_ram_rdata1[14]
port 849 nsew signal input
rlabel metal2 s 143538 352563 143594 353363 6 tag_array_ext_ram_rdata1[15]
port 850 nsew signal input
rlabel metal2 s 144550 352563 144606 353363 6 tag_array_ext_ram_rdata1[16]
port 851 nsew signal input
rlabel metal2 s 145654 352563 145710 353363 6 tag_array_ext_ram_rdata1[17]
port 852 nsew signal input
rlabel metal2 s 146666 352563 146722 353363 6 tag_array_ext_ram_rdata1[18]
port 853 nsew signal input
rlabel metal2 s 147770 352563 147826 353363 6 tag_array_ext_ram_rdata1[19]
port 854 nsew signal input
rlabel metal2 s 128542 352563 128598 353363 6 tag_array_ext_ram_rdata1[1]
port 855 nsew signal input
rlabel metal2 s 148874 352563 148930 353363 6 tag_array_ext_ram_rdata1[20]
port 856 nsew signal input
rlabel metal2 s 149886 352563 149942 353363 6 tag_array_ext_ram_rdata1[21]
port 857 nsew signal input
rlabel metal2 s 150990 352563 151046 353363 6 tag_array_ext_ram_rdata1[22]
port 858 nsew signal input
rlabel metal2 s 152002 352563 152058 353363 6 tag_array_ext_ram_rdata1[23]
port 859 nsew signal input
rlabel metal2 s 153106 352563 153162 353363 6 tag_array_ext_ram_rdata1[24]
port 860 nsew signal input
rlabel metal2 s 154210 352563 154266 353363 6 tag_array_ext_ram_rdata1[25]
port 861 nsew signal input
rlabel metal2 s 155222 352563 155278 353363 6 tag_array_ext_ram_rdata1[26]
port 862 nsew signal input
rlabel metal2 s 156326 352563 156382 353363 6 tag_array_ext_ram_rdata1[27]
port 863 nsew signal input
rlabel metal2 s 157338 352563 157394 353363 6 tag_array_ext_ram_rdata1[28]
port 864 nsew signal input
rlabel metal2 s 158442 352563 158498 353363 6 tag_array_ext_ram_rdata1[29]
port 865 nsew signal input
rlabel metal2 s 129646 352563 129702 353363 6 tag_array_ext_ram_rdata1[2]
port 866 nsew signal input
rlabel metal2 s 159546 352563 159602 353363 6 tag_array_ext_ram_rdata1[30]
port 867 nsew signal input
rlabel metal2 s 160558 352563 160614 353363 6 tag_array_ext_ram_rdata1[31]
port 868 nsew signal input
rlabel metal2 s 130658 352563 130714 353363 6 tag_array_ext_ram_rdata1[3]
port 869 nsew signal input
rlabel metal2 s 131762 352563 131818 353363 6 tag_array_ext_ram_rdata1[4]
port 870 nsew signal input
rlabel metal2 s 132866 352563 132922 353363 6 tag_array_ext_ram_rdata1[5]
port 871 nsew signal input
rlabel metal2 s 133878 352563 133934 353363 6 tag_array_ext_ram_rdata1[6]
port 872 nsew signal input
rlabel metal2 s 134982 352563 135038 353363 6 tag_array_ext_ram_rdata1[7]
port 873 nsew signal input
rlabel metal2 s 135994 352563 136050 353363 6 tag_array_ext_ram_rdata1[8]
port 874 nsew signal input
rlabel metal2 s 137098 352563 137154 353363 6 tag_array_ext_ram_rdata1[9]
port 875 nsew signal input
rlabel metal2 s 44178 352563 44234 353363 6 tag_array_ext_ram_wdata[0]
port 876 nsew signal output
rlabel metal2 s 54850 352563 54906 353363 6 tag_array_ext_ram_wdata[10]
port 877 nsew signal output
rlabel metal2 s 55954 352563 56010 353363 6 tag_array_ext_ram_wdata[11]
port 878 nsew signal output
rlabel metal2 s 57058 352563 57114 353363 6 tag_array_ext_ram_wdata[12]
port 879 nsew signal output
rlabel metal2 s 58070 352563 58126 353363 6 tag_array_ext_ram_wdata[13]
port 880 nsew signal output
rlabel metal2 s 59174 352563 59230 353363 6 tag_array_ext_ram_wdata[14]
port 881 nsew signal output
rlabel metal2 s 60186 352563 60242 353363 6 tag_array_ext_ram_wdata[15]
port 882 nsew signal output
rlabel metal2 s 61290 352563 61346 353363 6 tag_array_ext_ram_wdata[16]
port 883 nsew signal output
rlabel metal2 s 62394 352563 62450 353363 6 tag_array_ext_ram_wdata[17]
port 884 nsew signal output
rlabel metal2 s 63406 352563 63462 353363 6 tag_array_ext_ram_wdata[18]
port 885 nsew signal output
rlabel metal2 s 64510 352563 64566 353363 6 tag_array_ext_ram_wdata[19]
port 886 nsew signal output
rlabel metal2 s 45282 352563 45338 353363 6 tag_array_ext_ram_wdata[1]
port 887 nsew signal output
rlabel metal2 s 65522 352563 65578 353363 6 tag_array_ext_ram_wdata[20]
port 888 nsew signal output
rlabel metal2 s 66626 352563 66682 353363 6 tag_array_ext_ram_wdata[21]
port 889 nsew signal output
rlabel metal2 s 67730 352563 67786 353363 6 tag_array_ext_ram_wdata[22]
port 890 nsew signal output
rlabel metal2 s 68742 352563 68798 353363 6 tag_array_ext_ram_wdata[23]
port 891 nsew signal output
rlabel metal2 s 69846 352563 69902 353363 6 tag_array_ext_ram_wdata[24]
port 892 nsew signal output
rlabel metal2 s 70858 352563 70914 353363 6 tag_array_ext_ram_wdata[25]
port 893 nsew signal output
rlabel metal2 s 71962 352563 72018 353363 6 tag_array_ext_ram_wdata[26]
port 894 nsew signal output
rlabel metal2 s 73066 352563 73122 353363 6 tag_array_ext_ram_wdata[27]
port 895 nsew signal output
rlabel metal2 s 74078 352563 74134 353363 6 tag_array_ext_ram_wdata[28]
port 896 nsew signal output
rlabel metal2 s 75182 352563 75238 353363 6 tag_array_ext_ram_wdata[29]
port 897 nsew signal output
rlabel metal2 s 46386 352563 46442 353363 6 tag_array_ext_ram_wdata[2]
port 898 nsew signal output
rlabel metal2 s 76194 352563 76250 353363 6 tag_array_ext_ram_wdata[30]
port 899 nsew signal output
rlabel metal2 s 77298 352563 77354 353363 6 tag_array_ext_ram_wdata[31]
port 900 nsew signal output
rlabel metal2 s 78402 352563 78458 353363 6 tag_array_ext_ram_wdata[32]
port 901 nsew signal output
rlabel metal2 s 79414 352563 79470 353363 6 tag_array_ext_ram_wdata[33]
port 902 nsew signal output
rlabel metal2 s 80518 352563 80574 353363 6 tag_array_ext_ram_wdata[34]
port 903 nsew signal output
rlabel metal2 s 81530 352563 81586 353363 6 tag_array_ext_ram_wdata[35]
port 904 nsew signal output
rlabel metal2 s 82634 352563 82690 353363 6 tag_array_ext_ram_wdata[36]
port 905 nsew signal output
rlabel metal2 s 83738 352563 83794 353363 6 tag_array_ext_ram_wdata[37]
port 906 nsew signal output
rlabel metal2 s 84750 352563 84806 353363 6 tag_array_ext_ram_wdata[38]
port 907 nsew signal output
rlabel metal2 s 85854 352563 85910 353363 6 tag_array_ext_ram_wdata[39]
port 908 nsew signal output
rlabel metal2 s 47398 352563 47454 353363 6 tag_array_ext_ram_wdata[3]
port 909 nsew signal output
rlabel metal2 s 86866 352563 86922 353363 6 tag_array_ext_ram_wdata[40]
port 910 nsew signal output
rlabel metal2 s 87970 352563 88026 353363 6 tag_array_ext_ram_wdata[41]
port 911 nsew signal output
rlabel metal2 s 89074 352563 89130 353363 6 tag_array_ext_ram_wdata[42]
port 912 nsew signal output
rlabel metal2 s 90086 352563 90142 353363 6 tag_array_ext_ram_wdata[43]
port 913 nsew signal output
rlabel metal2 s 91190 352563 91246 353363 6 tag_array_ext_ram_wdata[44]
port 914 nsew signal output
rlabel metal2 s 92294 352563 92350 353363 6 tag_array_ext_ram_wdata[45]
port 915 nsew signal output
rlabel metal2 s 93306 352563 93362 353363 6 tag_array_ext_ram_wdata[46]
port 916 nsew signal output
rlabel metal2 s 94410 352563 94466 353363 6 tag_array_ext_ram_wdata[47]
port 917 nsew signal output
rlabel metal2 s 95422 352563 95478 353363 6 tag_array_ext_ram_wdata[48]
port 918 nsew signal output
rlabel metal2 s 96526 352563 96582 353363 6 tag_array_ext_ram_wdata[49]
port 919 nsew signal output
rlabel metal2 s 48502 352563 48558 353363 6 tag_array_ext_ram_wdata[4]
port 920 nsew signal output
rlabel metal2 s 97630 352563 97686 353363 6 tag_array_ext_ram_wdata[50]
port 921 nsew signal output
rlabel metal2 s 98642 352563 98698 353363 6 tag_array_ext_ram_wdata[51]
port 922 nsew signal output
rlabel metal2 s 99746 352563 99802 353363 6 tag_array_ext_ram_wdata[52]
port 923 nsew signal output
rlabel metal2 s 100758 352563 100814 353363 6 tag_array_ext_ram_wdata[53]
port 924 nsew signal output
rlabel metal2 s 101862 352563 101918 353363 6 tag_array_ext_ram_wdata[54]
port 925 nsew signal output
rlabel metal2 s 102966 352563 103022 353363 6 tag_array_ext_ram_wdata[55]
port 926 nsew signal output
rlabel metal2 s 103978 352563 104034 353363 6 tag_array_ext_ram_wdata[56]
port 927 nsew signal output
rlabel metal2 s 105082 352563 105138 353363 6 tag_array_ext_ram_wdata[57]
port 928 nsew signal output
rlabel metal2 s 106094 352563 106150 353363 6 tag_array_ext_ram_wdata[58]
port 929 nsew signal output
rlabel metal2 s 107198 352563 107254 353363 6 tag_array_ext_ram_wdata[59]
port 930 nsew signal output
rlabel metal2 s 49514 352563 49570 353363 6 tag_array_ext_ram_wdata[5]
port 931 nsew signal output
rlabel metal2 s 108302 352563 108358 353363 6 tag_array_ext_ram_wdata[60]
port 932 nsew signal output
rlabel metal2 s 109314 352563 109370 353363 6 tag_array_ext_ram_wdata[61]
port 933 nsew signal output
rlabel metal2 s 110418 352563 110474 353363 6 tag_array_ext_ram_wdata[62]
port 934 nsew signal output
rlabel metal2 s 111430 352563 111486 353363 6 tag_array_ext_ram_wdata[63]
port 935 nsew signal output
rlabel metal2 s 50618 352563 50674 353363 6 tag_array_ext_ram_wdata[6]
port 936 nsew signal output
rlabel metal2 s 51722 352563 51778 353363 6 tag_array_ext_ram_wdata[7]
port 937 nsew signal output
rlabel metal2 s 52734 352563 52790 353363 6 tag_array_ext_ram_wdata[8]
port 938 nsew signal output
rlabel metal2 s 53838 352563 53894 353363 6 tag_array_ext_ram_wdata[9]
port 939 nsew signal output
rlabel metal2 s 115754 352563 115810 353363 6 tag_array_ext_ram_web
port 940 nsew signal output
rlabel metal2 s 112534 352563 112590 353363 6 tag_array_ext_ram_wmask[0]
port 941 nsew signal output
rlabel metal2 s 113638 352563 113694 353363 6 tag_array_ext_ram_wmask[1]
port 942 nsew signal output
rlabel metal4 s 4208 2128 4528 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 34928 2128 35248 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 65648 2128 65968 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 96368 2128 96688 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 127088 2128 127408 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 157808 2128 158128 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 188528 2128 188848 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 219248 2128 219568 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 249968 2128 250288 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 280688 2128 281008 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 311408 2128 311728 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 342128 2128 342448 350928 6 vccd1
port 943 nsew power input
rlabel metal4 s 19568 2128 19888 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 50288 2128 50608 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 81008 2128 81328 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 111728 2128 112048 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 142448 2128 142768 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 173168 2128 173488 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 203888 2128 204208 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 234608 2128 234928 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 265328 2128 265648 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 296048 2128 296368 350928 6 vssd1
port 944 nsew ground input
rlabel metal4 s 326768 2128 327088 350928 6 vssd1
port 944 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 945 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 946 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_ack_o
port 947 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[0]
port 948 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[10]
port 949 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[11]
port 950 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[12]
port 951 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_adr_i[13]
port 952 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[14]
port 953 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_adr_i[15]
port 954 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_adr_i[16]
port 955 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[17]
port 956 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_adr_i[18]
port 957 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 wbs_adr_i[19]
port 958 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[1]
port 959 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[20]
port 960 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 wbs_adr_i[21]
port 961 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_adr_i[22]
port 962 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_adr_i[23]
port 963 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_adr_i[24]
port 964 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_adr_i[25]
port 965 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 wbs_adr_i[26]
port 966 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_adr_i[27]
port 967 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 wbs_adr_i[28]
port 968 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 wbs_adr_i[29]
port 969 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[2]
port 970 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 wbs_adr_i[30]
port 971 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 wbs_adr_i[31]
port 972 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[3]
port 973 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[4]
port 974 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[5]
port 975 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[6]
port 976 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_adr_i[7]
port 977 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[8]
port 978 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_adr_i[9]
port 979 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_cyc_i
port 980 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_i[0]
port 981 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[10]
port 982 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[11]
port 983 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[12]
port 984 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_i[13]
port 985 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[14]
port 986 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[15]
port 987 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 wbs_dat_i[16]
port 988 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_dat_i[17]
port 989 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_i[18]
port 990 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_dat_i[19]
port 991 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[1]
port 992 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[20]
port 993 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_i[21]
port 994 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[22]
port 995 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_i[23]
port 996 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 wbs_dat_i[24]
port 997 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_dat_i[25]
port 998 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 wbs_dat_i[26]
port 999 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_i[27]
port 1000 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 wbs_dat_i[28]
port 1001 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 wbs_dat_i[29]
port 1002 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[2]
port 1003 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 wbs_dat_i[30]
port 1004 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 wbs_dat_i[31]
port 1005 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[3]
port 1006 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[4]
port 1007 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[5]
port 1008 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_i[6]
port 1009 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[7]
port 1010 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[8]
port 1011 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_i[9]
port 1012 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[0]
port 1013 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_o[10]
port 1014 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[11]
port 1015 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[12]
port 1016 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_o[13]
port 1017 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_o[14]
port 1018 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[15]
port 1019 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[16]
port 1020 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_o[17]
port 1021 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_o[18]
port 1022 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_o[19]
port 1023 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[1]
port 1024 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_o[20]
port 1025 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 wbs_dat_o[21]
port 1026 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 wbs_dat_o[22]
port 1027 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_o[23]
port 1028 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_o[24]
port 1029 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 wbs_dat_o[25]
port 1030 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 wbs_dat_o[26]
port 1031 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 wbs_dat_o[27]
port 1032 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 wbs_dat_o[28]
port 1033 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 wbs_dat_o[29]
port 1034 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[2]
port 1035 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 wbs_dat_o[30]
port 1036 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 wbs_dat_o[31]
port 1037 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[3]
port 1038 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[4]
port 1039 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[5]
port 1040 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[6]
port 1041 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_o[7]
port 1042 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[8]
port 1043 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_o[9]
port 1044 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_sel_i[0]
port 1045 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_sel_i[1]
port 1046 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_sel_i[2]
port 1047 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_sel_i[3]
port 1048 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_stb_i
port 1049 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_we_i
port 1050 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 351219 353363
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 310714600
string GDS_FILE /home/shc/Development/efabless/marmot_asic/openlane/marmot/runs/marmot/results/finishing/Marmot.magic.gds
string GDS_START 1960534
<< end >>

