magic
tech sky130A
magscale 1 2
timestamp 1647805847
<< obsli1 >>
rect 1104 2159 352360 353073
<< obsm1 >>
rect 198 8 353450 354748
<< metal2 >>
rect 1490 354823 1546 355623
rect 4526 354823 4582 355623
rect 7654 354823 7710 355623
rect 10782 354823 10838 355623
rect 13818 354823 13874 355623
rect 16946 354823 17002 355623
rect 20074 354823 20130 355623
rect 23110 354823 23166 355623
rect 26238 354823 26294 355623
rect 29366 354823 29422 355623
rect 32494 354823 32550 355623
rect 35530 354823 35586 355623
rect 38658 354823 38714 355623
rect 41786 354823 41842 355623
rect 44822 354823 44878 355623
rect 47950 354823 48006 355623
rect 51078 354823 51134 355623
rect 54114 354823 54170 355623
rect 57242 354823 57298 355623
rect 60370 354823 60426 355623
rect 63498 354823 63554 355623
rect 66534 354823 66590 355623
rect 69662 354823 69718 355623
rect 72790 354823 72846 355623
rect 75826 354823 75882 355623
rect 78954 354823 79010 355623
rect 82082 354823 82138 355623
rect 85118 354823 85174 355623
rect 88246 354823 88302 355623
rect 91374 354823 91430 355623
rect 94502 354823 94558 355623
rect 97538 354823 97594 355623
rect 100666 354823 100722 355623
rect 103794 354823 103850 355623
rect 106830 354823 106886 355623
rect 109958 354823 110014 355623
rect 113086 354823 113142 355623
rect 116122 354823 116178 355623
rect 119250 354823 119306 355623
rect 122378 354823 122434 355623
rect 125506 354823 125562 355623
rect 128542 354823 128598 355623
rect 131670 354823 131726 355623
rect 134798 354823 134854 355623
rect 137834 354823 137890 355623
rect 140962 354823 141018 355623
rect 144090 354823 144146 355623
rect 147126 354823 147182 355623
rect 150254 354823 150310 355623
rect 153382 354823 153438 355623
rect 156510 354823 156566 355623
rect 159546 354823 159602 355623
rect 162674 354823 162730 355623
rect 165802 354823 165858 355623
rect 168838 354823 168894 355623
rect 171966 354823 172022 355623
rect 175094 354823 175150 355623
rect 178222 354823 178278 355623
rect 181258 354823 181314 355623
rect 184386 354823 184442 355623
rect 187514 354823 187570 355623
rect 190550 354823 190606 355623
rect 193678 354823 193734 355623
rect 196806 354823 196862 355623
rect 199842 354823 199898 355623
rect 202970 354823 203026 355623
rect 206098 354823 206154 355623
rect 209226 354823 209282 355623
rect 212262 354823 212318 355623
rect 215390 354823 215446 355623
rect 218518 354823 218574 355623
rect 221554 354823 221610 355623
rect 224682 354823 224738 355623
rect 227810 354823 227866 355623
rect 230846 354823 230902 355623
rect 233974 354823 234030 355623
rect 237102 354823 237158 355623
rect 240230 354823 240286 355623
rect 243266 354823 243322 355623
rect 246394 354823 246450 355623
rect 249522 354823 249578 355623
rect 252558 354823 252614 355623
rect 255686 354823 255742 355623
rect 258814 354823 258870 355623
rect 261850 354823 261906 355623
rect 264978 354823 265034 355623
rect 268106 354823 268162 355623
rect 271234 354823 271290 355623
rect 274270 354823 274326 355623
rect 277398 354823 277454 355623
rect 280526 354823 280582 355623
rect 283562 354823 283618 355623
rect 286690 354823 286746 355623
rect 289818 354823 289874 355623
rect 292854 354823 292910 355623
rect 295982 354823 296038 355623
rect 299110 354823 299166 355623
rect 302238 354823 302294 355623
rect 305274 354823 305330 355623
rect 308402 354823 308458 355623
rect 311530 354823 311586 355623
rect 314566 354823 314622 355623
rect 317694 354823 317750 355623
rect 320822 354823 320878 355623
rect 323858 354823 323914 355623
rect 326986 354823 327042 355623
rect 330114 354823 330170 355623
rect 333242 354823 333298 355623
rect 336278 354823 336334 355623
rect 339406 354823 339462 355623
rect 342534 354823 342590 355623
rect 345570 354823 345626 355623
rect 348698 354823 348754 355623
rect 351826 354823 351882 355623
rect 294 0 350 800
rect 938 0 994 800
rect 1674 0 1730 800
rect 2410 0 2466 800
rect 3146 0 3202 800
rect 3790 0 3846 800
rect 4526 0 4582 800
rect 5262 0 5318 800
rect 5998 0 6054 800
rect 6734 0 6790 800
rect 7378 0 7434 800
rect 8114 0 8170 800
rect 8850 0 8906 800
rect 9586 0 9642 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11702 0 11758 800
rect 12438 0 12494 800
rect 13174 0 13230 800
rect 13910 0 13966 800
rect 14554 0 14610 800
rect 15290 0 15346 800
rect 16026 0 16082 800
rect 16762 0 16818 800
rect 17498 0 17554 800
rect 18142 0 18198 800
rect 18878 0 18934 800
rect 19614 0 19670 800
rect 20350 0 20406 800
rect 21086 0 21142 800
rect 21730 0 21786 800
rect 22466 0 22522 800
rect 23202 0 23258 800
rect 23938 0 23994 800
rect 24582 0 24638 800
rect 25318 0 25374 800
rect 26054 0 26110 800
rect 26790 0 26846 800
rect 27526 0 27582 800
rect 28170 0 28226 800
rect 28906 0 28962 800
rect 29642 0 29698 800
rect 30378 0 30434 800
rect 31114 0 31170 800
rect 31758 0 31814 800
rect 32494 0 32550 800
rect 33230 0 33286 800
rect 33966 0 34022 800
rect 34702 0 34758 800
rect 35346 0 35402 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37554 0 37610 800
rect 38290 0 38346 800
rect 38934 0 38990 800
rect 39670 0 39726 800
rect 40406 0 40462 800
rect 41142 0 41198 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43258 0 43314 800
rect 43994 0 44050 800
rect 44730 0 44786 800
rect 45374 0 45430 800
rect 46110 0 46166 800
rect 46846 0 46902 800
rect 47582 0 47638 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49698 0 49754 800
rect 50434 0 50490 800
rect 51170 0 51226 800
rect 51906 0 51962 800
rect 52550 0 52606 800
rect 53286 0 53342 800
rect 54022 0 54078 800
rect 54758 0 54814 800
rect 55494 0 55550 800
rect 56138 0 56194 800
rect 56874 0 56930 800
rect 57610 0 57666 800
rect 58346 0 58402 800
rect 59082 0 59138 800
rect 59726 0 59782 800
rect 60462 0 60518 800
rect 61198 0 61254 800
rect 61934 0 61990 800
rect 62670 0 62726 800
rect 63314 0 63370 800
rect 64050 0 64106 800
rect 64786 0 64842 800
rect 65522 0 65578 800
rect 66166 0 66222 800
rect 66902 0 66958 800
rect 67638 0 67694 800
rect 68374 0 68430 800
rect 69110 0 69166 800
rect 69754 0 69810 800
rect 70490 0 70546 800
rect 71226 0 71282 800
rect 71962 0 72018 800
rect 72698 0 72754 800
rect 73342 0 73398 800
rect 74078 0 74134 800
rect 74814 0 74870 800
rect 75550 0 75606 800
rect 76286 0 76342 800
rect 76930 0 76986 800
rect 77666 0 77722 800
rect 78402 0 78458 800
rect 79138 0 79194 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81254 0 81310 800
rect 81990 0 82046 800
rect 82726 0 82782 800
rect 83462 0 83518 800
rect 84106 0 84162 800
rect 84842 0 84898 800
rect 85578 0 85634 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 87694 0 87750 800
rect 88430 0 88486 800
rect 89166 0 89222 800
rect 89902 0 89958 800
rect 90546 0 90602 800
rect 91282 0 91338 800
rect 92018 0 92074 800
rect 92754 0 92810 800
rect 93490 0 93546 800
rect 94134 0 94190 800
rect 94870 0 94926 800
rect 95606 0 95662 800
rect 96342 0 96398 800
rect 97078 0 97134 800
rect 97722 0 97778 800
rect 98458 0 98514 800
rect 99194 0 99250 800
rect 99930 0 99986 800
rect 100666 0 100722 800
rect 101310 0 101366 800
rect 102046 0 102102 800
rect 102782 0 102838 800
rect 103518 0 103574 800
rect 104254 0 104310 800
rect 104898 0 104954 800
rect 105634 0 105690 800
rect 106370 0 106426 800
rect 107106 0 107162 800
rect 107750 0 107806 800
rect 108486 0 108542 800
rect 109222 0 109278 800
rect 109958 0 110014 800
rect 110694 0 110750 800
rect 111338 0 111394 800
rect 112074 0 112130 800
rect 112810 0 112866 800
rect 113546 0 113602 800
rect 114282 0 114338 800
rect 114926 0 114982 800
rect 115662 0 115718 800
rect 116398 0 116454 800
rect 117134 0 117190 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119250 0 119306 800
rect 119986 0 120042 800
rect 120722 0 120778 800
rect 121458 0 121514 800
rect 122102 0 122158 800
rect 122838 0 122894 800
rect 123574 0 123630 800
rect 124310 0 124366 800
rect 125046 0 125102 800
rect 125690 0 125746 800
rect 126426 0 126482 800
rect 127162 0 127218 800
rect 127898 0 127954 800
rect 128542 0 128598 800
rect 129278 0 129334 800
rect 130014 0 130070 800
rect 130750 0 130806 800
rect 131486 0 131542 800
rect 132130 0 132186 800
rect 132866 0 132922 800
rect 133602 0 133658 800
rect 134338 0 134394 800
rect 135074 0 135130 800
rect 135718 0 135774 800
rect 136454 0 136510 800
rect 137190 0 137246 800
rect 137926 0 137982 800
rect 138662 0 138718 800
rect 139306 0 139362 800
rect 140042 0 140098 800
rect 140778 0 140834 800
rect 141514 0 141570 800
rect 142250 0 142306 800
rect 142894 0 142950 800
rect 143630 0 143686 800
rect 144366 0 144422 800
rect 145102 0 145158 800
rect 145838 0 145894 800
rect 146482 0 146538 800
rect 147218 0 147274 800
rect 147954 0 148010 800
rect 148690 0 148746 800
rect 149334 0 149390 800
rect 150070 0 150126 800
rect 150806 0 150862 800
rect 151542 0 151598 800
rect 152278 0 152334 800
rect 152922 0 152978 800
rect 153658 0 153714 800
rect 154394 0 154450 800
rect 155130 0 155186 800
rect 155866 0 155922 800
rect 156510 0 156566 800
rect 157246 0 157302 800
rect 157982 0 158038 800
rect 158718 0 158774 800
rect 159454 0 159510 800
rect 160098 0 160154 800
rect 160834 0 160890 800
rect 161570 0 161626 800
rect 162306 0 162362 800
rect 163042 0 163098 800
rect 163686 0 163742 800
rect 164422 0 164478 800
rect 165158 0 165214 800
rect 165894 0 165950 800
rect 166630 0 166686 800
rect 167274 0 167330 800
rect 168010 0 168066 800
rect 168746 0 168802 800
rect 169482 0 169538 800
rect 170126 0 170182 800
rect 170862 0 170918 800
rect 171598 0 171654 800
rect 172334 0 172390 800
rect 173070 0 173126 800
rect 173714 0 173770 800
rect 174450 0 174506 800
rect 175186 0 175242 800
rect 175922 0 175978 800
rect 176658 0 176714 800
rect 177302 0 177358 800
rect 178038 0 178094 800
rect 178774 0 178830 800
rect 179510 0 179566 800
rect 180246 0 180302 800
rect 180890 0 180946 800
rect 181626 0 181682 800
rect 182362 0 182418 800
rect 183098 0 183154 800
rect 183834 0 183890 800
rect 184478 0 184534 800
rect 185214 0 185270 800
rect 185950 0 186006 800
rect 186686 0 186742 800
rect 187422 0 187478 800
rect 188066 0 188122 800
rect 188802 0 188858 800
rect 189538 0 189594 800
rect 190274 0 190330 800
rect 190918 0 190974 800
rect 191654 0 191710 800
rect 192390 0 192446 800
rect 193126 0 193182 800
rect 193862 0 193918 800
rect 194506 0 194562 800
rect 195242 0 195298 800
rect 195978 0 196034 800
rect 196714 0 196770 800
rect 197450 0 197506 800
rect 198094 0 198150 800
rect 198830 0 198886 800
rect 199566 0 199622 800
rect 200302 0 200358 800
rect 201038 0 201094 800
rect 201682 0 201738 800
rect 202418 0 202474 800
rect 203154 0 203210 800
rect 203890 0 203946 800
rect 204626 0 204682 800
rect 205270 0 205326 800
rect 206006 0 206062 800
rect 206742 0 206798 800
rect 207478 0 207534 800
rect 208214 0 208270 800
rect 208858 0 208914 800
rect 209594 0 209650 800
rect 210330 0 210386 800
rect 211066 0 211122 800
rect 211710 0 211766 800
rect 212446 0 212502 800
rect 213182 0 213238 800
rect 213918 0 213974 800
rect 214654 0 214710 800
rect 215298 0 215354 800
rect 216034 0 216090 800
rect 216770 0 216826 800
rect 217506 0 217562 800
rect 218242 0 218298 800
rect 218886 0 218942 800
rect 219622 0 219678 800
rect 220358 0 220414 800
rect 221094 0 221150 800
rect 221830 0 221886 800
rect 222474 0 222530 800
rect 223210 0 223266 800
rect 223946 0 224002 800
rect 224682 0 224738 800
rect 225418 0 225474 800
rect 226062 0 226118 800
rect 226798 0 226854 800
rect 227534 0 227590 800
rect 228270 0 228326 800
rect 229006 0 229062 800
rect 229650 0 229706 800
rect 230386 0 230442 800
rect 231122 0 231178 800
rect 231858 0 231914 800
rect 232502 0 232558 800
rect 233238 0 233294 800
rect 233974 0 234030 800
rect 234710 0 234766 800
rect 235446 0 235502 800
rect 236090 0 236146 800
rect 236826 0 236882 800
rect 237562 0 237618 800
rect 238298 0 238354 800
rect 239034 0 239090 800
rect 239678 0 239734 800
rect 240414 0 240470 800
rect 241150 0 241206 800
rect 241886 0 241942 800
rect 242622 0 242678 800
rect 243266 0 243322 800
rect 244002 0 244058 800
rect 244738 0 244794 800
rect 245474 0 245530 800
rect 246210 0 246266 800
rect 246854 0 246910 800
rect 247590 0 247646 800
rect 248326 0 248382 800
rect 249062 0 249118 800
rect 249798 0 249854 800
rect 250442 0 250498 800
rect 251178 0 251234 800
rect 251914 0 251970 800
rect 252650 0 252706 800
rect 253294 0 253350 800
rect 254030 0 254086 800
rect 254766 0 254822 800
rect 255502 0 255558 800
rect 256238 0 256294 800
rect 256882 0 256938 800
rect 257618 0 257674 800
rect 258354 0 258410 800
rect 259090 0 259146 800
rect 259826 0 259882 800
rect 260470 0 260526 800
rect 261206 0 261262 800
rect 261942 0 261998 800
rect 262678 0 262734 800
rect 263414 0 263470 800
rect 264058 0 264114 800
rect 264794 0 264850 800
rect 265530 0 265586 800
rect 266266 0 266322 800
rect 267002 0 267058 800
rect 267646 0 267702 800
rect 268382 0 268438 800
rect 269118 0 269174 800
rect 269854 0 269910 800
rect 270590 0 270646 800
rect 271234 0 271290 800
rect 271970 0 272026 800
rect 272706 0 272762 800
rect 273442 0 273498 800
rect 274086 0 274142 800
rect 274822 0 274878 800
rect 275558 0 275614 800
rect 276294 0 276350 800
rect 277030 0 277086 800
rect 277674 0 277730 800
rect 278410 0 278466 800
rect 279146 0 279202 800
rect 279882 0 279938 800
rect 280618 0 280674 800
rect 281262 0 281318 800
rect 281998 0 282054 800
rect 282734 0 282790 800
rect 283470 0 283526 800
rect 284206 0 284262 800
rect 284850 0 284906 800
rect 285586 0 285642 800
rect 286322 0 286378 800
rect 287058 0 287114 800
rect 287794 0 287850 800
rect 288438 0 288494 800
rect 289174 0 289230 800
rect 289910 0 289966 800
rect 290646 0 290702 800
rect 291382 0 291438 800
rect 292026 0 292082 800
rect 292762 0 292818 800
rect 293498 0 293554 800
rect 294234 0 294290 800
rect 294878 0 294934 800
rect 295614 0 295670 800
rect 296350 0 296406 800
rect 297086 0 297142 800
rect 297822 0 297878 800
rect 298466 0 298522 800
rect 299202 0 299258 800
rect 299938 0 299994 800
rect 300674 0 300730 800
rect 301410 0 301466 800
rect 302054 0 302110 800
rect 302790 0 302846 800
rect 303526 0 303582 800
rect 304262 0 304318 800
rect 304998 0 305054 800
rect 305642 0 305698 800
rect 306378 0 306434 800
rect 307114 0 307170 800
rect 307850 0 307906 800
rect 308586 0 308642 800
rect 309230 0 309286 800
rect 309966 0 310022 800
rect 310702 0 310758 800
rect 311438 0 311494 800
rect 312174 0 312230 800
rect 312818 0 312874 800
rect 313554 0 313610 800
rect 314290 0 314346 800
rect 315026 0 315082 800
rect 315670 0 315726 800
rect 316406 0 316462 800
rect 317142 0 317198 800
rect 317878 0 317934 800
rect 318614 0 318670 800
rect 319258 0 319314 800
rect 319994 0 320050 800
rect 320730 0 320786 800
rect 321466 0 321522 800
rect 322202 0 322258 800
rect 322846 0 322902 800
rect 323582 0 323638 800
rect 324318 0 324374 800
rect 325054 0 325110 800
rect 325790 0 325846 800
rect 326434 0 326490 800
rect 327170 0 327226 800
rect 327906 0 327962 800
rect 328642 0 328698 800
rect 329378 0 329434 800
rect 330022 0 330078 800
rect 330758 0 330814 800
rect 331494 0 331550 800
rect 332230 0 332286 800
rect 332966 0 333022 800
rect 333610 0 333666 800
rect 334346 0 334402 800
rect 335082 0 335138 800
rect 335818 0 335874 800
rect 336462 0 336518 800
rect 337198 0 337254 800
rect 337934 0 337990 800
rect 338670 0 338726 800
rect 339406 0 339462 800
rect 340050 0 340106 800
rect 340786 0 340842 800
rect 341522 0 341578 800
rect 342258 0 342314 800
rect 342994 0 343050 800
rect 343638 0 343694 800
rect 344374 0 344430 800
rect 345110 0 345166 800
rect 345846 0 345902 800
rect 346582 0 346638 800
rect 347226 0 347282 800
rect 347962 0 348018 800
rect 348698 0 348754 800
rect 349434 0 349490 800
rect 350170 0 350226 800
rect 350814 0 350870 800
rect 351550 0 351606 800
rect 352286 0 352342 800
rect 353022 0 353078 800
<< obsm2 >>
rect 204 354767 1434 354906
rect 1602 354767 4470 354906
rect 4638 354767 7598 354906
rect 7766 354767 10726 354906
rect 10894 354767 13762 354906
rect 13930 354767 16890 354906
rect 17058 354767 20018 354906
rect 20186 354767 23054 354906
rect 23222 354767 26182 354906
rect 26350 354767 29310 354906
rect 29478 354767 32438 354906
rect 32606 354767 35474 354906
rect 35642 354767 38602 354906
rect 38770 354767 41730 354906
rect 41898 354767 44766 354906
rect 44934 354767 47894 354906
rect 48062 354767 51022 354906
rect 51190 354767 54058 354906
rect 54226 354767 57186 354906
rect 57354 354767 60314 354906
rect 60482 354767 63442 354906
rect 63610 354767 66478 354906
rect 66646 354767 69606 354906
rect 69774 354767 72734 354906
rect 72902 354767 75770 354906
rect 75938 354767 78898 354906
rect 79066 354767 82026 354906
rect 82194 354767 85062 354906
rect 85230 354767 88190 354906
rect 88358 354767 91318 354906
rect 91486 354767 94446 354906
rect 94614 354767 97482 354906
rect 97650 354767 100610 354906
rect 100778 354767 103738 354906
rect 103906 354767 106774 354906
rect 106942 354767 109902 354906
rect 110070 354767 113030 354906
rect 113198 354767 116066 354906
rect 116234 354767 119194 354906
rect 119362 354767 122322 354906
rect 122490 354767 125450 354906
rect 125618 354767 128486 354906
rect 128654 354767 131614 354906
rect 131782 354767 134742 354906
rect 134910 354767 137778 354906
rect 137946 354767 140906 354906
rect 141074 354767 144034 354906
rect 144202 354767 147070 354906
rect 147238 354767 150198 354906
rect 150366 354767 153326 354906
rect 153494 354767 156454 354906
rect 156622 354767 159490 354906
rect 159658 354767 162618 354906
rect 162786 354767 165746 354906
rect 165914 354767 168782 354906
rect 168950 354767 171910 354906
rect 172078 354767 175038 354906
rect 175206 354767 178166 354906
rect 178334 354767 181202 354906
rect 181370 354767 184330 354906
rect 184498 354767 187458 354906
rect 187626 354767 190494 354906
rect 190662 354767 193622 354906
rect 193790 354767 196750 354906
rect 196918 354767 199786 354906
rect 199954 354767 202914 354906
rect 203082 354767 206042 354906
rect 206210 354767 209170 354906
rect 209338 354767 212206 354906
rect 212374 354767 215334 354906
rect 215502 354767 218462 354906
rect 218630 354767 221498 354906
rect 221666 354767 224626 354906
rect 224794 354767 227754 354906
rect 227922 354767 230790 354906
rect 230958 354767 233918 354906
rect 234086 354767 237046 354906
rect 237214 354767 240174 354906
rect 240342 354767 243210 354906
rect 243378 354767 246338 354906
rect 246506 354767 249466 354906
rect 249634 354767 252502 354906
rect 252670 354767 255630 354906
rect 255798 354767 258758 354906
rect 258926 354767 261794 354906
rect 261962 354767 264922 354906
rect 265090 354767 268050 354906
rect 268218 354767 271178 354906
rect 271346 354767 274214 354906
rect 274382 354767 277342 354906
rect 277510 354767 280470 354906
rect 280638 354767 283506 354906
rect 283674 354767 286634 354906
rect 286802 354767 289762 354906
rect 289930 354767 292798 354906
rect 292966 354767 295926 354906
rect 296094 354767 299054 354906
rect 299222 354767 302182 354906
rect 302350 354767 305218 354906
rect 305386 354767 308346 354906
rect 308514 354767 311474 354906
rect 311642 354767 314510 354906
rect 314678 354767 317638 354906
rect 317806 354767 320766 354906
rect 320934 354767 323802 354906
rect 323970 354767 326930 354906
rect 327098 354767 330058 354906
rect 330226 354767 333186 354906
rect 333354 354767 336222 354906
rect 336390 354767 339350 354906
rect 339518 354767 342478 354906
rect 342646 354767 345514 354906
rect 345682 354767 348642 354906
rect 348810 354767 351770 354906
rect 351938 354767 353446 354906
rect 204 856 353446 354767
rect 204 2 238 856
rect 406 2 882 856
rect 1050 2 1618 856
rect 1786 2 2354 856
rect 2522 2 3090 856
rect 3258 2 3734 856
rect 3902 2 4470 856
rect 4638 2 5206 856
rect 5374 2 5942 856
rect 6110 2 6678 856
rect 6846 2 7322 856
rect 7490 2 8058 856
rect 8226 2 8794 856
rect 8962 2 9530 856
rect 9698 2 10266 856
rect 10434 2 10910 856
rect 11078 2 11646 856
rect 11814 2 12382 856
rect 12550 2 13118 856
rect 13286 2 13854 856
rect 14022 2 14498 856
rect 14666 2 15234 856
rect 15402 2 15970 856
rect 16138 2 16706 856
rect 16874 2 17442 856
rect 17610 2 18086 856
rect 18254 2 18822 856
rect 18990 2 19558 856
rect 19726 2 20294 856
rect 20462 2 21030 856
rect 21198 2 21674 856
rect 21842 2 22410 856
rect 22578 2 23146 856
rect 23314 2 23882 856
rect 24050 2 24526 856
rect 24694 2 25262 856
rect 25430 2 25998 856
rect 26166 2 26734 856
rect 26902 2 27470 856
rect 27638 2 28114 856
rect 28282 2 28850 856
rect 29018 2 29586 856
rect 29754 2 30322 856
rect 30490 2 31058 856
rect 31226 2 31702 856
rect 31870 2 32438 856
rect 32606 2 33174 856
rect 33342 2 33910 856
rect 34078 2 34646 856
rect 34814 2 35290 856
rect 35458 2 36026 856
rect 36194 2 36762 856
rect 36930 2 37498 856
rect 37666 2 38234 856
rect 38402 2 38878 856
rect 39046 2 39614 856
rect 39782 2 40350 856
rect 40518 2 41086 856
rect 41254 2 41822 856
rect 41990 2 42466 856
rect 42634 2 43202 856
rect 43370 2 43938 856
rect 44106 2 44674 856
rect 44842 2 45318 856
rect 45486 2 46054 856
rect 46222 2 46790 856
rect 46958 2 47526 856
rect 47694 2 48262 856
rect 48430 2 48906 856
rect 49074 2 49642 856
rect 49810 2 50378 856
rect 50546 2 51114 856
rect 51282 2 51850 856
rect 52018 2 52494 856
rect 52662 2 53230 856
rect 53398 2 53966 856
rect 54134 2 54702 856
rect 54870 2 55438 856
rect 55606 2 56082 856
rect 56250 2 56818 856
rect 56986 2 57554 856
rect 57722 2 58290 856
rect 58458 2 59026 856
rect 59194 2 59670 856
rect 59838 2 60406 856
rect 60574 2 61142 856
rect 61310 2 61878 856
rect 62046 2 62614 856
rect 62782 2 63258 856
rect 63426 2 63994 856
rect 64162 2 64730 856
rect 64898 2 65466 856
rect 65634 2 66110 856
rect 66278 2 66846 856
rect 67014 2 67582 856
rect 67750 2 68318 856
rect 68486 2 69054 856
rect 69222 2 69698 856
rect 69866 2 70434 856
rect 70602 2 71170 856
rect 71338 2 71906 856
rect 72074 2 72642 856
rect 72810 2 73286 856
rect 73454 2 74022 856
rect 74190 2 74758 856
rect 74926 2 75494 856
rect 75662 2 76230 856
rect 76398 2 76874 856
rect 77042 2 77610 856
rect 77778 2 78346 856
rect 78514 2 79082 856
rect 79250 2 79818 856
rect 79986 2 80462 856
rect 80630 2 81198 856
rect 81366 2 81934 856
rect 82102 2 82670 856
rect 82838 2 83406 856
rect 83574 2 84050 856
rect 84218 2 84786 856
rect 84954 2 85522 856
rect 85690 2 86258 856
rect 86426 2 86902 856
rect 87070 2 87638 856
rect 87806 2 88374 856
rect 88542 2 89110 856
rect 89278 2 89846 856
rect 90014 2 90490 856
rect 90658 2 91226 856
rect 91394 2 91962 856
rect 92130 2 92698 856
rect 92866 2 93434 856
rect 93602 2 94078 856
rect 94246 2 94814 856
rect 94982 2 95550 856
rect 95718 2 96286 856
rect 96454 2 97022 856
rect 97190 2 97666 856
rect 97834 2 98402 856
rect 98570 2 99138 856
rect 99306 2 99874 856
rect 100042 2 100610 856
rect 100778 2 101254 856
rect 101422 2 101990 856
rect 102158 2 102726 856
rect 102894 2 103462 856
rect 103630 2 104198 856
rect 104366 2 104842 856
rect 105010 2 105578 856
rect 105746 2 106314 856
rect 106482 2 107050 856
rect 107218 2 107694 856
rect 107862 2 108430 856
rect 108598 2 109166 856
rect 109334 2 109902 856
rect 110070 2 110638 856
rect 110806 2 111282 856
rect 111450 2 112018 856
rect 112186 2 112754 856
rect 112922 2 113490 856
rect 113658 2 114226 856
rect 114394 2 114870 856
rect 115038 2 115606 856
rect 115774 2 116342 856
rect 116510 2 117078 856
rect 117246 2 117814 856
rect 117982 2 118458 856
rect 118626 2 119194 856
rect 119362 2 119930 856
rect 120098 2 120666 856
rect 120834 2 121402 856
rect 121570 2 122046 856
rect 122214 2 122782 856
rect 122950 2 123518 856
rect 123686 2 124254 856
rect 124422 2 124990 856
rect 125158 2 125634 856
rect 125802 2 126370 856
rect 126538 2 127106 856
rect 127274 2 127842 856
rect 128010 2 128486 856
rect 128654 2 129222 856
rect 129390 2 129958 856
rect 130126 2 130694 856
rect 130862 2 131430 856
rect 131598 2 132074 856
rect 132242 2 132810 856
rect 132978 2 133546 856
rect 133714 2 134282 856
rect 134450 2 135018 856
rect 135186 2 135662 856
rect 135830 2 136398 856
rect 136566 2 137134 856
rect 137302 2 137870 856
rect 138038 2 138606 856
rect 138774 2 139250 856
rect 139418 2 139986 856
rect 140154 2 140722 856
rect 140890 2 141458 856
rect 141626 2 142194 856
rect 142362 2 142838 856
rect 143006 2 143574 856
rect 143742 2 144310 856
rect 144478 2 145046 856
rect 145214 2 145782 856
rect 145950 2 146426 856
rect 146594 2 147162 856
rect 147330 2 147898 856
rect 148066 2 148634 856
rect 148802 2 149278 856
rect 149446 2 150014 856
rect 150182 2 150750 856
rect 150918 2 151486 856
rect 151654 2 152222 856
rect 152390 2 152866 856
rect 153034 2 153602 856
rect 153770 2 154338 856
rect 154506 2 155074 856
rect 155242 2 155810 856
rect 155978 2 156454 856
rect 156622 2 157190 856
rect 157358 2 157926 856
rect 158094 2 158662 856
rect 158830 2 159398 856
rect 159566 2 160042 856
rect 160210 2 160778 856
rect 160946 2 161514 856
rect 161682 2 162250 856
rect 162418 2 162986 856
rect 163154 2 163630 856
rect 163798 2 164366 856
rect 164534 2 165102 856
rect 165270 2 165838 856
rect 166006 2 166574 856
rect 166742 2 167218 856
rect 167386 2 167954 856
rect 168122 2 168690 856
rect 168858 2 169426 856
rect 169594 2 170070 856
rect 170238 2 170806 856
rect 170974 2 171542 856
rect 171710 2 172278 856
rect 172446 2 173014 856
rect 173182 2 173658 856
rect 173826 2 174394 856
rect 174562 2 175130 856
rect 175298 2 175866 856
rect 176034 2 176602 856
rect 176770 2 177246 856
rect 177414 2 177982 856
rect 178150 2 178718 856
rect 178886 2 179454 856
rect 179622 2 180190 856
rect 180358 2 180834 856
rect 181002 2 181570 856
rect 181738 2 182306 856
rect 182474 2 183042 856
rect 183210 2 183778 856
rect 183946 2 184422 856
rect 184590 2 185158 856
rect 185326 2 185894 856
rect 186062 2 186630 856
rect 186798 2 187366 856
rect 187534 2 188010 856
rect 188178 2 188746 856
rect 188914 2 189482 856
rect 189650 2 190218 856
rect 190386 2 190862 856
rect 191030 2 191598 856
rect 191766 2 192334 856
rect 192502 2 193070 856
rect 193238 2 193806 856
rect 193974 2 194450 856
rect 194618 2 195186 856
rect 195354 2 195922 856
rect 196090 2 196658 856
rect 196826 2 197394 856
rect 197562 2 198038 856
rect 198206 2 198774 856
rect 198942 2 199510 856
rect 199678 2 200246 856
rect 200414 2 200982 856
rect 201150 2 201626 856
rect 201794 2 202362 856
rect 202530 2 203098 856
rect 203266 2 203834 856
rect 204002 2 204570 856
rect 204738 2 205214 856
rect 205382 2 205950 856
rect 206118 2 206686 856
rect 206854 2 207422 856
rect 207590 2 208158 856
rect 208326 2 208802 856
rect 208970 2 209538 856
rect 209706 2 210274 856
rect 210442 2 211010 856
rect 211178 2 211654 856
rect 211822 2 212390 856
rect 212558 2 213126 856
rect 213294 2 213862 856
rect 214030 2 214598 856
rect 214766 2 215242 856
rect 215410 2 215978 856
rect 216146 2 216714 856
rect 216882 2 217450 856
rect 217618 2 218186 856
rect 218354 2 218830 856
rect 218998 2 219566 856
rect 219734 2 220302 856
rect 220470 2 221038 856
rect 221206 2 221774 856
rect 221942 2 222418 856
rect 222586 2 223154 856
rect 223322 2 223890 856
rect 224058 2 224626 856
rect 224794 2 225362 856
rect 225530 2 226006 856
rect 226174 2 226742 856
rect 226910 2 227478 856
rect 227646 2 228214 856
rect 228382 2 228950 856
rect 229118 2 229594 856
rect 229762 2 230330 856
rect 230498 2 231066 856
rect 231234 2 231802 856
rect 231970 2 232446 856
rect 232614 2 233182 856
rect 233350 2 233918 856
rect 234086 2 234654 856
rect 234822 2 235390 856
rect 235558 2 236034 856
rect 236202 2 236770 856
rect 236938 2 237506 856
rect 237674 2 238242 856
rect 238410 2 238978 856
rect 239146 2 239622 856
rect 239790 2 240358 856
rect 240526 2 241094 856
rect 241262 2 241830 856
rect 241998 2 242566 856
rect 242734 2 243210 856
rect 243378 2 243946 856
rect 244114 2 244682 856
rect 244850 2 245418 856
rect 245586 2 246154 856
rect 246322 2 246798 856
rect 246966 2 247534 856
rect 247702 2 248270 856
rect 248438 2 249006 856
rect 249174 2 249742 856
rect 249910 2 250386 856
rect 250554 2 251122 856
rect 251290 2 251858 856
rect 252026 2 252594 856
rect 252762 2 253238 856
rect 253406 2 253974 856
rect 254142 2 254710 856
rect 254878 2 255446 856
rect 255614 2 256182 856
rect 256350 2 256826 856
rect 256994 2 257562 856
rect 257730 2 258298 856
rect 258466 2 259034 856
rect 259202 2 259770 856
rect 259938 2 260414 856
rect 260582 2 261150 856
rect 261318 2 261886 856
rect 262054 2 262622 856
rect 262790 2 263358 856
rect 263526 2 264002 856
rect 264170 2 264738 856
rect 264906 2 265474 856
rect 265642 2 266210 856
rect 266378 2 266946 856
rect 267114 2 267590 856
rect 267758 2 268326 856
rect 268494 2 269062 856
rect 269230 2 269798 856
rect 269966 2 270534 856
rect 270702 2 271178 856
rect 271346 2 271914 856
rect 272082 2 272650 856
rect 272818 2 273386 856
rect 273554 2 274030 856
rect 274198 2 274766 856
rect 274934 2 275502 856
rect 275670 2 276238 856
rect 276406 2 276974 856
rect 277142 2 277618 856
rect 277786 2 278354 856
rect 278522 2 279090 856
rect 279258 2 279826 856
rect 279994 2 280562 856
rect 280730 2 281206 856
rect 281374 2 281942 856
rect 282110 2 282678 856
rect 282846 2 283414 856
rect 283582 2 284150 856
rect 284318 2 284794 856
rect 284962 2 285530 856
rect 285698 2 286266 856
rect 286434 2 287002 856
rect 287170 2 287738 856
rect 287906 2 288382 856
rect 288550 2 289118 856
rect 289286 2 289854 856
rect 290022 2 290590 856
rect 290758 2 291326 856
rect 291494 2 291970 856
rect 292138 2 292706 856
rect 292874 2 293442 856
rect 293610 2 294178 856
rect 294346 2 294822 856
rect 294990 2 295558 856
rect 295726 2 296294 856
rect 296462 2 297030 856
rect 297198 2 297766 856
rect 297934 2 298410 856
rect 298578 2 299146 856
rect 299314 2 299882 856
rect 300050 2 300618 856
rect 300786 2 301354 856
rect 301522 2 301998 856
rect 302166 2 302734 856
rect 302902 2 303470 856
rect 303638 2 304206 856
rect 304374 2 304942 856
rect 305110 2 305586 856
rect 305754 2 306322 856
rect 306490 2 307058 856
rect 307226 2 307794 856
rect 307962 2 308530 856
rect 308698 2 309174 856
rect 309342 2 309910 856
rect 310078 2 310646 856
rect 310814 2 311382 856
rect 311550 2 312118 856
rect 312286 2 312762 856
rect 312930 2 313498 856
rect 313666 2 314234 856
rect 314402 2 314970 856
rect 315138 2 315614 856
rect 315782 2 316350 856
rect 316518 2 317086 856
rect 317254 2 317822 856
rect 317990 2 318558 856
rect 318726 2 319202 856
rect 319370 2 319938 856
rect 320106 2 320674 856
rect 320842 2 321410 856
rect 321578 2 322146 856
rect 322314 2 322790 856
rect 322958 2 323526 856
rect 323694 2 324262 856
rect 324430 2 324998 856
rect 325166 2 325734 856
rect 325902 2 326378 856
rect 326546 2 327114 856
rect 327282 2 327850 856
rect 328018 2 328586 856
rect 328754 2 329322 856
rect 329490 2 329966 856
rect 330134 2 330702 856
rect 330870 2 331438 856
rect 331606 2 332174 856
rect 332342 2 332910 856
rect 333078 2 333554 856
rect 333722 2 334290 856
rect 334458 2 335026 856
rect 335194 2 335762 856
rect 335930 2 336406 856
rect 336574 2 337142 856
rect 337310 2 337878 856
rect 338046 2 338614 856
rect 338782 2 339350 856
rect 339518 2 339994 856
rect 340162 2 340730 856
rect 340898 2 341466 856
rect 341634 2 342202 856
rect 342370 2 342938 856
rect 343106 2 343582 856
rect 343750 2 344318 856
rect 344486 2 345054 856
rect 345222 2 345790 856
rect 345958 2 346526 856
rect 346694 2 347170 856
rect 347338 2 347906 856
rect 348074 2 348642 856
rect 348810 2 349378 856
rect 349546 2 350114 856
rect 350282 2 350758 856
rect 350926 2 351494 856
rect 351662 2 352230 856
rect 352398 2 352966 856
rect 353134 2 353446 856
<< metal3 >>
rect 0 355104 800 355224
rect 0 354424 800 354544
rect 352679 354560 353479 354680
rect 0 353744 800 353864
rect 0 353064 800 353184
rect 352679 352792 353479 352912
rect 0 352384 800 352504
rect 0 351568 800 351688
rect 0 350888 800 351008
rect 352679 351024 353479 351144
rect 0 350208 800 350328
rect 0 349528 800 349648
rect 352679 349256 353479 349376
rect 0 348848 800 348968
rect 0 348168 800 348288
rect 0 347352 800 347472
rect 352679 347488 353479 347608
rect 0 346672 800 346792
rect 0 345992 800 346112
rect 352679 345720 353479 345840
rect 0 345312 800 345432
rect 0 344632 800 344752
rect 0 343816 800 343936
rect 352679 343952 353479 344072
rect 0 343136 800 343256
rect 0 342456 800 342576
rect 352679 342184 353479 342304
rect 0 341776 800 341896
rect 0 341096 800 341216
rect 0 340416 800 340536
rect 352679 340416 353479 340536
rect 0 339600 800 339720
rect 0 338920 800 339040
rect 352679 338648 353479 338768
rect 0 338240 800 338360
rect 0 337560 800 337680
rect 0 336880 800 337000
rect 352679 336880 353479 337000
rect 0 336200 800 336320
rect 0 335384 800 335504
rect 352679 335112 353479 335232
rect 0 334704 800 334824
rect 0 334024 800 334144
rect 0 333344 800 333464
rect 352679 333344 353479 333464
rect 0 332664 800 332784
rect 0 331848 800 331968
rect 352679 331440 353479 331560
rect 0 331168 800 331288
rect 0 330488 800 330608
rect 0 329808 800 329928
rect 352679 329672 353479 329792
rect 0 329128 800 329248
rect 0 328448 800 328568
rect 352679 327904 353479 328024
rect 0 327632 800 327752
rect 0 326952 800 327072
rect 0 326272 800 326392
rect 352679 326136 353479 326256
rect 0 325592 800 325712
rect 0 324912 800 325032
rect 352679 324368 353479 324488
rect 0 324096 800 324216
rect 0 323416 800 323536
rect 0 322736 800 322856
rect 352679 322600 353479 322720
rect 0 322056 800 322176
rect 0 321376 800 321496
rect 0 320696 800 320816
rect 352679 320832 353479 320952
rect 0 319880 800 320000
rect 0 319200 800 319320
rect 352679 319064 353479 319184
rect 0 318520 800 318640
rect 0 317840 800 317960
rect 0 317160 800 317280
rect 352679 317296 353479 317416
rect 0 316480 800 316600
rect 0 315664 800 315784
rect 352679 315528 353479 315648
rect 0 314984 800 315104
rect 0 314304 800 314424
rect 0 313624 800 313744
rect 352679 313760 353479 313880
rect 0 312944 800 313064
rect 0 312128 800 312248
rect 352679 311992 353479 312112
rect 0 311448 800 311568
rect 0 310768 800 310888
rect 0 310088 800 310208
rect 352679 310224 353479 310344
rect 0 309408 800 309528
rect 0 308728 800 308848
rect 352679 308320 353479 308440
rect 0 307912 800 308032
rect 0 307232 800 307352
rect 0 306552 800 306672
rect 352679 306552 353479 306672
rect 0 305872 800 305992
rect 0 305192 800 305312
rect 352679 304784 353479 304904
rect 0 304376 800 304496
rect 0 303696 800 303816
rect 0 303016 800 303136
rect 352679 303016 353479 303136
rect 0 302336 800 302456
rect 0 301656 800 301776
rect 352679 301248 353479 301368
rect 0 300976 800 301096
rect 0 300160 800 300280
rect 0 299480 800 299600
rect 352679 299480 353479 299600
rect 0 298800 800 298920
rect 0 298120 800 298240
rect 352679 297712 353479 297832
rect 0 297440 800 297560
rect 0 296760 800 296880
rect 0 295944 800 296064
rect 352679 295944 353479 296064
rect 0 295264 800 295384
rect 0 294584 800 294704
rect 352679 294176 353479 294296
rect 0 293904 800 294024
rect 0 293224 800 293344
rect 0 292408 800 292528
rect 352679 292408 353479 292528
rect 0 291728 800 291848
rect 0 291048 800 291168
rect 352679 290640 353479 290760
rect 0 290368 800 290488
rect 0 289688 800 289808
rect 0 289008 800 289128
rect 352679 288872 353479 288992
rect 0 288192 800 288312
rect 0 287512 800 287632
rect 352679 287104 353479 287224
rect 0 286832 800 286952
rect 0 286152 800 286272
rect 0 285472 800 285592
rect 352679 285336 353479 285456
rect 0 284792 800 284912
rect 0 283976 800 284096
rect 0 283296 800 283416
rect 352679 283432 353479 283552
rect 0 282616 800 282736
rect 0 281936 800 282056
rect 352679 281664 353479 281784
rect 0 281256 800 281376
rect 0 280440 800 280560
rect 0 279760 800 279880
rect 352679 279896 353479 280016
rect 0 279080 800 279200
rect 0 278400 800 278520
rect 352679 278128 353479 278248
rect 0 277720 800 277840
rect 0 277040 800 277160
rect 0 276224 800 276344
rect 352679 276360 353479 276480
rect 0 275544 800 275664
rect 0 274864 800 274984
rect 352679 274592 353479 274712
rect 0 274184 800 274304
rect 0 273504 800 273624
rect 0 272688 800 272808
rect 352679 272824 353479 272944
rect 0 272008 800 272128
rect 0 271328 800 271448
rect 352679 271056 353479 271176
rect 0 270648 800 270768
rect 0 269968 800 270088
rect 0 269288 800 269408
rect 352679 269288 353479 269408
rect 0 268472 800 268592
rect 0 267792 800 267912
rect 352679 267520 353479 267640
rect 0 267112 800 267232
rect 0 266432 800 266552
rect 0 265752 800 265872
rect 352679 265752 353479 265872
rect 0 265072 800 265192
rect 0 264256 800 264376
rect 352679 263984 353479 264104
rect 0 263576 800 263696
rect 0 262896 800 263016
rect 0 262216 800 262336
rect 352679 262216 353479 262336
rect 0 261536 800 261656
rect 0 260720 800 260840
rect 352679 260312 353479 260432
rect 0 260040 800 260160
rect 0 259360 800 259480
rect 0 258680 800 258800
rect 352679 258544 353479 258664
rect 0 258000 800 258120
rect 0 257320 800 257440
rect 352679 256776 353479 256896
rect 0 256504 800 256624
rect 0 255824 800 255944
rect 0 255144 800 255264
rect 352679 255008 353479 255128
rect 0 254464 800 254584
rect 0 253784 800 253904
rect 352679 253240 353479 253360
rect 0 252968 800 253088
rect 0 252288 800 252408
rect 0 251608 800 251728
rect 352679 251472 353479 251592
rect 0 250928 800 251048
rect 0 250248 800 250368
rect 0 249568 800 249688
rect 352679 249704 353479 249824
rect 0 248752 800 248872
rect 0 248072 800 248192
rect 352679 247936 353479 248056
rect 0 247392 800 247512
rect 0 246712 800 246832
rect 0 246032 800 246152
rect 352679 246168 353479 246288
rect 0 245352 800 245472
rect 0 244536 800 244656
rect 352679 244400 353479 244520
rect 0 243856 800 243976
rect 0 243176 800 243296
rect 0 242496 800 242616
rect 352679 242632 353479 242752
rect 0 241816 800 241936
rect 0 241000 800 241120
rect 352679 240864 353479 240984
rect 0 240320 800 240440
rect 0 239640 800 239760
rect 0 238960 800 239080
rect 352679 239096 353479 239216
rect 0 238280 800 238400
rect 0 237600 800 237720
rect 352679 237192 353479 237312
rect 0 236784 800 236904
rect 0 236104 800 236224
rect 0 235424 800 235544
rect 352679 235424 353479 235544
rect 0 234744 800 234864
rect 0 234064 800 234184
rect 352679 233656 353479 233776
rect 0 233248 800 233368
rect 0 232568 800 232688
rect 0 231888 800 232008
rect 352679 231888 353479 232008
rect 0 231208 800 231328
rect 0 230528 800 230648
rect 352679 230120 353479 230240
rect 0 229848 800 229968
rect 0 229032 800 229152
rect 0 228352 800 228472
rect 352679 228352 353479 228472
rect 0 227672 800 227792
rect 0 226992 800 227112
rect 352679 226584 353479 226704
rect 0 226312 800 226432
rect 0 225632 800 225752
rect 0 224816 800 224936
rect 352679 224816 353479 224936
rect 0 224136 800 224256
rect 0 223456 800 223576
rect 352679 223048 353479 223168
rect 0 222776 800 222896
rect 0 222096 800 222216
rect 0 221280 800 221400
rect 352679 221280 353479 221400
rect 0 220600 800 220720
rect 0 219920 800 220040
rect 352679 219512 353479 219632
rect 0 219240 800 219360
rect 0 218560 800 218680
rect 0 217880 800 218000
rect 352679 217744 353479 217864
rect 0 217064 800 217184
rect 0 216384 800 216504
rect 352679 215976 353479 216096
rect 0 215704 800 215824
rect 0 215024 800 215144
rect 0 214344 800 214464
rect 352679 214208 353479 214328
rect 0 213664 800 213784
rect 0 212848 800 212968
rect 0 212168 800 212288
rect 352679 212304 353479 212424
rect 0 211488 800 211608
rect 0 210808 800 210928
rect 352679 210536 353479 210656
rect 0 210128 800 210248
rect 0 209312 800 209432
rect 0 208632 800 208752
rect 352679 208768 353479 208888
rect 0 207952 800 208072
rect 0 207272 800 207392
rect 352679 207000 353479 207120
rect 0 206592 800 206712
rect 0 205912 800 206032
rect 0 205096 800 205216
rect 352679 205232 353479 205352
rect 0 204416 800 204536
rect 0 203736 800 203856
rect 352679 203464 353479 203584
rect 0 203056 800 203176
rect 0 202376 800 202496
rect 0 201560 800 201680
rect 352679 201696 353479 201816
rect 0 200880 800 201000
rect 0 200200 800 200320
rect 352679 199928 353479 200048
rect 0 199520 800 199640
rect 0 198840 800 198960
rect 0 198160 800 198280
rect 352679 198160 353479 198280
rect 0 197344 800 197464
rect 0 196664 800 196784
rect 352679 196392 353479 196512
rect 0 195984 800 196104
rect 0 195304 800 195424
rect 0 194624 800 194744
rect 352679 194624 353479 194744
rect 0 193944 800 194064
rect 0 193128 800 193248
rect 352679 192856 353479 192976
rect 0 192448 800 192568
rect 0 191768 800 191888
rect 0 191088 800 191208
rect 352679 191088 353479 191208
rect 0 190408 800 190528
rect 0 189592 800 189712
rect 352679 189184 353479 189304
rect 0 188912 800 189032
rect 0 188232 800 188352
rect 0 187552 800 187672
rect 352679 187416 353479 187536
rect 0 186872 800 186992
rect 0 186192 800 186312
rect 352679 185648 353479 185768
rect 0 185376 800 185496
rect 0 184696 800 184816
rect 0 184016 800 184136
rect 352679 183880 353479 184000
rect 0 183336 800 183456
rect 0 182656 800 182776
rect 352679 182112 353479 182232
rect 0 181840 800 181960
rect 0 181160 800 181280
rect 0 180480 800 180600
rect 352679 180344 353479 180464
rect 0 179800 800 179920
rect 0 179120 800 179240
rect 0 178440 800 178560
rect 352679 178576 353479 178696
rect 0 177624 800 177744
rect 0 176944 800 177064
rect 352679 176808 353479 176928
rect 0 176264 800 176384
rect 0 175584 800 175704
rect 0 174904 800 175024
rect 352679 175040 353479 175160
rect 0 174224 800 174344
rect 0 173408 800 173528
rect 352679 173272 353479 173392
rect 0 172728 800 172848
rect 0 172048 800 172168
rect 0 171368 800 171488
rect 352679 171504 353479 171624
rect 0 170688 800 170808
rect 0 169872 800 169992
rect 352679 169736 353479 169856
rect 0 169192 800 169312
rect 0 168512 800 168632
rect 0 167832 800 167952
rect 352679 167968 353479 168088
rect 0 167152 800 167272
rect 0 166472 800 166592
rect 352679 166064 353479 166184
rect 0 165656 800 165776
rect 0 164976 800 165096
rect 0 164296 800 164416
rect 352679 164296 353479 164416
rect 0 163616 800 163736
rect 0 162936 800 163056
rect 352679 162528 353479 162648
rect 0 162120 800 162240
rect 0 161440 800 161560
rect 0 160760 800 160880
rect 352679 160760 353479 160880
rect 0 160080 800 160200
rect 0 159400 800 159520
rect 352679 158992 353479 159112
rect 0 158720 800 158840
rect 0 157904 800 158024
rect 0 157224 800 157344
rect 352679 157224 353479 157344
rect 0 156544 800 156664
rect 0 155864 800 155984
rect 352679 155456 353479 155576
rect 0 155184 800 155304
rect 0 154504 800 154624
rect 0 153688 800 153808
rect 352679 153688 353479 153808
rect 0 153008 800 153128
rect 0 152328 800 152448
rect 352679 151920 353479 152040
rect 0 151648 800 151768
rect 0 150968 800 151088
rect 0 150152 800 150272
rect 352679 150152 353479 150272
rect 0 149472 800 149592
rect 0 148792 800 148912
rect 352679 148384 353479 148504
rect 0 148112 800 148232
rect 0 147432 800 147552
rect 0 146752 800 146872
rect 352679 146616 353479 146736
rect 0 145936 800 146056
rect 0 145256 800 145376
rect 352679 144848 353479 144968
rect 0 144576 800 144696
rect 0 143896 800 144016
rect 0 143216 800 143336
rect 352679 143080 353479 143200
rect 0 142536 800 142656
rect 0 141720 800 141840
rect 0 141040 800 141160
rect 352679 141176 353479 141296
rect 0 140360 800 140480
rect 0 139680 800 139800
rect 352679 139408 353479 139528
rect 0 139000 800 139120
rect 0 138184 800 138304
rect 0 137504 800 137624
rect 352679 137640 353479 137760
rect 0 136824 800 136944
rect 0 136144 800 136264
rect 352679 135872 353479 135992
rect 0 135464 800 135584
rect 0 134784 800 134904
rect 0 133968 800 134088
rect 352679 134104 353479 134224
rect 0 133288 800 133408
rect 0 132608 800 132728
rect 352679 132336 353479 132456
rect 0 131928 800 132048
rect 0 131248 800 131368
rect 0 130432 800 130552
rect 352679 130568 353479 130688
rect 0 129752 800 129872
rect 0 129072 800 129192
rect 352679 128800 353479 128920
rect 0 128392 800 128512
rect 0 127712 800 127832
rect 0 127032 800 127152
rect 352679 127032 353479 127152
rect 0 126216 800 126336
rect 0 125536 800 125656
rect 352679 125264 353479 125384
rect 0 124856 800 124976
rect 0 124176 800 124296
rect 0 123496 800 123616
rect 352679 123496 353479 123616
rect 0 122816 800 122936
rect 0 122000 800 122120
rect 352679 121728 353479 121848
rect 0 121320 800 121440
rect 0 120640 800 120760
rect 0 119960 800 120080
rect 352679 119960 353479 120080
rect 0 119280 800 119400
rect 0 118464 800 118584
rect 352679 118056 353479 118176
rect 0 117784 800 117904
rect 0 117104 800 117224
rect 0 116424 800 116544
rect 352679 116288 353479 116408
rect 0 115744 800 115864
rect 0 115064 800 115184
rect 352679 114520 353479 114640
rect 0 114248 800 114368
rect 0 113568 800 113688
rect 0 112888 800 113008
rect 352679 112752 353479 112872
rect 0 112208 800 112328
rect 0 111528 800 111648
rect 352679 110984 353479 111104
rect 0 110712 800 110832
rect 0 110032 800 110152
rect 0 109352 800 109472
rect 352679 109216 353479 109336
rect 0 108672 800 108792
rect 0 107992 800 108112
rect 0 107312 800 107432
rect 352679 107448 353479 107568
rect 0 106496 800 106616
rect 0 105816 800 105936
rect 352679 105680 353479 105800
rect 0 105136 800 105256
rect 0 104456 800 104576
rect 0 103776 800 103896
rect 352679 103912 353479 104032
rect 0 103096 800 103216
rect 0 102280 800 102400
rect 352679 102144 353479 102264
rect 0 101600 800 101720
rect 0 100920 800 101040
rect 0 100240 800 100360
rect 352679 100376 353479 100496
rect 0 99560 800 99680
rect 0 98744 800 98864
rect 352679 98608 353479 98728
rect 0 98064 800 98184
rect 0 97384 800 97504
rect 0 96704 800 96824
rect 352679 96840 353479 96960
rect 0 96024 800 96144
rect 0 95344 800 95464
rect 352679 94936 353479 95056
rect 0 94528 800 94648
rect 0 93848 800 93968
rect 0 93168 800 93288
rect 352679 93168 353479 93288
rect 0 92488 800 92608
rect 0 91808 800 91928
rect 352679 91400 353479 91520
rect 0 90992 800 91112
rect 0 90312 800 90432
rect 0 89632 800 89752
rect 352679 89632 353479 89752
rect 0 88952 800 89072
rect 0 88272 800 88392
rect 352679 87864 353479 87984
rect 0 87592 800 87712
rect 0 86776 800 86896
rect 0 86096 800 86216
rect 352679 86096 353479 86216
rect 0 85416 800 85536
rect 0 84736 800 84856
rect 352679 84328 353479 84448
rect 0 84056 800 84176
rect 0 83376 800 83496
rect 0 82560 800 82680
rect 352679 82560 353479 82680
rect 0 81880 800 82000
rect 0 81200 800 81320
rect 352679 80792 353479 80912
rect 0 80520 800 80640
rect 0 79840 800 79960
rect 0 79024 800 79144
rect 352679 79024 353479 79144
rect 0 78344 800 78464
rect 0 77664 800 77784
rect 352679 77256 353479 77376
rect 0 76984 800 77104
rect 0 76304 800 76424
rect 0 75624 800 75744
rect 352679 75488 353479 75608
rect 0 74808 800 74928
rect 0 74128 800 74248
rect 352679 73720 353479 73840
rect 0 73448 800 73568
rect 0 72768 800 72888
rect 0 72088 800 72208
rect 352679 71952 353479 72072
rect 0 71408 800 71528
rect 0 70592 800 70712
rect 0 69912 800 70032
rect 352679 70048 353479 70168
rect 0 69232 800 69352
rect 0 68552 800 68672
rect 352679 68280 353479 68400
rect 0 67872 800 67992
rect 0 67056 800 67176
rect 0 66376 800 66496
rect 352679 66512 353479 66632
rect 0 65696 800 65816
rect 0 65016 800 65136
rect 352679 64744 353479 64864
rect 0 64336 800 64456
rect 0 63656 800 63776
rect 0 62840 800 62960
rect 352679 62976 353479 63096
rect 0 62160 800 62280
rect 0 61480 800 61600
rect 352679 61208 353479 61328
rect 0 60800 800 60920
rect 0 60120 800 60240
rect 0 59304 800 59424
rect 352679 59440 353479 59560
rect 0 58624 800 58744
rect 0 57944 800 58064
rect 352679 57672 353479 57792
rect 0 57264 800 57384
rect 0 56584 800 56704
rect 0 55904 800 56024
rect 352679 55904 353479 56024
rect 0 55088 800 55208
rect 0 54408 800 54528
rect 352679 54136 353479 54256
rect 0 53728 800 53848
rect 0 53048 800 53168
rect 0 52368 800 52488
rect 352679 52368 353479 52488
rect 0 51688 800 51808
rect 0 50872 800 50992
rect 352679 50600 353479 50720
rect 0 50192 800 50312
rect 0 49512 800 49632
rect 0 48832 800 48952
rect 352679 48832 353479 48952
rect 0 48152 800 48272
rect 0 47336 800 47456
rect 352679 46928 353479 47048
rect 0 46656 800 46776
rect 0 45976 800 46096
rect 0 45296 800 45416
rect 352679 45160 353479 45280
rect 0 44616 800 44736
rect 0 43936 800 44056
rect 352679 43392 353479 43512
rect 0 43120 800 43240
rect 0 42440 800 42560
rect 0 41760 800 41880
rect 352679 41624 353479 41744
rect 0 41080 800 41200
rect 0 40400 800 40520
rect 352679 39856 353479 39976
rect 0 39584 800 39704
rect 0 38904 800 39024
rect 0 38224 800 38344
rect 352679 38088 353479 38208
rect 0 37544 800 37664
rect 0 36864 800 36984
rect 0 36184 800 36304
rect 352679 36320 353479 36440
rect 0 35368 800 35488
rect 0 34688 800 34808
rect 352679 34552 353479 34672
rect 0 34008 800 34128
rect 0 33328 800 33448
rect 0 32648 800 32768
rect 352679 32784 353479 32904
rect 0 31968 800 32088
rect 0 31152 800 31272
rect 352679 31016 353479 31136
rect 0 30472 800 30592
rect 0 29792 800 29912
rect 0 29112 800 29232
rect 352679 29248 353479 29368
rect 0 28432 800 28552
rect 0 27616 800 27736
rect 352679 27480 353479 27600
rect 0 26936 800 27056
rect 0 26256 800 26376
rect 0 25576 800 25696
rect 352679 25712 353479 25832
rect 0 24896 800 25016
rect 0 24216 800 24336
rect 352679 23808 353479 23928
rect 0 23400 800 23520
rect 0 22720 800 22840
rect 0 22040 800 22160
rect 352679 22040 353479 22160
rect 0 21360 800 21480
rect 0 20680 800 20800
rect 352679 20272 353479 20392
rect 0 19864 800 19984
rect 0 19184 800 19304
rect 0 18504 800 18624
rect 352679 18504 353479 18624
rect 0 17824 800 17944
rect 0 17144 800 17264
rect 352679 16736 353479 16856
rect 0 16464 800 16584
rect 0 15648 800 15768
rect 0 14968 800 15088
rect 352679 14968 353479 15088
rect 0 14288 800 14408
rect 0 13608 800 13728
rect 352679 13200 353479 13320
rect 0 12928 800 13048
rect 0 12248 800 12368
rect 0 11432 800 11552
rect 352679 11432 353479 11552
rect 0 10752 800 10872
rect 0 10072 800 10192
rect 352679 9664 353479 9784
rect 0 9392 800 9512
rect 0 8712 800 8832
rect 0 7896 800 8016
rect 352679 7896 353479 8016
rect 0 7216 800 7336
rect 0 6536 800 6656
rect 352679 6128 353479 6248
rect 0 5856 800 5976
rect 0 5176 800 5296
rect 0 4496 800 4616
rect 352679 4360 353479 4480
rect 0 3680 800 3800
rect 0 3000 800 3120
rect 352679 2592 353479 2712
rect 0 2320 800 2440
rect 0 1640 800 1760
rect 0 960 800 1080
rect 352679 824 353479 944
rect 0 280 800 400
<< obsm3 >>
rect 289 354624 352599 354653
rect 880 354480 352599 354624
rect 880 354344 353451 354480
rect 289 353944 353451 354344
rect 880 353664 353451 353944
rect 289 353264 353451 353664
rect 880 352992 353451 353264
rect 880 352984 352599 352992
rect 289 352712 352599 352984
rect 289 352584 353451 352712
rect 880 352304 353451 352584
rect 289 351768 353451 352304
rect 880 351488 353451 351768
rect 289 351224 353451 351488
rect 289 351088 352599 351224
rect 880 350944 352599 351088
rect 880 350808 353451 350944
rect 289 350408 353451 350808
rect 880 350128 353451 350408
rect 289 349728 353451 350128
rect 880 349456 353451 349728
rect 880 349448 352599 349456
rect 289 349176 352599 349448
rect 289 349048 353451 349176
rect 880 348768 353451 349048
rect 289 348368 353451 348768
rect 880 348088 353451 348368
rect 289 347688 353451 348088
rect 289 347552 352599 347688
rect 880 347408 352599 347552
rect 880 347272 353451 347408
rect 289 346872 353451 347272
rect 880 346592 353451 346872
rect 289 346192 353451 346592
rect 880 345920 353451 346192
rect 880 345912 352599 345920
rect 289 345640 352599 345912
rect 289 345512 353451 345640
rect 880 345232 353451 345512
rect 289 344832 353451 345232
rect 880 344552 353451 344832
rect 289 344152 353451 344552
rect 289 344016 352599 344152
rect 880 343872 352599 344016
rect 880 343736 353451 343872
rect 289 343336 353451 343736
rect 880 343056 353451 343336
rect 289 342656 353451 343056
rect 880 342384 353451 342656
rect 880 342376 352599 342384
rect 289 342104 352599 342376
rect 289 341976 353451 342104
rect 880 341696 353451 341976
rect 289 341296 353451 341696
rect 880 341016 353451 341296
rect 289 340616 353451 341016
rect 880 340336 352599 340616
rect 289 339800 353451 340336
rect 880 339520 353451 339800
rect 289 339120 353451 339520
rect 880 338848 353451 339120
rect 880 338840 352599 338848
rect 289 338568 352599 338840
rect 289 338440 353451 338568
rect 880 338160 353451 338440
rect 289 337760 353451 338160
rect 880 337480 353451 337760
rect 289 337080 353451 337480
rect 880 336800 352599 337080
rect 289 336400 353451 336800
rect 880 336120 353451 336400
rect 289 335584 353451 336120
rect 880 335312 353451 335584
rect 880 335304 352599 335312
rect 289 335032 352599 335304
rect 289 334904 353451 335032
rect 880 334624 353451 334904
rect 289 334224 353451 334624
rect 880 333944 353451 334224
rect 289 333544 353451 333944
rect 880 333264 352599 333544
rect 289 332864 353451 333264
rect 880 332584 353451 332864
rect 289 332048 353451 332584
rect 880 331768 353451 332048
rect 289 331640 353451 331768
rect 289 331368 352599 331640
rect 880 331360 352599 331368
rect 880 331088 353451 331360
rect 289 330688 353451 331088
rect 880 330408 353451 330688
rect 289 330008 353451 330408
rect 880 329872 353451 330008
rect 880 329728 352599 329872
rect 289 329592 352599 329728
rect 289 329328 353451 329592
rect 880 329048 353451 329328
rect 289 328648 353451 329048
rect 880 328368 353451 328648
rect 289 328104 353451 328368
rect 289 327832 352599 328104
rect 880 327824 352599 327832
rect 880 327552 353451 327824
rect 289 327152 353451 327552
rect 880 326872 353451 327152
rect 289 326472 353451 326872
rect 880 326336 353451 326472
rect 880 326192 352599 326336
rect 289 326056 352599 326192
rect 289 325792 353451 326056
rect 880 325512 353451 325792
rect 289 325112 353451 325512
rect 880 324832 353451 325112
rect 289 324568 353451 324832
rect 289 324296 352599 324568
rect 880 324288 352599 324296
rect 880 324016 353451 324288
rect 289 323616 353451 324016
rect 880 323336 353451 323616
rect 289 322936 353451 323336
rect 880 322800 353451 322936
rect 880 322656 352599 322800
rect 289 322520 352599 322656
rect 289 322256 353451 322520
rect 880 321976 353451 322256
rect 289 321576 353451 321976
rect 880 321296 353451 321576
rect 289 321032 353451 321296
rect 289 320896 352599 321032
rect 880 320752 352599 320896
rect 880 320616 353451 320752
rect 289 320080 353451 320616
rect 880 319800 353451 320080
rect 289 319400 353451 319800
rect 880 319264 353451 319400
rect 880 319120 352599 319264
rect 289 318984 352599 319120
rect 289 318720 353451 318984
rect 880 318440 353451 318720
rect 289 318040 353451 318440
rect 880 317760 353451 318040
rect 289 317496 353451 317760
rect 289 317360 352599 317496
rect 880 317216 352599 317360
rect 880 317080 353451 317216
rect 289 316680 353451 317080
rect 880 316400 353451 316680
rect 289 315864 353451 316400
rect 880 315728 353451 315864
rect 880 315584 352599 315728
rect 289 315448 352599 315584
rect 289 315184 353451 315448
rect 880 314904 353451 315184
rect 289 314504 353451 314904
rect 880 314224 353451 314504
rect 289 313960 353451 314224
rect 289 313824 352599 313960
rect 880 313680 352599 313824
rect 880 313544 353451 313680
rect 289 313144 353451 313544
rect 880 312864 353451 313144
rect 289 312328 353451 312864
rect 880 312192 353451 312328
rect 880 312048 352599 312192
rect 289 311912 352599 312048
rect 289 311648 353451 311912
rect 880 311368 353451 311648
rect 289 310968 353451 311368
rect 880 310688 353451 310968
rect 289 310424 353451 310688
rect 289 310288 352599 310424
rect 880 310144 352599 310288
rect 880 310008 353451 310144
rect 289 309608 353451 310008
rect 880 309328 353451 309608
rect 289 308928 353451 309328
rect 880 308648 353451 308928
rect 289 308520 353451 308648
rect 289 308240 352599 308520
rect 289 308112 353451 308240
rect 880 307832 353451 308112
rect 289 307432 353451 307832
rect 880 307152 353451 307432
rect 289 306752 353451 307152
rect 880 306472 352599 306752
rect 289 306072 353451 306472
rect 880 305792 353451 306072
rect 289 305392 353451 305792
rect 880 305112 353451 305392
rect 289 304984 353451 305112
rect 289 304704 352599 304984
rect 289 304576 353451 304704
rect 880 304296 353451 304576
rect 289 303896 353451 304296
rect 880 303616 353451 303896
rect 289 303216 353451 303616
rect 880 302936 352599 303216
rect 289 302536 353451 302936
rect 880 302256 353451 302536
rect 289 301856 353451 302256
rect 880 301576 353451 301856
rect 289 301448 353451 301576
rect 289 301176 352599 301448
rect 880 301168 352599 301176
rect 880 300896 353451 301168
rect 289 300360 353451 300896
rect 880 300080 353451 300360
rect 289 299680 353451 300080
rect 880 299400 352599 299680
rect 289 299000 353451 299400
rect 880 298720 353451 299000
rect 289 298320 353451 298720
rect 880 298040 353451 298320
rect 289 297912 353451 298040
rect 289 297640 352599 297912
rect 880 297632 352599 297640
rect 880 297360 353451 297632
rect 289 296960 353451 297360
rect 880 296680 353451 296960
rect 289 296144 353451 296680
rect 880 295864 352599 296144
rect 289 295464 353451 295864
rect 880 295184 353451 295464
rect 289 294784 353451 295184
rect 880 294504 353451 294784
rect 289 294376 353451 294504
rect 289 294104 352599 294376
rect 880 294096 352599 294104
rect 880 293824 353451 294096
rect 289 293424 353451 293824
rect 880 293144 353451 293424
rect 289 292608 353451 293144
rect 880 292328 352599 292608
rect 289 291928 353451 292328
rect 880 291648 353451 291928
rect 289 291248 353451 291648
rect 880 290968 353451 291248
rect 289 290840 353451 290968
rect 289 290568 352599 290840
rect 880 290560 352599 290568
rect 880 290288 353451 290560
rect 289 289888 353451 290288
rect 880 289608 353451 289888
rect 289 289208 353451 289608
rect 880 289072 353451 289208
rect 880 288928 352599 289072
rect 289 288792 352599 288928
rect 289 288392 353451 288792
rect 880 288112 353451 288392
rect 289 287712 353451 288112
rect 880 287432 353451 287712
rect 289 287304 353451 287432
rect 289 287032 352599 287304
rect 880 287024 352599 287032
rect 880 286752 353451 287024
rect 289 286352 353451 286752
rect 880 286072 353451 286352
rect 289 285672 353451 286072
rect 880 285536 353451 285672
rect 880 285392 352599 285536
rect 289 285256 352599 285392
rect 289 284992 353451 285256
rect 880 284712 353451 284992
rect 289 284176 353451 284712
rect 880 283896 353451 284176
rect 289 283632 353451 283896
rect 289 283496 352599 283632
rect 880 283352 352599 283496
rect 880 283216 353451 283352
rect 289 282816 353451 283216
rect 880 282536 353451 282816
rect 289 282136 353451 282536
rect 880 281864 353451 282136
rect 880 281856 352599 281864
rect 289 281584 352599 281856
rect 289 281456 353451 281584
rect 880 281176 353451 281456
rect 289 280640 353451 281176
rect 880 280360 353451 280640
rect 289 280096 353451 280360
rect 289 279960 352599 280096
rect 880 279816 352599 279960
rect 880 279680 353451 279816
rect 289 279280 353451 279680
rect 880 279000 353451 279280
rect 289 278600 353451 279000
rect 880 278328 353451 278600
rect 880 278320 352599 278328
rect 289 278048 352599 278320
rect 289 277920 353451 278048
rect 880 277640 353451 277920
rect 289 277240 353451 277640
rect 880 276960 353451 277240
rect 289 276560 353451 276960
rect 289 276424 352599 276560
rect 880 276280 352599 276424
rect 880 276144 353451 276280
rect 289 275744 353451 276144
rect 880 275464 353451 275744
rect 289 275064 353451 275464
rect 880 274792 353451 275064
rect 880 274784 352599 274792
rect 289 274512 352599 274784
rect 289 274384 353451 274512
rect 880 274104 353451 274384
rect 289 273704 353451 274104
rect 880 273424 353451 273704
rect 289 273024 353451 273424
rect 289 272888 352599 273024
rect 880 272744 352599 272888
rect 880 272608 353451 272744
rect 289 272208 353451 272608
rect 880 271928 353451 272208
rect 289 271528 353451 271928
rect 880 271256 353451 271528
rect 880 271248 352599 271256
rect 289 270976 352599 271248
rect 289 270848 353451 270976
rect 880 270568 353451 270848
rect 289 270168 353451 270568
rect 880 269888 353451 270168
rect 289 269488 353451 269888
rect 880 269208 352599 269488
rect 289 268672 353451 269208
rect 880 268392 353451 268672
rect 289 267992 353451 268392
rect 880 267720 353451 267992
rect 880 267712 352599 267720
rect 289 267440 352599 267712
rect 289 267312 353451 267440
rect 880 267032 353451 267312
rect 289 266632 353451 267032
rect 880 266352 353451 266632
rect 289 265952 353451 266352
rect 880 265672 352599 265952
rect 289 265272 353451 265672
rect 880 264992 353451 265272
rect 289 264456 353451 264992
rect 880 264184 353451 264456
rect 880 264176 352599 264184
rect 289 263904 352599 264176
rect 289 263776 353451 263904
rect 880 263496 353451 263776
rect 289 263096 353451 263496
rect 880 262816 353451 263096
rect 289 262416 353451 262816
rect 880 262136 352599 262416
rect 289 261736 353451 262136
rect 880 261456 353451 261736
rect 289 260920 353451 261456
rect 880 260640 353451 260920
rect 289 260512 353451 260640
rect 289 260240 352599 260512
rect 880 260232 352599 260240
rect 880 259960 353451 260232
rect 289 259560 353451 259960
rect 880 259280 353451 259560
rect 289 258880 353451 259280
rect 880 258744 353451 258880
rect 880 258600 352599 258744
rect 289 258464 352599 258600
rect 289 258200 353451 258464
rect 880 257920 353451 258200
rect 289 257520 353451 257920
rect 880 257240 353451 257520
rect 289 256976 353451 257240
rect 289 256704 352599 256976
rect 880 256696 352599 256704
rect 880 256424 353451 256696
rect 289 256024 353451 256424
rect 880 255744 353451 256024
rect 289 255344 353451 255744
rect 880 255208 353451 255344
rect 880 255064 352599 255208
rect 289 254928 352599 255064
rect 289 254664 353451 254928
rect 880 254384 353451 254664
rect 289 253984 353451 254384
rect 880 253704 353451 253984
rect 289 253440 353451 253704
rect 289 253168 352599 253440
rect 880 253160 352599 253168
rect 880 252888 353451 253160
rect 289 252488 353451 252888
rect 880 252208 353451 252488
rect 289 251808 353451 252208
rect 880 251672 353451 251808
rect 880 251528 352599 251672
rect 289 251392 352599 251528
rect 289 251128 353451 251392
rect 880 250848 353451 251128
rect 289 250448 353451 250848
rect 880 250168 353451 250448
rect 289 249904 353451 250168
rect 289 249768 352599 249904
rect 880 249624 352599 249768
rect 880 249488 353451 249624
rect 289 248952 353451 249488
rect 880 248672 353451 248952
rect 289 248272 353451 248672
rect 880 248136 353451 248272
rect 880 247992 352599 248136
rect 289 247856 352599 247992
rect 289 247592 353451 247856
rect 880 247312 353451 247592
rect 289 246912 353451 247312
rect 880 246632 353451 246912
rect 289 246368 353451 246632
rect 289 246232 352599 246368
rect 880 246088 352599 246232
rect 880 245952 353451 246088
rect 289 245552 353451 245952
rect 880 245272 353451 245552
rect 289 244736 353451 245272
rect 880 244600 353451 244736
rect 880 244456 352599 244600
rect 289 244320 352599 244456
rect 289 244056 353451 244320
rect 880 243776 353451 244056
rect 289 243376 353451 243776
rect 880 243096 353451 243376
rect 289 242832 353451 243096
rect 289 242696 352599 242832
rect 880 242552 352599 242696
rect 880 242416 353451 242552
rect 289 242016 353451 242416
rect 880 241736 353451 242016
rect 289 241200 353451 241736
rect 880 241064 353451 241200
rect 880 240920 352599 241064
rect 289 240784 352599 240920
rect 289 240520 353451 240784
rect 880 240240 353451 240520
rect 289 239840 353451 240240
rect 880 239560 353451 239840
rect 289 239296 353451 239560
rect 289 239160 352599 239296
rect 880 239016 352599 239160
rect 880 238880 353451 239016
rect 289 238480 353451 238880
rect 880 238200 353451 238480
rect 289 237800 353451 238200
rect 880 237520 353451 237800
rect 289 237392 353451 237520
rect 289 237112 352599 237392
rect 289 236984 353451 237112
rect 880 236704 353451 236984
rect 289 236304 353451 236704
rect 880 236024 353451 236304
rect 289 235624 353451 236024
rect 880 235344 352599 235624
rect 289 234944 353451 235344
rect 880 234664 353451 234944
rect 289 234264 353451 234664
rect 880 233984 353451 234264
rect 289 233856 353451 233984
rect 289 233576 352599 233856
rect 289 233448 353451 233576
rect 880 233168 353451 233448
rect 289 232768 353451 233168
rect 880 232488 353451 232768
rect 289 232088 353451 232488
rect 880 231808 352599 232088
rect 289 231408 353451 231808
rect 880 231128 353451 231408
rect 289 230728 353451 231128
rect 880 230448 353451 230728
rect 289 230320 353451 230448
rect 289 230048 352599 230320
rect 880 230040 352599 230048
rect 880 229768 353451 230040
rect 289 229232 353451 229768
rect 880 228952 353451 229232
rect 289 228552 353451 228952
rect 880 228272 352599 228552
rect 289 227872 353451 228272
rect 880 227592 353451 227872
rect 289 227192 353451 227592
rect 880 226912 353451 227192
rect 289 226784 353451 226912
rect 289 226512 352599 226784
rect 880 226504 352599 226512
rect 880 226232 353451 226504
rect 289 225832 353451 226232
rect 880 225552 353451 225832
rect 289 225016 353451 225552
rect 880 224736 352599 225016
rect 289 224336 353451 224736
rect 880 224056 353451 224336
rect 289 223656 353451 224056
rect 880 223376 353451 223656
rect 289 223248 353451 223376
rect 289 222976 352599 223248
rect 880 222968 352599 222976
rect 880 222696 353451 222968
rect 289 222296 353451 222696
rect 880 222016 353451 222296
rect 289 221480 353451 222016
rect 880 221200 352599 221480
rect 289 220800 353451 221200
rect 880 220520 353451 220800
rect 289 220120 353451 220520
rect 880 219840 353451 220120
rect 289 219712 353451 219840
rect 289 219440 352599 219712
rect 880 219432 352599 219440
rect 880 219160 353451 219432
rect 289 218760 353451 219160
rect 880 218480 353451 218760
rect 289 218080 353451 218480
rect 880 217944 353451 218080
rect 880 217800 352599 217944
rect 289 217664 352599 217800
rect 289 217264 353451 217664
rect 880 216984 353451 217264
rect 289 216584 353451 216984
rect 880 216304 353451 216584
rect 289 216176 353451 216304
rect 289 215904 352599 216176
rect 880 215896 352599 215904
rect 880 215624 353451 215896
rect 289 215224 353451 215624
rect 880 214944 353451 215224
rect 289 214544 353451 214944
rect 880 214408 353451 214544
rect 880 214264 352599 214408
rect 289 214128 352599 214264
rect 289 213864 353451 214128
rect 880 213584 353451 213864
rect 289 213048 353451 213584
rect 880 212768 353451 213048
rect 289 212504 353451 212768
rect 289 212368 352599 212504
rect 880 212224 352599 212368
rect 880 212088 353451 212224
rect 289 211688 353451 212088
rect 880 211408 353451 211688
rect 289 211008 353451 211408
rect 880 210736 353451 211008
rect 880 210728 352599 210736
rect 289 210456 352599 210728
rect 289 210328 353451 210456
rect 880 210048 353451 210328
rect 289 209512 353451 210048
rect 880 209232 353451 209512
rect 289 208968 353451 209232
rect 289 208832 352599 208968
rect 880 208688 352599 208832
rect 880 208552 353451 208688
rect 289 208152 353451 208552
rect 880 207872 353451 208152
rect 289 207472 353451 207872
rect 880 207200 353451 207472
rect 880 207192 352599 207200
rect 289 206920 352599 207192
rect 289 206792 353451 206920
rect 880 206512 353451 206792
rect 289 206112 353451 206512
rect 880 205832 353451 206112
rect 289 205432 353451 205832
rect 289 205296 352599 205432
rect 880 205152 352599 205296
rect 880 205016 353451 205152
rect 289 204616 353451 205016
rect 880 204336 353451 204616
rect 289 203936 353451 204336
rect 880 203664 353451 203936
rect 880 203656 352599 203664
rect 289 203384 352599 203656
rect 289 203256 353451 203384
rect 880 202976 353451 203256
rect 289 202576 353451 202976
rect 880 202296 353451 202576
rect 289 201896 353451 202296
rect 289 201760 352599 201896
rect 880 201616 352599 201760
rect 880 201480 353451 201616
rect 289 201080 353451 201480
rect 880 200800 353451 201080
rect 289 200400 353451 200800
rect 880 200128 353451 200400
rect 880 200120 352599 200128
rect 289 199848 352599 200120
rect 289 199720 353451 199848
rect 880 199440 353451 199720
rect 289 199040 353451 199440
rect 880 198760 353451 199040
rect 289 198360 353451 198760
rect 880 198080 352599 198360
rect 289 197544 353451 198080
rect 880 197264 353451 197544
rect 289 196864 353451 197264
rect 880 196592 353451 196864
rect 880 196584 352599 196592
rect 289 196312 352599 196584
rect 289 196184 353451 196312
rect 880 195904 353451 196184
rect 289 195504 353451 195904
rect 880 195224 353451 195504
rect 289 194824 353451 195224
rect 880 194544 352599 194824
rect 289 194144 353451 194544
rect 880 193864 353451 194144
rect 289 193328 353451 193864
rect 880 193056 353451 193328
rect 880 193048 352599 193056
rect 289 192776 352599 193048
rect 289 192648 353451 192776
rect 880 192368 353451 192648
rect 289 191968 353451 192368
rect 880 191688 353451 191968
rect 289 191288 353451 191688
rect 880 191008 352599 191288
rect 289 190608 353451 191008
rect 880 190328 353451 190608
rect 289 189792 353451 190328
rect 880 189512 353451 189792
rect 289 189384 353451 189512
rect 289 189112 352599 189384
rect 880 189104 352599 189112
rect 880 188832 353451 189104
rect 289 188432 353451 188832
rect 880 188152 353451 188432
rect 289 187752 353451 188152
rect 880 187616 353451 187752
rect 880 187472 352599 187616
rect 289 187336 352599 187472
rect 289 187072 353451 187336
rect 880 186792 353451 187072
rect 289 186392 353451 186792
rect 880 186112 353451 186392
rect 289 185848 353451 186112
rect 289 185576 352599 185848
rect 880 185568 352599 185576
rect 880 185296 353451 185568
rect 289 184896 353451 185296
rect 880 184616 353451 184896
rect 289 184216 353451 184616
rect 880 184080 353451 184216
rect 880 183936 352599 184080
rect 289 183800 352599 183936
rect 289 183536 353451 183800
rect 880 183256 353451 183536
rect 289 182856 353451 183256
rect 880 182576 353451 182856
rect 289 182312 353451 182576
rect 289 182040 352599 182312
rect 880 182032 352599 182040
rect 880 181760 353451 182032
rect 289 181360 353451 181760
rect 880 181080 353451 181360
rect 289 180680 353451 181080
rect 880 180544 353451 180680
rect 880 180400 352599 180544
rect 289 180264 352599 180400
rect 289 180000 353451 180264
rect 880 179720 353451 180000
rect 289 179320 353451 179720
rect 880 179040 353451 179320
rect 289 178776 353451 179040
rect 289 178640 352599 178776
rect 880 178496 352599 178640
rect 880 178360 353451 178496
rect 289 177824 353451 178360
rect 880 177544 353451 177824
rect 289 177144 353451 177544
rect 880 177008 353451 177144
rect 880 176864 352599 177008
rect 289 176728 352599 176864
rect 289 176464 353451 176728
rect 880 176184 353451 176464
rect 289 175784 353451 176184
rect 880 175504 353451 175784
rect 289 175240 353451 175504
rect 289 175104 352599 175240
rect 880 174960 352599 175104
rect 880 174824 353451 174960
rect 289 174424 353451 174824
rect 880 174144 353451 174424
rect 289 173608 353451 174144
rect 880 173472 353451 173608
rect 880 173328 352599 173472
rect 289 173192 352599 173328
rect 289 172928 353451 173192
rect 880 172648 353451 172928
rect 289 172248 353451 172648
rect 880 171968 353451 172248
rect 289 171704 353451 171968
rect 289 171568 352599 171704
rect 880 171424 352599 171568
rect 880 171288 353451 171424
rect 289 170888 353451 171288
rect 880 170608 353451 170888
rect 289 170072 353451 170608
rect 880 169936 353451 170072
rect 880 169792 352599 169936
rect 289 169656 352599 169792
rect 289 169392 353451 169656
rect 880 169112 353451 169392
rect 289 168712 353451 169112
rect 880 168432 353451 168712
rect 289 168168 353451 168432
rect 289 168032 352599 168168
rect 880 167888 352599 168032
rect 880 167752 353451 167888
rect 289 167352 353451 167752
rect 880 167072 353451 167352
rect 289 166672 353451 167072
rect 880 166392 353451 166672
rect 289 166264 353451 166392
rect 289 165984 352599 166264
rect 289 165856 353451 165984
rect 880 165576 353451 165856
rect 289 165176 353451 165576
rect 880 164896 353451 165176
rect 289 164496 353451 164896
rect 880 164216 352599 164496
rect 289 163816 353451 164216
rect 880 163536 353451 163816
rect 289 163136 353451 163536
rect 880 162856 353451 163136
rect 289 162728 353451 162856
rect 289 162448 352599 162728
rect 289 162320 353451 162448
rect 880 162040 353451 162320
rect 289 161640 353451 162040
rect 880 161360 353451 161640
rect 289 160960 353451 161360
rect 880 160680 352599 160960
rect 289 160280 353451 160680
rect 880 160000 353451 160280
rect 289 159600 353451 160000
rect 880 159320 353451 159600
rect 289 159192 353451 159320
rect 289 158920 352599 159192
rect 880 158912 352599 158920
rect 880 158640 353451 158912
rect 289 158104 353451 158640
rect 880 157824 353451 158104
rect 289 157424 353451 157824
rect 880 157144 352599 157424
rect 289 156744 353451 157144
rect 880 156464 353451 156744
rect 289 156064 353451 156464
rect 880 155784 353451 156064
rect 289 155656 353451 155784
rect 289 155384 352599 155656
rect 880 155376 352599 155384
rect 880 155104 353451 155376
rect 289 154704 353451 155104
rect 880 154424 353451 154704
rect 289 153888 353451 154424
rect 880 153608 352599 153888
rect 289 153208 353451 153608
rect 880 152928 353451 153208
rect 289 152528 353451 152928
rect 880 152248 353451 152528
rect 289 152120 353451 152248
rect 289 151848 352599 152120
rect 880 151840 352599 151848
rect 880 151568 353451 151840
rect 289 151168 353451 151568
rect 880 150888 353451 151168
rect 289 150352 353451 150888
rect 880 150072 352599 150352
rect 289 149672 353451 150072
rect 880 149392 353451 149672
rect 289 148992 353451 149392
rect 880 148712 353451 148992
rect 289 148584 353451 148712
rect 289 148312 352599 148584
rect 880 148304 352599 148312
rect 880 148032 353451 148304
rect 289 147632 353451 148032
rect 880 147352 353451 147632
rect 289 146952 353451 147352
rect 880 146816 353451 146952
rect 880 146672 352599 146816
rect 289 146536 352599 146672
rect 289 146136 353451 146536
rect 880 145856 353451 146136
rect 289 145456 353451 145856
rect 880 145176 353451 145456
rect 289 145048 353451 145176
rect 289 144776 352599 145048
rect 880 144768 352599 144776
rect 880 144496 353451 144768
rect 289 144096 353451 144496
rect 880 143816 353451 144096
rect 289 143416 353451 143816
rect 880 143280 353451 143416
rect 880 143136 352599 143280
rect 289 143000 352599 143136
rect 289 142736 353451 143000
rect 880 142456 353451 142736
rect 289 141920 353451 142456
rect 880 141640 353451 141920
rect 289 141376 353451 141640
rect 289 141240 352599 141376
rect 880 141096 352599 141240
rect 880 140960 353451 141096
rect 289 140560 353451 140960
rect 880 140280 353451 140560
rect 289 139880 353451 140280
rect 880 139608 353451 139880
rect 880 139600 352599 139608
rect 289 139328 352599 139600
rect 289 139200 353451 139328
rect 880 138920 353451 139200
rect 289 138384 353451 138920
rect 880 138104 353451 138384
rect 289 137840 353451 138104
rect 289 137704 352599 137840
rect 880 137560 352599 137704
rect 880 137424 353451 137560
rect 289 137024 353451 137424
rect 880 136744 353451 137024
rect 289 136344 353451 136744
rect 880 136072 353451 136344
rect 880 136064 352599 136072
rect 289 135792 352599 136064
rect 289 135664 353451 135792
rect 880 135384 353451 135664
rect 289 134984 353451 135384
rect 880 134704 353451 134984
rect 289 134304 353451 134704
rect 289 134168 352599 134304
rect 880 134024 352599 134168
rect 880 133888 353451 134024
rect 289 133488 353451 133888
rect 880 133208 353451 133488
rect 289 132808 353451 133208
rect 880 132536 353451 132808
rect 880 132528 352599 132536
rect 289 132256 352599 132528
rect 289 132128 353451 132256
rect 880 131848 353451 132128
rect 289 131448 353451 131848
rect 880 131168 353451 131448
rect 289 130768 353451 131168
rect 289 130632 352599 130768
rect 880 130488 352599 130632
rect 880 130352 353451 130488
rect 289 129952 353451 130352
rect 880 129672 353451 129952
rect 289 129272 353451 129672
rect 880 129000 353451 129272
rect 880 128992 352599 129000
rect 289 128720 352599 128992
rect 289 128592 353451 128720
rect 880 128312 353451 128592
rect 289 127912 353451 128312
rect 880 127632 353451 127912
rect 289 127232 353451 127632
rect 880 126952 352599 127232
rect 289 126416 353451 126952
rect 880 126136 353451 126416
rect 289 125736 353451 126136
rect 880 125464 353451 125736
rect 880 125456 352599 125464
rect 289 125184 352599 125456
rect 289 125056 353451 125184
rect 880 124776 353451 125056
rect 289 124376 353451 124776
rect 880 124096 353451 124376
rect 289 123696 353451 124096
rect 880 123416 352599 123696
rect 289 123016 353451 123416
rect 880 122736 353451 123016
rect 289 122200 353451 122736
rect 880 121928 353451 122200
rect 880 121920 352599 121928
rect 289 121648 352599 121920
rect 289 121520 353451 121648
rect 880 121240 353451 121520
rect 289 120840 353451 121240
rect 880 120560 353451 120840
rect 289 120160 353451 120560
rect 880 119880 352599 120160
rect 289 119480 353451 119880
rect 880 119200 353451 119480
rect 289 118664 353451 119200
rect 880 118384 353451 118664
rect 289 118256 353451 118384
rect 289 117984 352599 118256
rect 880 117976 352599 117984
rect 880 117704 353451 117976
rect 289 117304 353451 117704
rect 880 117024 353451 117304
rect 289 116624 353451 117024
rect 880 116488 353451 116624
rect 880 116344 352599 116488
rect 289 116208 352599 116344
rect 289 115944 353451 116208
rect 880 115664 353451 115944
rect 289 115264 353451 115664
rect 880 114984 353451 115264
rect 289 114720 353451 114984
rect 289 114448 352599 114720
rect 880 114440 352599 114448
rect 880 114168 353451 114440
rect 289 113768 353451 114168
rect 880 113488 353451 113768
rect 289 113088 353451 113488
rect 880 112952 353451 113088
rect 880 112808 352599 112952
rect 289 112672 352599 112808
rect 289 112408 353451 112672
rect 880 112128 353451 112408
rect 289 111728 353451 112128
rect 880 111448 353451 111728
rect 289 111184 353451 111448
rect 289 110912 352599 111184
rect 880 110904 352599 110912
rect 880 110632 353451 110904
rect 289 110232 353451 110632
rect 880 109952 353451 110232
rect 289 109552 353451 109952
rect 880 109416 353451 109552
rect 880 109272 352599 109416
rect 289 109136 352599 109272
rect 289 108872 353451 109136
rect 880 108592 353451 108872
rect 289 108192 353451 108592
rect 880 107912 353451 108192
rect 289 107648 353451 107912
rect 289 107512 352599 107648
rect 880 107368 352599 107512
rect 880 107232 353451 107368
rect 289 106696 353451 107232
rect 880 106416 353451 106696
rect 289 106016 353451 106416
rect 880 105880 353451 106016
rect 880 105736 352599 105880
rect 289 105600 352599 105736
rect 289 105336 353451 105600
rect 880 105056 353451 105336
rect 289 104656 353451 105056
rect 880 104376 353451 104656
rect 289 104112 353451 104376
rect 289 103976 352599 104112
rect 880 103832 352599 103976
rect 880 103696 353451 103832
rect 289 103296 353451 103696
rect 880 103016 353451 103296
rect 289 102480 353451 103016
rect 880 102344 353451 102480
rect 880 102200 352599 102344
rect 289 102064 352599 102200
rect 289 101800 353451 102064
rect 880 101520 353451 101800
rect 289 101120 353451 101520
rect 880 100840 353451 101120
rect 289 100576 353451 100840
rect 289 100440 352599 100576
rect 880 100296 352599 100440
rect 880 100160 353451 100296
rect 289 99760 353451 100160
rect 880 99480 353451 99760
rect 289 98944 353451 99480
rect 880 98808 353451 98944
rect 880 98664 352599 98808
rect 289 98528 352599 98664
rect 289 98264 353451 98528
rect 880 97984 353451 98264
rect 289 97584 353451 97984
rect 880 97304 353451 97584
rect 289 97040 353451 97304
rect 289 96904 352599 97040
rect 880 96760 352599 96904
rect 880 96624 353451 96760
rect 289 96224 353451 96624
rect 880 95944 353451 96224
rect 289 95544 353451 95944
rect 880 95264 353451 95544
rect 289 95136 353451 95264
rect 289 94856 352599 95136
rect 289 94728 353451 94856
rect 880 94448 353451 94728
rect 289 94048 353451 94448
rect 880 93768 353451 94048
rect 289 93368 353451 93768
rect 880 93088 352599 93368
rect 289 92688 353451 93088
rect 880 92408 353451 92688
rect 289 92008 353451 92408
rect 880 91728 353451 92008
rect 289 91600 353451 91728
rect 289 91320 352599 91600
rect 289 91192 353451 91320
rect 880 90912 353451 91192
rect 289 90512 353451 90912
rect 880 90232 353451 90512
rect 289 89832 353451 90232
rect 880 89552 352599 89832
rect 289 89152 353451 89552
rect 880 88872 353451 89152
rect 289 88472 353451 88872
rect 880 88192 353451 88472
rect 289 88064 353451 88192
rect 289 87792 352599 88064
rect 880 87784 352599 87792
rect 880 87512 353451 87784
rect 289 86976 353451 87512
rect 880 86696 353451 86976
rect 289 86296 353451 86696
rect 880 86016 352599 86296
rect 289 85616 353451 86016
rect 880 85336 353451 85616
rect 289 84936 353451 85336
rect 880 84656 353451 84936
rect 289 84528 353451 84656
rect 289 84256 352599 84528
rect 880 84248 352599 84256
rect 880 83976 353451 84248
rect 289 83576 353451 83976
rect 880 83296 353451 83576
rect 289 82760 353451 83296
rect 880 82480 352599 82760
rect 289 82080 353451 82480
rect 880 81800 353451 82080
rect 289 81400 353451 81800
rect 880 81120 353451 81400
rect 289 80992 353451 81120
rect 289 80720 352599 80992
rect 880 80712 352599 80720
rect 880 80440 353451 80712
rect 289 80040 353451 80440
rect 880 79760 353451 80040
rect 289 79224 353451 79760
rect 880 78944 352599 79224
rect 289 78544 353451 78944
rect 880 78264 353451 78544
rect 289 77864 353451 78264
rect 880 77584 353451 77864
rect 289 77456 353451 77584
rect 289 77184 352599 77456
rect 880 77176 352599 77184
rect 880 76904 353451 77176
rect 289 76504 353451 76904
rect 880 76224 353451 76504
rect 289 75824 353451 76224
rect 880 75688 353451 75824
rect 880 75544 352599 75688
rect 289 75408 352599 75544
rect 289 75008 353451 75408
rect 880 74728 353451 75008
rect 289 74328 353451 74728
rect 880 74048 353451 74328
rect 289 73920 353451 74048
rect 289 73648 352599 73920
rect 880 73640 352599 73648
rect 880 73368 353451 73640
rect 289 72968 353451 73368
rect 880 72688 353451 72968
rect 289 72288 353451 72688
rect 880 72152 353451 72288
rect 880 72008 352599 72152
rect 289 71872 352599 72008
rect 289 71608 353451 71872
rect 880 71328 353451 71608
rect 289 70792 353451 71328
rect 880 70512 353451 70792
rect 289 70248 353451 70512
rect 289 70112 352599 70248
rect 880 69968 352599 70112
rect 880 69832 353451 69968
rect 289 69432 353451 69832
rect 880 69152 353451 69432
rect 289 68752 353451 69152
rect 880 68480 353451 68752
rect 880 68472 352599 68480
rect 289 68200 352599 68472
rect 289 68072 353451 68200
rect 880 67792 353451 68072
rect 289 67256 353451 67792
rect 880 66976 353451 67256
rect 289 66712 353451 66976
rect 289 66576 352599 66712
rect 880 66432 352599 66576
rect 880 66296 353451 66432
rect 289 65896 353451 66296
rect 880 65616 353451 65896
rect 289 65216 353451 65616
rect 880 64944 353451 65216
rect 880 64936 352599 64944
rect 289 64664 352599 64936
rect 289 64536 353451 64664
rect 880 64256 353451 64536
rect 289 63856 353451 64256
rect 880 63576 353451 63856
rect 289 63176 353451 63576
rect 289 63040 352599 63176
rect 880 62896 352599 63040
rect 880 62760 353451 62896
rect 289 62360 353451 62760
rect 880 62080 353451 62360
rect 289 61680 353451 62080
rect 880 61408 353451 61680
rect 880 61400 352599 61408
rect 289 61128 352599 61400
rect 289 61000 353451 61128
rect 880 60720 353451 61000
rect 289 60320 353451 60720
rect 880 60040 353451 60320
rect 289 59640 353451 60040
rect 289 59504 352599 59640
rect 880 59360 352599 59504
rect 880 59224 353451 59360
rect 289 58824 353451 59224
rect 880 58544 353451 58824
rect 289 58144 353451 58544
rect 880 57872 353451 58144
rect 880 57864 352599 57872
rect 289 57592 352599 57864
rect 289 57464 353451 57592
rect 880 57184 353451 57464
rect 289 56784 353451 57184
rect 880 56504 353451 56784
rect 289 56104 353451 56504
rect 880 55824 352599 56104
rect 289 55288 353451 55824
rect 880 55008 353451 55288
rect 289 54608 353451 55008
rect 880 54336 353451 54608
rect 880 54328 352599 54336
rect 289 54056 352599 54328
rect 289 53928 353451 54056
rect 880 53648 353451 53928
rect 289 53248 353451 53648
rect 880 52968 353451 53248
rect 289 52568 353451 52968
rect 880 52288 352599 52568
rect 289 51888 353451 52288
rect 880 51608 353451 51888
rect 289 51072 353451 51608
rect 880 50800 353451 51072
rect 880 50792 352599 50800
rect 289 50520 352599 50792
rect 289 50392 353451 50520
rect 880 50112 353451 50392
rect 289 49712 353451 50112
rect 880 49432 353451 49712
rect 289 49032 353451 49432
rect 880 48752 352599 49032
rect 289 48352 353451 48752
rect 880 48072 353451 48352
rect 289 47536 353451 48072
rect 880 47256 353451 47536
rect 289 47128 353451 47256
rect 289 46856 352599 47128
rect 880 46848 352599 46856
rect 880 46576 353451 46848
rect 289 46176 353451 46576
rect 880 45896 353451 46176
rect 289 45496 353451 45896
rect 880 45360 353451 45496
rect 880 45216 352599 45360
rect 289 45080 352599 45216
rect 289 44816 353451 45080
rect 880 44536 353451 44816
rect 289 44136 353451 44536
rect 880 43856 353451 44136
rect 289 43592 353451 43856
rect 289 43320 352599 43592
rect 880 43312 352599 43320
rect 880 43040 353451 43312
rect 289 42640 353451 43040
rect 880 42360 353451 42640
rect 289 41960 353451 42360
rect 880 41824 353451 41960
rect 880 41680 352599 41824
rect 289 41544 352599 41680
rect 289 41280 353451 41544
rect 880 41000 353451 41280
rect 289 40600 353451 41000
rect 880 40320 353451 40600
rect 289 40056 353451 40320
rect 289 39784 352599 40056
rect 880 39776 352599 39784
rect 880 39504 353451 39776
rect 289 39104 353451 39504
rect 880 38824 353451 39104
rect 289 38424 353451 38824
rect 880 38288 353451 38424
rect 880 38144 352599 38288
rect 289 38008 352599 38144
rect 289 37744 353451 38008
rect 880 37464 353451 37744
rect 289 37064 353451 37464
rect 880 36784 353451 37064
rect 289 36520 353451 36784
rect 289 36384 352599 36520
rect 880 36240 352599 36384
rect 880 36104 353451 36240
rect 289 35568 353451 36104
rect 880 35288 353451 35568
rect 289 34888 353451 35288
rect 880 34752 353451 34888
rect 880 34608 352599 34752
rect 289 34472 352599 34608
rect 289 34208 353451 34472
rect 880 33928 353451 34208
rect 289 33528 353451 33928
rect 880 33248 353451 33528
rect 289 32984 353451 33248
rect 289 32848 352599 32984
rect 880 32704 352599 32848
rect 880 32568 353451 32704
rect 289 32168 353451 32568
rect 880 31888 353451 32168
rect 289 31352 353451 31888
rect 880 31216 353451 31352
rect 880 31072 352599 31216
rect 289 30936 352599 31072
rect 289 30672 353451 30936
rect 880 30392 353451 30672
rect 289 29992 353451 30392
rect 880 29712 353451 29992
rect 289 29448 353451 29712
rect 289 29312 352599 29448
rect 880 29168 352599 29312
rect 880 29032 353451 29168
rect 289 28632 353451 29032
rect 880 28352 353451 28632
rect 289 27816 353451 28352
rect 880 27680 353451 27816
rect 880 27536 352599 27680
rect 289 27400 352599 27536
rect 289 27136 353451 27400
rect 880 26856 353451 27136
rect 289 26456 353451 26856
rect 880 26176 353451 26456
rect 289 25912 353451 26176
rect 289 25776 352599 25912
rect 880 25632 352599 25776
rect 880 25496 353451 25632
rect 289 25096 353451 25496
rect 880 24816 353451 25096
rect 289 24416 353451 24816
rect 880 24136 353451 24416
rect 289 24008 353451 24136
rect 289 23728 352599 24008
rect 289 23600 353451 23728
rect 880 23320 353451 23600
rect 289 22920 353451 23320
rect 880 22640 353451 22920
rect 289 22240 353451 22640
rect 880 21960 352599 22240
rect 289 21560 353451 21960
rect 880 21280 353451 21560
rect 289 20880 353451 21280
rect 880 20600 353451 20880
rect 289 20472 353451 20600
rect 289 20192 352599 20472
rect 289 20064 353451 20192
rect 880 19784 353451 20064
rect 289 19384 353451 19784
rect 880 19104 353451 19384
rect 289 18704 353451 19104
rect 880 18424 352599 18704
rect 289 18024 353451 18424
rect 880 17744 353451 18024
rect 289 17344 353451 17744
rect 880 17064 353451 17344
rect 289 16936 353451 17064
rect 289 16664 352599 16936
rect 880 16656 352599 16664
rect 880 16384 353451 16656
rect 289 15848 353451 16384
rect 880 15568 353451 15848
rect 289 15168 353451 15568
rect 880 14888 352599 15168
rect 289 14488 353451 14888
rect 880 14208 353451 14488
rect 289 13808 353451 14208
rect 880 13528 353451 13808
rect 289 13400 353451 13528
rect 289 13128 352599 13400
rect 880 13120 352599 13128
rect 880 12848 353451 13120
rect 289 12448 353451 12848
rect 880 12168 353451 12448
rect 289 11632 353451 12168
rect 880 11352 352599 11632
rect 289 10952 353451 11352
rect 880 10672 353451 10952
rect 289 10272 353451 10672
rect 880 9992 353451 10272
rect 289 9864 353451 9992
rect 289 9592 352599 9864
rect 880 9584 352599 9592
rect 880 9312 353451 9584
rect 289 8912 353451 9312
rect 880 8632 353451 8912
rect 289 8096 353451 8632
rect 880 7816 352599 8096
rect 289 7416 353451 7816
rect 880 7136 353451 7416
rect 289 6736 353451 7136
rect 880 6456 353451 6736
rect 289 6328 353451 6456
rect 289 6056 352599 6328
rect 880 6048 352599 6056
rect 880 5776 353451 6048
rect 289 5376 353451 5776
rect 880 5096 353451 5376
rect 289 4696 353451 5096
rect 880 4560 353451 4696
rect 880 4416 352599 4560
rect 289 4280 352599 4416
rect 289 3880 353451 4280
rect 880 3600 353451 3880
rect 289 3200 353451 3600
rect 880 2920 353451 3200
rect 289 2792 353451 2920
rect 289 2520 352599 2792
rect 880 2512 352599 2520
rect 880 2240 353451 2512
rect 289 1840 353451 2240
rect 880 1560 353451 1840
rect 289 1160 353451 1560
rect 880 1024 353451 1160
rect 880 880 352599 1024
rect 289 744 352599 880
rect 289 480 353451 744
rect 880 307 353451 480
<< metal4 >>
rect 4208 2128 4528 353104
rect 19568 2128 19888 353104
rect 34928 2128 35248 353104
rect 50288 2128 50608 353104
rect 65648 2128 65968 353104
rect 81008 2128 81328 353104
rect 96368 2128 96688 353104
rect 111728 2128 112048 353104
rect 127088 2128 127408 353104
rect 142448 2128 142768 353104
rect 157808 2128 158128 353104
rect 173168 2128 173488 353104
rect 188528 2128 188848 353104
rect 203888 2128 204208 353104
rect 219248 2128 219568 353104
rect 234608 2128 234928 353104
rect 249968 2128 250288 353104
rect 265328 2128 265648 353104
rect 280688 2128 281008 353104
rect 296048 2128 296368 353104
rect 311408 2128 311728 353104
rect 326768 2128 327088 353104
rect 342128 2128 342448 353104
<< obsm4 >>
rect 795 353184 353037 353565
rect 795 2048 4128 353184
rect 4608 2048 19488 353184
rect 19968 2048 34848 353184
rect 35328 2048 50208 353184
rect 50688 2048 65568 353184
rect 66048 2048 80928 353184
rect 81408 2048 96288 353184
rect 96768 2048 111648 353184
rect 112128 2048 127008 353184
rect 127488 2048 142368 353184
rect 142848 2048 157728 353184
rect 158208 2048 173088 353184
rect 173568 2048 188448 353184
rect 188928 2048 203808 353184
rect 204288 2048 219168 353184
rect 219648 2048 234528 353184
rect 235008 2048 249888 353184
rect 250368 2048 265248 353184
rect 265728 2048 280608 353184
rect 281088 2048 295968 353184
rect 296448 2048 311328 353184
rect 311808 2048 326688 353184
rect 327168 2048 342048 353184
rect 342528 2048 353037 353184
rect 795 1803 353037 2048
<< labels >>
rlabel metal3 s 0 153008 800 153128 6 data_arrays_0_0_ext_ram_addr1[0]
port 1 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 data_arrays_0_0_ext_ram_addr1[1]
port 2 nsew signal output
rlabel metal3 s 0 154504 800 154624 6 data_arrays_0_0_ext_ram_addr1[2]
port 3 nsew signal output
rlabel metal3 s 0 155184 800 155304 6 data_arrays_0_0_ext_ram_addr1[3]
port 4 nsew signal output
rlabel metal3 s 0 155864 800 155984 6 data_arrays_0_0_ext_ram_addr1[4]
port 5 nsew signal output
rlabel metal3 s 0 156544 800 156664 6 data_arrays_0_0_ext_ram_addr1[5]
port 6 nsew signal output
rlabel metal3 s 0 157224 800 157344 6 data_arrays_0_0_ext_ram_addr1[6]
port 7 nsew signal output
rlabel metal3 s 0 157904 800 158024 6 data_arrays_0_0_ext_ram_addr1[7]
port 8 nsew signal output
rlabel metal3 s 0 158720 800 158840 6 data_arrays_0_0_ext_ram_addr1[8]
port 9 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 data_arrays_0_0_ext_ram_addr[0]
port 10 nsew signal output
rlabel metal3 s 0 90992 800 91112 6 data_arrays_0_0_ext_ram_addr[1]
port 11 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 data_arrays_0_0_ext_ram_addr[2]
port 12 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 data_arrays_0_0_ext_ram_addr[3]
port 13 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 data_arrays_0_0_ext_ram_addr[4]
port 14 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 data_arrays_0_0_ext_ram_addr[5]
port 15 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 data_arrays_0_0_ext_ram_addr[6]
port 16 nsew signal output
rlabel metal3 s 0 95344 800 95464 6 data_arrays_0_0_ext_ram_addr[7]
port 17 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 data_arrays_0_0_ext_ram_addr[8]
port 18 nsew signal output
rlabel metal3 s 0 96704 800 96824 6 data_arrays_0_0_ext_ram_clk
port 19 nsew signal output
rlabel metal3 s 0 147432 800 147552 6 data_arrays_0_0_ext_ram_csb1[0]
port 20 nsew signal output
rlabel metal3 s 0 148112 800 148232 6 data_arrays_0_0_ext_ram_csb1[1]
port 21 nsew signal output
rlabel metal3 s 0 148792 800 148912 6 data_arrays_0_0_ext_ram_csb1[2]
port 22 nsew signal output
rlabel metal3 s 0 149472 800 149592 6 data_arrays_0_0_ext_ram_csb1[3]
port 23 nsew signal output
rlabel metal3 s 0 150152 800 150272 6 data_arrays_0_0_ext_ram_csb1[4]
port 24 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 data_arrays_0_0_ext_ram_csb1[5]
port 25 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 data_arrays_0_0_ext_ram_csb1[6]
port 26 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 data_arrays_0_0_ext_ram_csb1[7]
port 27 nsew signal output
rlabel metal3 s 0 143896 800 144016 6 data_arrays_0_0_ext_ram_csb[0]
port 28 nsew signal output
rlabel metal3 s 0 144576 800 144696 6 data_arrays_0_0_ext_ram_csb[1]
port 29 nsew signal output
rlabel metal3 s 0 145256 800 145376 6 data_arrays_0_0_ext_ram_csb[2]
port 30 nsew signal output
rlabel metal3 s 0 145936 800 146056 6 data_arrays_0_0_ext_ram_csb[3]
port 31 nsew signal output
rlabel metal3 s 0 280 800 400 6 data_arrays_0_0_ext_ram_rdata0[0]
port 32 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 data_arrays_0_0_ext_ram_rdata0[10]
port 33 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 data_arrays_0_0_ext_ram_rdata0[11]
port 34 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 data_arrays_0_0_ext_ram_rdata0[12]
port 35 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 data_arrays_0_0_ext_ram_rdata0[13]
port 36 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 data_arrays_0_0_ext_ram_rdata0[14]
port 37 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 data_arrays_0_0_ext_ram_rdata0[15]
port 38 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 data_arrays_0_0_ext_ram_rdata0[16]
port 39 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 data_arrays_0_0_ext_ram_rdata0[17]
port 40 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 data_arrays_0_0_ext_ram_rdata0[18]
port 41 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 data_arrays_0_0_ext_ram_rdata0[19]
port 42 nsew signal input
rlabel metal3 s 0 960 800 1080 6 data_arrays_0_0_ext_ram_rdata0[1]
port 43 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 data_arrays_0_0_ext_ram_rdata0[20]
port 44 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 data_arrays_0_0_ext_ram_rdata0[21]
port 45 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 data_arrays_0_0_ext_ram_rdata0[22]
port 46 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 data_arrays_0_0_ext_ram_rdata0[23]
port 47 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 data_arrays_0_0_ext_ram_rdata0[24]
port 48 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 data_arrays_0_0_ext_ram_rdata0[25]
port 49 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 data_arrays_0_0_ext_ram_rdata0[26]
port 50 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 data_arrays_0_0_ext_ram_rdata0[27]
port 51 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 data_arrays_0_0_ext_ram_rdata0[28]
port 52 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 data_arrays_0_0_ext_ram_rdata0[29]
port 53 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 data_arrays_0_0_ext_ram_rdata0[2]
port 54 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 data_arrays_0_0_ext_ram_rdata0[30]
port 55 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 data_arrays_0_0_ext_ram_rdata0[31]
port 56 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 data_arrays_0_0_ext_ram_rdata0[32]
port 57 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 data_arrays_0_0_ext_ram_rdata0[33]
port 58 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 data_arrays_0_0_ext_ram_rdata0[34]
port 59 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 data_arrays_0_0_ext_ram_rdata0[35]
port 60 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 data_arrays_0_0_ext_ram_rdata0[36]
port 61 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 data_arrays_0_0_ext_ram_rdata0[37]
port 62 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 data_arrays_0_0_ext_ram_rdata0[38]
port 63 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 data_arrays_0_0_ext_ram_rdata0[39]
port 64 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 data_arrays_0_0_ext_ram_rdata0[3]
port 65 nsew signal input
rlabel metal3 s 0 28432 800 28552 6 data_arrays_0_0_ext_ram_rdata0[40]
port 66 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 data_arrays_0_0_ext_ram_rdata0[41]
port 67 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 data_arrays_0_0_ext_ram_rdata0[42]
port 68 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 data_arrays_0_0_ext_ram_rdata0[43]
port 69 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 data_arrays_0_0_ext_ram_rdata0[44]
port 70 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 data_arrays_0_0_ext_ram_rdata0[45]
port 71 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 data_arrays_0_0_ext_ram_rdata0[46]
port 72 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 data_arrays_0_0_ext_ram_rdata0[47]
port 73 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 data_arrays_0_0_ext_ram_rdata0[48]
port 74 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 data_arrays_0_0_ext_ram_rdata0[49]
port 75 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 data_arrays_0_0_ext_ram_rdata0[4]
port 76 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 data_arrays_0_0_ext_ram_rdata0[50]
port 77 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 data_arrays_0_0_ext_ram_rdata0[51]
port 78 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 data_arrays_0_0_ext_ram_rdata0[52]
port 79 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 data_arrays_0_0_ext_ram_rdata0[53]
port 80 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 data_arrays_0_0_ext_ram_rdata0[54]
port 81 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 data_arrays_0_0_ext_ram_rdata0[55]
port 82 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 data_arrays_0_0_ext_ram_rdata0[56]
port 83 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 data_arrays_0_0_ext_ram_rdata0[57]
port 84 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 data_arrays_0_0_ext_ram_rdata0[58]
port 85 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 data_arrays_0_0_ext_ram_rdata0[59]
port 86 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 data_arrays_0_0_ext_ram_rdata0[5]
port 87 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 data_arrays_0_0_ext_ram_rdata0[60]
port 88 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 data_arrays_0_0_ext_ram_rdata0[61]
port 89 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 data_arrays_0_0_ext_ram_rdata0[62]
port 90 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 data_arrays_0_0_ext_ram_rdata0[63]
port 91 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 data_arrays_0_0_ext_ram_rdata0[6]
port 92 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 data_arrays_0_0_ext_ram_rdata0[7]
port 93 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 data_arrays_0_0_ext_ram_rdata0[8]
port 94 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 data_arrays_0_0_ext_ram_rdata0[9]
port 95 nsew signal input
rlabel metal3 s 0 45296 800 45416 6 data_arrays_0_0_ext_ram_rdata1[0]
port 96 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 data_arrays_0_0_ext_ram_rdata1[10]
port 97 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 data_arrays_0_0_ext_ram_rdata1[11]
port 98 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 data_arrays_0_0_ext_ram_rdata1[12]
port 99 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 data_arrays_0_0_ext_ram_rdata1[13]
port 100 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 data_arrays_0_0_ext_ram_rdata1[14]
port 101 nsew signal input
rlabel metal3 s 0 55904 800 56024 6 data_arrays_0_0_ext_ram_rdata1[15]
port 102 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 data_arrays_0_0_ext_ram_rdata1[16]
port 103 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 data_arrays_0_0_ext_ram_rdata1[17]
port 104 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 data_arrays_0_0_ext_ram_rdata1[18]
port 105 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 data_arrays_0_0_ext_ram_rdata1[19]
port 106 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 data_arrays_0_0_ext_ram_rdata1[1]
port 107 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 data_arrays_0_0_ext_ram_rdata1[20]
port 108 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 data_arrays_0_0_ext_ram_rdata1[21]
port 109 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 data_arrays_0_0_ext_ram_rdata1[22]
port 110 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 data_arrays_0_0_ext_ram_rdata1[23]
port 111 nsew signal input
rlabel metal3 s 0 62160 800 62280 6 data_arrays_0_0_ext_ram_rdata1[24]
port 112 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 data_arrays_0_0_ext_ram_rdata1[25]
port 113 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 data_arrays_0_0_ext_ram_rdata1[26]
port 114 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 data_arrays_0_0_ext_ram_rdata1[27]
port 115 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 data_arrays_0_0_ext_ram_rdata1[28]
port 116 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 data_arrays_0_0_ext_ram_rdata1[29]
port 117 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 data_arrays_0_0_ext_ram_rdata1[2]
port 118 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 data_arrays_0_0_ext_ram_rdata1[30]
port 119 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 data_arrays_0_0_ext_ram_rdata1[31]
port 120 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 data_arrays_0_0_ext_ram_rdata1[32]
port 121 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 data_arrays_0_0_ext_ram_rdata1[33]
port 122 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 data_arrays_0_0_ext_ram_rdata1[34]
port 123 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 data_arrays_0_0_ext_ram_rdata1[35]
port 124 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 data_arrays_0_0_ext_ram_rdata1[36]
port 125 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 data_arrays_0_0_ext_ram_rdata1[37]
port 126 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 data_arrays_0_0_ext_ram_rdata1[38]
port 127 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 data_arrays_0_0_ext_ram_rdata1[39]
port 128 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 data_arrays_0_0_ext_ram_rdata1[3]
port 129 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 data_arrays_0_0_ext_ram_rdata1[40]
port 130 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 data_arrays_0_0_ext_ram_rdata1[41]
port 131 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 data_arrays_0_0_ext_ram_rdata1[42]
port 132 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 data_arrays_0_0_ext_ram_rdata1[43]
port 133 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 data_arrays_0_0_ext_ram_rdata1[44]
port 134 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 data_arrays_0_0_ext_ram_rdata1[45]
port 135 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 data_arrays_0_0_ext_ram_rdata1[46]
port 136 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 data_arrays_0_0_ext_ram_rdata1[47]
port 137 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 data_arrays_0_0_ext_ram_rdata1[48]
port 138 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 data_arrays_0_0_ext_ram_rdata1[49]
port 139 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 data_arrays_0_0_ext_ram_rdata1[4]
port 140 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 data_arrays_0_0_ext_ram_rdata1[50]
port 141 nsew signal input
rlabel metal3 s 0 81200 800 81320 6 data_arrays_0_0_ext_ram_rdata1[51]
port 142 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 data_arrays_0_0_ext_ram_rdata1[52]
port 143 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 data_arrays_0_0_ext_ram_rdata1[53]
port 144 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 data_arrays_0_0_ext_ram_rdata1[54]
port 145 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 data_arrays_0_0_ext_ram_rdata1[55]
port 146 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 data_arrays_0_0_ext_ram_rdata1[56]
port 147 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 data_arrays_0_0_ext_ram_rdata1[57]
port 148 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 data_arrays_0_0_ext_ram_rdata1[58]
port 149 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 data_arrays_0_0_ext_ram_rdata1[59]
port 150 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 data_arrays_0_0_ext_ram_rdata1[5]
port 151 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 data_arrays_0_0_ext_ram_rdata1[60]
port 152 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 data_arrays_0_0_ext_ram_rdata1[61]
port 153 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 data_arrays_0_0_ext_ram_rdata1[62]
port 154 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 data_arrays_0_0_ext_ram_rdata1[63]
port 155 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 data_arrays_0_0_ext_ram_rdata1[6]
port 156 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 data_arrays_0_0_ext_ram_rdata1[7]
port 157 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 data_arrays_0_0_ext_ram_rdata1[8]
port 158 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 data_arrays_0_0_ext_ram_rdata1[9]
port 159 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 data_arrays_0_0_ext_ram_rdata2[0]
port 160 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 data_arrays_0_0_ext_ram_rdata2[10]
port 161 nsew signal input
rlabel metal3 s 0 167152 800 167272 6 data_arrays_0_0_ext_ram_rdata2[11]
port 162 nsew signal input
rlabel metal3 s 0 167832 800 167952 6 data_arrays_0_0_ext_ram_rdata2[12]
port 163 nsew signal input
rlabel metal3 s 0 168512 800 168632 6 data_arrays_0_0_ext_ram_rdata2[13]
port 164 nsew signal input
rlabel metal3 s 0 169192 800 169312 6 data_arrays_0_0_ext_ram_rdata2[14]
port 165 nsew signal input
rlabel metal3 s 0 169872 800 169992 6 data_arrays_0_0_ext_ram_rdata2[15]
port 166 nsew signal input
rlabel metal3 s 0 170688 800 170808 6 data_arrays_0_0_ext_ram_rdata2[16]
port 167 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 data_arrays_0_0_ext_ram_rdata2[17]
port 168 nsew signal input
rlabel metal3 s 0 172048 800 172168 6 data_arrays_0_0_ext_ram_rdata2[18]
port 169 nsew signal input
rlabel metal3 s 0 172728 800 172848 6 data_arrays_0_0_ext_ram_rdata2[19]
port 170 nsew signal input
rlabel metal3 s 0 160080 800 160200 6 data_arrays_0_0_ext_ram_rdata2[1]
port 171 nsew signal input
rlabel metal3 s 0 173408 800 173528 6 data_arrays_0_0_ext_ram_rdata2[20]
port 172 nsew signal input
rlabel metal3 s 0 174224 800 174344 6 data_arrays_0_0_ext_ram_rdata2[21]
port 173 nsew signal input
rlabel metal3 s 0 174904 800 175024 6 data_arrays_0_0_ext_ram_rdata2[22]
port 174 nsew signal input
rlabel metal3 s 0 175584 800 175704 6 data_arrays_0_0_ext_ram_rdata2[23]
port 175 nsew signal input
rlabel metal3 s 0 176264 800 176384 6 data_arrays_0_0_ext_ram_rdata2[24]
port 176 nsew signal input
rlabel metal3 s 0 176944 800 177064 6 data_arrays_0_0_ext_ram_rdata2[25]
port 177 nsew signal input
rlabel metal3 s 0 177624 800 177744 6 data_arrays_0_0_ext_ram_rdata2[26]
port 178 nsew signal input
rlabel metal3 s 0 178440 800 178560 6 data_arrays_0_0_ext_ram_rdata2[27]
port 179 nsew signal input
rlabel metal3 s 0 179120 800 179240 6 data_arrays_0_0_ext_ram_rdata2[28]
port 180 nsew signal input
rlabel metal3 s 0 179800 800 179920 6 data_arrays_0_0_ext_ram_rdata2[29]
port 181 nsew signal input
rlabel metal3 s 0 160760 800 160880 6 data_arrays_0_0_ext_ram_rdata2[2]
port 182 nsew signal input
rlabel metal3 s 0 180480 800 180600 6 data_arrays_0_0_ext_ram_rdata2[30]
port 183 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 data_arrays_0_0_ext_ram_rdata2[31]
port 184 nsew signal input
rlabel metal3 s 0 181840 800 181960 6 data_arrays_0_0_ext_ram_rdata2[32]
port 185 nsew signal input
rlabel metal3 s 0 182656 800 182776 6 data_arrays_0_0_ext_ram_rdata2[33]
port 186 nsew signal input
rlabel metal3 s 0 183336 800 183456 6 data_arrays_0_0_ext_ram_rdata2[34]
port 187 nsew signal input
rlabel metal3 s 0 184016 800 184136 6 data_arrays_0_0_ext_ram_rdata2[35]
port 188 nsew signal input
rlabel metal3 s 0 184696 800 184816 6 data_arrays_0_0_ext_ram_rdata2[36]
port 189 nsew signal input
rlabel metal3 s 0 185376 800 185496 6 data_arrays_0_0_ext_ram_rdata2[37]
port 190 nsew signal input
rlabel metal3 s 0 186192 800 186312 6 data_arrays_0_0_ext_ram_rdata2[38]
port 191 nsew signal input
rlabel metal3 s 0 186872 800 186992 6 data_arrays_0_0_ext_ram_rdata2[39]
port 192 nsew signal input
rlabel metal3 s 0 161440 800 161560 6 data_arrays_0_0_ext_ram_rdata2[3]
port 193 nsew signal input
rlabel metal3 s 0 187552 800 187672 6 data_arrays_0_0_ext_ram_rdata2[40]
port 194 nsew signal input
rlabel metal3 s 0 188232 800 188352 6 data_arrays_0_0_ext_ram_rdata2[41]
port 195 nsew signal input
rlabel metal3 s 0 188912 800 189032 6 data_arrays_0_0_ext_ram_rdata2[42]
port 196 nsew signal input
rlabel metal3 s 0 189592 800 189712 6 data_arrays_0_0_ext_ram_rdata2[43]
port 197 nsew signal input
rlabel metal3 s 0 190408 800 190528 6 data_arrays_0_0_ext_ram_rdata2[44]
port 198 nsew signal input
rlabel metal3 s 0 191088 800 191208 6 data_arrays_0_0_ext_ram_rdata2[45]
port 199 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 data_arrays_0_0_ext_ram_rdata2[46]
port 200 nsew signal input
rlabel metal3 s 0 192448 800 192568 6 data_arrays_0_0_ext_ram_rdata2[47]
port 201 nsew signal input
rlabel metal3 s 0 193128 800 193248 6 data_arrays_0_0_ext_ram_rdata2[48]
port 202 nsew signal input
rlabel metal3 s 0 193944 800 194064 6 data_arrays_0_0_ext_ram_rdata2[49]
port 203 nsew signal input
rlabel metal3 s 0 162120 800 162240 6 data_arrays_0_0_ext_ram_rdata2[4]
port 204 nsew signal input
rlabel metal3 s 0 194624 800 194744 6 data_arrays_0_0_ext_ram_rdata2[50]
port 205 nsew signal input
rlabel metal3 s 0 195304 800 195424 6 data_arrays_0_0_ext_ram_rdata2[51]
port 206 nsew signal input
rlabel metal3 s 0 195984 800 196104 6 data_arrays_0_0_ext_ram_rdata2[52]
port 207 nsew signal input
rlabel metal3 s 0 196664 800 196784 6 data_arrays_0_0_ext_ram_rdata2[53]
port 208 nsew signal input
rlabel metal3 s 0 197344 800 197464 6 data_arrays_0_0_ext_ram_rdata2[54]
port 209 nsew signal input
rlabel metal3 s 0 198160 800 198280 6 data_arrays_0_0_ext_ram_rdata2[55]
port 210 nsew signal input
rlabel metal3 s 0 198840 800 198960 6 data_arrays_0_0_ext_ram_rdata2[56]
port 211 nsew signal input
rlabel metal3 s 0 199520 800 199640 6 data_arrays_0_0_ext_ram_rdata2[57]
port 212 nsew signal input
rlabel metal3 s 0 200200 800 200320 6 data_arrays_0_0_ext_ram_rdata2[58]
port 213 nsew signal input
rlabel metal3 s 0 200880 800 201000 6 data_arrays_0_0_ext_ram_rdata2[59]
port 214 nsew signal input
rlabel metal3 s 0 162936 800 163056 6 data_arrays_0_0_ext_ram_rdata2[5]
port 215 nsew signal input
rlabel metal3 s 0 201560 800 201680 6 data_arrays_0_0_ext_ram_rdata2[60]
port 216 nsew signal input
rlabel metal3 s 0 202376 800 202496 6 data_arrays_0_0_ext_ram_rdata2[61]
port 217 nsew signal input
rlabel metal3 s 0 203056 800 203176 6 data_arrays_0_0_ext_ram_rdata2[62]
port 218 nsew signal input
rlabel metal3 s 0 203736 800 203856 6 data_arrays_0_0_ext_ram_rdata2[63]
port 219 nsew signal input
rlabel metal3 s 0 163616 800 163736 6 data_arrays_0_0_ext_ram_rdata2[6]
port 220 nsew signal input
rlabel metal3 s 0 164296 800 164416 6 data_arrays_0_0_ext_ram_rdata2[7]
port 221 nsew signal input
rlabel metal3 s 0 164976 800 165096 6 data_arrays_0_0_ext_ram_rdata2[8]
port 222 nsew signal input
rlabel metal3 s 0 165656 800 165776 6 data_arrays_0_0_ext_ram_rdata2[9]
port 223 nsew signal input
rlabel metal3 s 0 204416 800 204536 6 data_arrays_0_0_ext_ram_rdata3[0]
port 224 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 data_arrays_0_0_ext_ram_rdata3[10]
port 225 nsew signal input
rlabel metal3 s 0 212168 800 212288 6 data_arrays_0_0_ext_ram_rdata3[11]
port 226 nsew signal input
rlabel metal3 s 0 212848 800 212968 6 data_arrays_0_0_ext_ram_rdata3[12]
port 227 nsew signal input
rlabel metal3 s 0 213664 800 213784 6 data_arrays_0_0_ext_ram_rdata3[13]
port 228 nsew signal input
rlabel metal3 s 0 214344 800 214464 6 data_arrays_0_0_ext_ram_rdata3[14]
port 229 nsew signal input
rlabel metal3 s 0 215024 800 215144 6 data_arrays_0_0_ext_ram_rdata3[15]
port 230 nsew signal input
rlabel metal3 s 0 215704 800 215824 6 data_arrays_0_0_ext_ram_rdata3[16]
port 231 nsew signal input
rlabel metal3 s 0 216384 800 216504 6 data_arrays_0_0_ext_ram_rdata3[17]
port 232 nsew signal input
rlabel metal3 s 0 217064 800 217184 6 data_arrays_0_0_ext_ram_rdata3[18]
port 233 nsew signal input
rlabel metal3 s 0 217880 800 218000 6 data_arrays_0_0_ext_ram_rdata3[19]
port 234 nsew signal input
rlabel metal3 s 0 205096 800 205216 6 data_arrays_0_0_ext_ram_rdata3[1]
port 235 nsew signal input
rlabel metal3 s 0 218560 800 218680 6 data_arrays_0_0_ext_ram_rdata3[20]
port 236 nsew signal input
rlabel metal3 s 0 219240 800 219360 6 data_arrays_0_0_ext_ram_rdata3[21]
port 237 nsew signal input
rlabel metal3 s 0 219920 800 220040 6 data_arrays_0_0_ext_ram_rdata3[22]
port 238 nsew signal input
rlabel metal3 s 0 220600 800 220720 6 data_arrays_0_0_ext_ram_rdata3[23]
port 239 nsew signal input
rlabel metal3 s 0 221280 800 221400 6 data_arrays_0_0_ext_ram_rdata3[24]
port 240 nsew signal input
rlabel metal3 s 0 222096 800 222216 6 data_arrays_0_0_ext_ram_rdata3[25]
port 241 nsew signal input
rlabel metal3 s 0 222776 800 222896 6 data_arrays_0_0_ext_ram_rdata3[26]
port 242 nsew signal input
rlabel metal3 s 0 223456 800 223576 6 data_arrays_0_0_ext_ram_rdata3[27]
port 243 nsew signal input
rlabel metal3 s 0 224136 800 224256 6 data_arrays_0_0_ext_ram_rdata3[28]
port 244 nsew signal input
rlabel metal3 s 0 224816 800 224936 6 data_arrays_0_0_ext_ram_rdata3[29]
port 245 nsew signal input
rlabel metal3 s 0 205912 800 206032 6 data_arrays_0_0_ext_ram_rdata3[2]
port 246 nsew signal input
rlabel metal3 s 0 225632 800 225752 6 data_arrays_0_0_ext_ram_rdata3[30]
port 247 nsew signal input
rlabel metal3 s 0 226312 800 226432 6 data_arrays_0_0_ext_ram_rdata3[31]
port 248 nsew signal input
rlabel metal3 s 0 226992 800 227112 6 data_arrays_0_0_ext_ram_rdata3[32]
port 249 nsew signal input
rlabel metal3 s 0 227672 800 227792 6 data_arrays_0_0_ext_ram_rdata3[33]
port 250 nsew signal input
rlabel metal3 s 0 228352 800 228472 6 data_arrays_0_0_ext_ram_rdata3[34]
port 251 nsew signal input
rlabel metal3 s 0 229032 800 229152 6 data_arrays_0_0_ext_ram_rdata3[35]
port 252 nsew signal input
rlabel metal3 s 0 229848 800 229968 6 data_arrays_0_0_ext_ram_rdata3[36]
port 253 nsew signal input
rlabel metal3 s 0 230528 800 230648 6 data_arrays_0_0_ext_ram_rdata3[37]
port 254 nsew signal input
rlabel metal3 s 0 231208 800 231328 6 data_arrays_0_0_ext_ram_rdata3[38]
port 255 nsew signal input
rlabel metal3 s 0 231888 800 232008 6 data_arrays_0_0_ext_ram_rdata3[39]
port 256 nsew signal input
rlabel metal3 s 0 206592 800 206712 6 data_arrays_0_0_ext_ram_rdata3[3]
port 257 nsew signal input
rlabel metal3 s 0 232568 800 232688 6 data_arrays_0_0_ext_ram_rdata3[40]
port 258 nsew signal input
rlabel metal3 s 0 233248 800 233368 6 data_arrays_0_0_ext_ram_rdata3[41]
port 259 nsew signal input
rlabel metal3 s 0 234064 800 234184 6 data_arrays_0_0_ext_ram_rdata3[42]
port 260 nsew signal input
rlabel metal3 s 0 234744 800 234864 6 data_arrays_0_0_ext_ram_rdata3[43]
port 261 nsew signal input
rlabel metal3 s 0 235424 800 235544 6 data_arrays_0_0_ext_ram_rdata3[44]
port 262 nsew signal input
rlabel metal3 s 0 236104 800 236224 6 data_arrays_0_0_ext_ram_rdata3[45]
port 263 nsew signal input
rlabel metal3 s 0 236784 800 236904 6 data_arrays_0_0_ext_ram_rdata3[46]
port 264 nsew signal input
rlabel metal3 s 0 237600 800 237720 6 data_arrays_0_0_ext_ram_rdata3[47]
port 265 nsew signal input
rlabel metal3 s 0 238280 800 238400 6 data_arrays_0_0_ext_ram_rdata3[48]
port 266 nsew signal input
rlabel metal3 s 0 238960 800 239080 6 data_arrays_0_0_ext_ram_rdata3[49]
port 267 nsew signal input
rlabel metal3 s 0 207272 800 207392 6 data_arrays_0_0_ext_ram_rdata3[4]
port 268 nsew signal input
rlabel metal3 s 0 239640 800 239760 6 data_arrays_0_0_ext_ram_rdata3[50]
port 269 nsew signal input
rlabel metal3 s 0 240320 800 240440 6 data_arrays_0_0_ext_ram_rdata3[51]
port 270 nsew signal input
rlabel metal3 s 0 241000 800 241120 6 data_arrays_0_0_ext_ram_rdata3[52]
port 271 nsew signal input
rlabel metal3 s 0 241816 800 241936 6 data_arrays_0_0_ext_ram_rdata3[53]
port 272 nsew signal input
rlabel metal3 s 0 242496 800 242616 6 data_arrays_0_0_ext_ram_rdata3[54]
port 273 nsew signal input
rlabel metal3 s 0 243176 800 243296 6 data_arrays_0_0_ext_ram_rdata3[55]
port 274 nsew signal input
rlabel metal3 s 0 243856 800 243976 6 data_arrays_0_0_ext_ram_rdata3[56]
port 275 nsew signal input
rlabel metal3 s 0 244536 800 244656 6 data_arrays_0_0_ext_ram_rdata3[57]
port 276 nsew signal input
rlabel metal3 s 0 245352 800 245472 6 data_arrays_0_0_ext_ram_rdata3[58]
port 277 nsew signal input
rlabel metal3 s 0 246032 800 246152 6 data_arrays_0_0_ext_ram_rdata3[59]
port 278 nsew signal input
rlabel metal3 s 0 207952 800 208072 6 data_arrays_0_0_ext_ram_rdata3[5]
port 279 nsew signal input
rlabel metal3 s 0 246712 800 246832 6 data_arrays_0_0_ext_ram_rdata3[60]
port 280 nsew signal input
rlabel metal3 s 0 247392 800 247512 6 data_arrays_0_0_ext_ram_rdata3[61]
port 281 nsew signal input
rlabel metal3 s 0 248072 800 248192 6 data_arrays_0_0_ext_ram_rdata3[62]
port 282 nsew signal input
rlabel metal3 s 0 248752 800 248872 6 data_arrays_0_0_ext_ram_rdata3[63]
port 283 nsew signal input
rlabel metal3 s 0 208632 800 208752 6 data_arrays_0_0_ext_ram_rdata3[6]
port 284 nsew signal input
rlabel metal3 s 0 209312 800 209432 6 data_arrays_0_0_ext_ram_rdata3[7]
port 285 nsew signal input
rlabel metal3 s 0 210128 800 210248 6 data_arrays_0_0_ext_ram_rdata3[8]
port 286 nsew signal input
rlabel metal3 s 0 210808 800 210928 6 data_arrays_0_0_ext_ram_rdata3[9]
port 287 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 data_arrays_0_0_ext_ram_wdata[0]
port 288 nsew signal output
rlabel metal3 s 0 104456 800 104576 6 data_arrays_0_0_ext_ram_wdata[10]
port 289 nsew signal output
rlabel metal3 s 0 105136 800 105256 6 data_arrays_0_0_ext_ram_wdata[11]
port 290 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 data_arrays_0_0_ext_ram_wdata[12]
port 291 nsew signal output
rlabel metal3 s 0 106496 800 106616 6 data_arrays_0_0_ext_ram_wdata[13]
port 292 nsew signal output
rlabel metal3 s 0 107312 800 107432 6 data_arrays_0_0_ext_ram_wdata[14]
port 293 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 data_arrays_0_0_ext_ram_wdata[15]
port 294 nsew signal output
rlabel metal3 s 0 108672 800 108792 6 data_arrays_0_0_ext_ram_wdata[16]
port 295 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 data_arrays_0_0_ext_ram_wdata[17]
port 296 nsew signal output
rlabel metal3 s 0 110032 800 110152 6 data_arrays_0_0_ext_ram_wdata[18]
port 297 nsew signal output
rlabel metal3 s 0 110712 800 110832 6 data_arrays_0_0_ext_ram_wdata[19]
port 298 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 data_arrays_0_0_ext_ram_wdata[1]
port 299 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 data_arrays_0_0_ext_ram_wdata[20]
port 300 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 data_arrays_0_0_ext_ram_wdata[21]
port 301 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 data_arrays_0_0_ext_ram_wdata[22]
port 302 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 data_arrays_0_0_ext_ram_wdata[23]
port 303 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 data_arrays_0_0_ext_ram_wdata[24]
port 304 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 data_arrays_0_0_ext_ram_wdata[25]
port 305 nsew signal output
rlabel metal3 s 0 115744 800 115864 6 data_arrays_0_0_ext_ram_wdata[26]
port 306 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 data_arrays_0_0_ext_ram_wdata[27]
port 307 nsew signal output
rlabel metal3 s 0 117104 800 117224 6 data_arrays_0_0_ext_ram_wdata[28]
port 308 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 data_arrays_0_0_ext_ram_wdata[29]
port 309 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 data_arrays_0_0_ext_ram_wdata[2]
port 310 nsew signal output
rlabel metal3 s 0 118464 800 118584 6 data_arrays_0_0_ext_ram_wdata[30]
port 311 nsew signal output
rlabel metal3 s 0 119280 800 119400 6 data_arrays_0_0_ext_ram_wdata[31]
port 312 nsew signal output
rlabel metal3 s 0 119960 800 120080 6 data_arrays_0_0_ext_ram_wdata[32]
port 313 nsew signal output
rlabel metal3 s 0 120640 800 120760 6 data_arrays_0_0_ext_ram_wdata[33]
port 314 nsew signal output
rlabel metal3 s 0 121320 800 121440 6 data_arrays_0_0_ext_ram_wdata[34]
port 315 nsew signal output
rlabel metal3 s 0 122000 800 122120 6 data_arrays_0_0_ext_ram_wdata[35]
port 316 nsew signal output
rlabel metal3 s 0 122816 800 122936 6 data_arrays_0_0_ext_ram_wdata[36]
port 317 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 data_arrays_0_0_ext_ram_wdata[37]
port 318 nsew signal output
rlabel metal3 s 0 124176 800 124296 6 data_arrays_0_0_ext_ram_wdata[38]
port 319 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 data_arrays_0_0_ext_ram_wdata[39]
port 320 nsew signal output
rlabel metal3 s 0 99560 800 99680 6 data_arrays_0_0_ext_ram_wdata[3]
port 321 nsew signal output
rlabel metal3 s 0 125536 800 125656 6 data_arrays_0_0_ext_ram_wdata[40]
port 322 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 data_arrays_0_0_ext_ram_wdata[41]
port 323 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 data_arrays_0_0_ext_ram_wdata[42]
port 324 nsew signal output
rlabel metal3 s 0 127712 800 127832 6 data_arrays_0_0_ext_ram_wdata[43]
port 325 nsew signal output
rlabel metal3 s 0 128392 800 128512 6 data_arrays_0_0_ext_ram_wdata[44]
port 326 nsew signal output
rlabel metal3 s 0 129072 800 129192 6 data_arrays_0_0_ext_ram_wdata[45]
port 327 nsew signal output
rlabel metal3 s 0 129752 800 129872 6 data_arrays_0_0_ext_ram_wdata[46]
port 328 nsew signal output
rlabel metal3 s 0 130432 800 130552 6 data_arrays_0_0_ext_ram_wdata[47]
port 329 nsew signal output
rlabel metal3 s 0 131248 800 131368 6 data_arrays_0_0_ext_ram_wdata[48]
port 330 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 data_arrays_0_0_ext_ram_wdata[49]
port 331 nsew signal output
rlabel metal3 s 0 100240 800 100360 6 data_arrays_0_0_ext_ram_wdata[4]
port 332 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 data_arrays_0_0_ext_ram_wdata[50]
port 333 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 data_arrays_0_0_ext_ram_wdata[51]
port 334 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 data_arrays_0_0_ext_ram_wdata[52]
port 335 nsew signal output
rlabel metal3 s 0 134784 800 134904 6 data_arrays_0_0_ext_ram_wdata[53]
port 336 nsew signal output
rlabel metal3 s 0 135464 800 135584 6 data_arrays_0_0_ext_ram_wdata[54]
port 337 nsew signal output
rlabel metal3 s 0 136144 800 136264 6 data_arrays_0_0_ext_ram_wdata[55]
port 338 nsew signal output
rlabel metal3 s 0 136824 800 136944 6 data_arrays_0_0_ext_ram_wdata[56]
port 339 nsew signal output
rlabel metal3 s 0 137504 800 137624 6 data_arrays_0_0_ext_ram_wdata[57]
port 340 nsew signal output
rlabel metal3 s 0 138184 800 138304 6 data_arrays_0_0_ext_ram_wdata[58]
port 341 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 data_arrays_0_0_ext_ram_wdata[59]
port 342 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 data_arrays_0_0_ext_ram_wdata[5]
port 343 nsew signal output
rlabel metal3 s 0 139680 800 139800 6 data_arrays_0_0_ext_ram_wdata[60]
port 344 nsew signal output
rlabel metal3 s 0 140360 800 140480 6 data_arrays_0_0_ext_ram_wdata[61]
port 345 nsew signal output
rlabel metal3 s 0 141040 800 141160 6 data_arrays_0_0_ext_ram_wdata[62]
port 346 nsew signal output
rlabel metal3 s 0 141720 800 141840 6 data_arrays_0_0_ext_ram_wdata[63]
port 347 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 data_arrays_0_0_ext_ram_wdata[6]
port 348 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 data_arrays_0_0_ext_ram_wdata[7]
port 349 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 data_arrays_0_0_ext_ram_wdata[8]
port 350 nsew signal output
rlabel metal3 s 0 103776 800 103896 6 data_arrays_0_0_ext_ram_wdata[9]
port 351 nsew signal output
rlabel metal3 s 0 146752 800 146872 6 data_arrays_0_0_ext_ram_web
port 352 nsew signal output
rlabel metal3 s 0 142536 800 142656 6 data_arrays_0_0_ext_ram_wmask[0]
port 353 nsew signal output
rlabel metal3 s 0 143216 800 143336 6 data_arrays_0_0_ext_ram_wmask[1]
port 354 nsew signal output
rlabel metal3 s 352679 340416 353479 340536 6 data_arrays_0_ext_ram_addr1[0]
port 355 nsew signal output
rlabel metal3 s 352679 342184 353479 342304 6 data_arrays_0_ext_ram_addr1[1]
port 356 nsew signal output
rlabel metal3 s 352679 343952 353479 344072 6 data_arrays_0_ext_ram_addr1[2]
port 357 nsew signal output
rlabel metal3 s 352679 345720 353479 345840 6 data_arrays_0_ext_ram_addr1[3]
port 358 nsew signal output
rlabel metal3 s 352679 347488 353479 347608 6 data_arrays_0_ext_ram_addr1[4]
port 359 nsew signal output
rlabel metal3 s 352679 349256 353479 349376 6 data_arrays_0_ext_ram_addr1[5]
port 360 nsew signal output
rlabel metal3 s 352679 351024 353479 351144 6 data_arrays_0_ext_ram_addr1[6]
port 361 nsew signal output
rlabel metal3 s 352679 352792 353479 352912 6 data_arrays_0_ext_ram_addr1[7]
port 362 nsew signal output
rlabel metal3 s 352679 354560 353479 354680 6 data_arrays_0_ext_ram_addr1[8]
port 363 nsew signal output
rlabel metal3 s 352679 228352 353479 228472 6 data_arrays_0_ext_ram_addr[0]
port 364 nsew signal output
rlabel metal3 s 352679 230120 353479 230240 6 data_arrays_0_ext_ram_addr[1]
port 365 nsew signal output
rlabel metal3 s 352679 231888 353479 232008 6 data_arrays_0_ext_ram_addr[2]
port 366 nsew signal output
rlabel metal3 s 352679 233656 353479 233776 6 data_arrays_0_ext_ram_addr[3]
port 367 nsew signal output
rlabel metal3 s 352679 235424 353479 235544 6 data_arrays_0_ext_ram_addr[4]
port 368 nsew signal output
rlabel metal3 s 352679 237192 353479 237312 6 data_arrays_0_ext_ram_addr[5]
port 369 nsew signal output
rlabel metal3 s 352679 239096 353479 239216 6 data_arrays_0_ext_ram_addr[6]
port 370 nsew signal output
rlabel metal3 s 352679 240864 353479 240984 6 data_arrays_0_ext_ram_addr[7]
port 371 nsew signal output
rlabel metal3 s 352679 242632 353479 242752 6 data_arrays_0_ext_ram_addr[8]
port 372 nsew signal output
rlabel metal3 s 352679 244400 353479 244520 6 data_arrays_0_ext_ram_clk
port 373 nsew signal output
rlabel metal3 s 352679 326136 353479 326256 6 data_arrays_0_ext_ram_csb1[0]
port 374 nsew signal output
rlabel metal3 s 352679 327904 353479 328024 6 data_arrays_0_ext_ram_csb1[1]
port 375 nsew signal output
rlabel metal3 s 352679 329672 353479 329792 6 data_arrays_0_ext_ram_csb1[2]
port 376 nsew signal output
rlabel metal3 s 352679 331440 353479 331560 6 data_arrays_0_ext_ram_csb1[3]
port 377 nsew signal output
rlabel metal3 s 352679 333344 353479 333464 6 data_arrays_0_ext_ram_csb1[4]
port 378 nsew signal output
rlabel metal3 s 352679 335112 353479 335232 6 data_arrays_0_ext_ram_csb1[5]
port 379 nsew signal output
rlabel metal3 s 352679 336880 353479 337000 6 data_arrays_0_ext_ram_csb1[6]
port 380 nsew signal output
rlabel metal3 s 352679 338648 353479 338768 6 data_arrays_0_ext_ram_csb1[7]
port 381 nsew signal output
rlabel metal3 s 352679 310224 353479 310344 6 data_arrays_0_ext_ram_csb[0]
port 382 nsew signal output
rlabel metal3 s 352679 311992 353479 312112 6 data_arrays_0_ext_ram_csb[1]
port 383 nsew signal output
rlabel metal3 s 352679 313760 353479 313880 6 data_arrays_0_ext_ram_csb[2]
port 384 nsew signal output
rlabel metal3 s 352679 315528 353479 315648 6 data_arrays_0_ext_ram_csb[3]
port 385 nsew signal output
rlabel metal3 s 352679 317296 353479 317416 6 data_arrays_0_ext_ram_csb[4]
port 386 nsew signal output
rlabel metal3 s 352679 319064 353479 319184 6 data_arrays_0_ext_ram_csb[5]
port 387 nsew signal output
rlabel metal3 s 352679 320832 353479 320952 6 data_arrays_0_ext_ram_csb[6]
port 388 nsew signal output
rlabel metal3 s 352679 322600 353479 322720 6 data_arrays_0_ext_ram_csb[7]
port 389 nsew signal output
rlabel metal3 s 352679 824 353479 944 6 data_arrays_0_ext_ram_rdata0[0]
port 390 nsew signal input
rlabel metal3 s 352679 18504 353479 18624 6 data_arrays_0_ext_ram_rdata0[10]
port 391 nsew signal input
rlabel metal3 s 352679 20272 353479 20392 6 data_arrays_0_ext_ram_rdata0[11]
port 392 nsew signal input
rlabel metal3 s 352679 22040 353479 22160 6 data_arrays_0_ext_ram_rdata0[12]
port 393 nsew signal input
rlabel metal3 s 352679 23808 353479 23928 6 data_arrays_0_ext_ram_rdata0[13]
port 394 nsew signal input
rlabel metal3 s 352679 25712 353479 25832 6 data_arrays_0_ext_ram_rdata0[14]
port 395 nsew signal input
rlabel metal3 s 352679 27480 353479 27600 6 data_arrays_0_ext_ram_rdata0[15]
port 396 nsew signal input
rlabel metal3 s 352679 29248 353479 29368 6 data_arrays_0_ext_ram_rdata0[16]
port 397 nsew signal input
rlabel metal3 s 352679 31016 353479 31136 6 data_arrays_0_ext_ram_rdata0[17]
port 398 nsew signal input
rlabel metal3 s 352679 32784 353479 32904 6 data_arrays_0_ext_ram_rdata0[18]
port 399 nsew signal input
rlabel metal3 s 352679 34552 353479 34672 6 data_arrays_0_ext_ram_rdata0[19]
port 400 nsew signal input
rlabel metal3 s 352679 2592 353479 2712 6 data_arrays_0_ext_ram_rdata0[1]
port 401 nsew signal input
rlabel metal3 s 352679 36320 353479 36440 6 data_arrays_0_ext_ram_rdata0[20]
port 402 nsew signal input
rlabel metal3 s 352679 38088 353479 38208 6 data_arrays_0_ext_ram_rdata0[21]
port 403 nsew signal input
rlabel metal3 s 352679 39856 353479 39976 6 data_arrays_0_ext_ram_rdata0[22]
port 404 nsew signal input
rlabel metal3 s 352679 41624 353479 41744 6 data_arrays_0_ext_ram_rdata0[23]
port 405 nsew signal input
rlabel metal3 s 352679 43392 353479 43512 6 data_arrays_0_ext_ram_rdata0[24]
port 406 nsew signal input
rlabel metal3 s 352679 45160 353479 45280 6 data_arrays_0_ext_ram_rdata0[25]
port 407 nsew signal input
rlabel metal3 s 352679 46928 353479 47048 6 data_arrays_0_ext_ram_rdata0[26]
port 408 nsew signal input
rlabel metal3 s 352679 48832 353479 48952 6 data_arrays_0_ext_ram_rdata0[27]
port 409 nsew signal input
rlabel metal3 s 352679 50600 353479 50720 6 data_arrays_0_ext_ram_rdata0[28]
port 410 nsew signal input
rlabel metal3 s 352679 52368 353479 52488 6 data_arrays_0_ext_ram_rdata0[29]
port 411 nsew signal input
rlabel metal3 s 352679 4360 353479 4480 6 data_arrays_0_ext_ram_rdata0[2]
port 412 nsew signal input
rlabel metal3 s 352679 54136 353479 54256 6 data_arrays_0_ext_ram_rdata0[30]
port 413 nsew signal input
rlabel metal3 s 352679 55904 353479 56024 6 data_arrays_0_ext_ram_rdata0[31]
port 414 nsew signal input
rlabel metal3 s 352679 6128 353479 6248 6 data_arrays_0_ext_ram_rdata0[3]
port 415 nsew signal input
rlabel metal3 s 352679 7896 353479 8016 6 data_arrays_0_ext_ram_rdata0[4]
port 416 nsew signal input
rlabel metal3 s 352679 9664 353479 9784 6 data_arrays_0_ext_ram_rdata0[5]
port 417 nsew signal input
rlabel metal3 s 352679 11432 353479 11552 6 data_arrays_0_ext_ram_rdata0[6]
port 418 nsew signal input
rlabel metal3 s 352679 13200 353479 13320 6 data_arrays_0_ext_ram_rdata0[7]
port 419 nsew signal input
rlabel metal3 s 352679 14968 353479 15088 6 data_arrays_0_ext_ram_rdata0[8]
port 420 nsew signal input
rlabel metal3 s 352679 16736 353479 16856 6 data_arrays_0_ext_ram_rdata0[9]
port 421 nsew signal input
rlabel metal3 s 352679 57672 353479 57792 6 data_arrays_0_ext_ram_rdata1[0]
port 422 nsew signal input
rlabel metal3 s 352679 75488 353479 75608 6 data_arrays_0_ext_ram_rdata1[10]
port 423 nsew signal input
rlabel metal3 s 352679 77256 353479 77376 6 data_arrays_0_ext_ram_rdata1[11]
port 424 nsew signal input
rlabel metal3 s 352679 79024 353479 79144 6 data_arrays_0_ext_ram_rdata1[12]
port 425 nsew signal input
rlabel metal3 s 352679 80792 353479 80912 6 data_arrays_0_ext_ram_rdata1[13]
port 426 nsew signal input
rlabel metal3 s 352679 82560 353479 82680 6 data_arrays_0_ext_ram_rdata1[14]
port 427 nsew signal input
rlabel metal3 s 352679 84328 353479 84448 6 data_arrays_0_ext_ram_rdata1[15]
port 428 nsew signal input
rlabel metal3 s 352679 86096 353479 86216 6 data_arrays_0_ext_ram_rdata1[16]
port 429 nsew signal input
rlabel metal3 s 352679 87864 353479 87984 6 data_arrays_0_ext_ram_rdata1[17]
port 430 nsew signal input
rlabel metal3 s 352679 89632 353479 89752 6 data_arrays_0_ext_ram_rdata1[18]
port 431 nsew signal input
rlabel metal3 s 352679 91400 353479 91520 6 data_arrays_0_ext_ram_rdata1[19]
port 432 nsew signal input
rlabel metal3 s 352679 59440 353479 59560 6 data_arrays_0_ext_ram_rdata1[1]
port 433 nsew signal input
rlabel metal3 s 352679 93168 353479 93288 6 data_arrays_0_ext_ram_rdata1[20]
port 434 nsew signal input
rlabel metal3 s 352679 94936 353479 95056 6 data_arrays_0_ext_ram_rdata1[21]
port 435 nsew signal input
rlabel metal3 s 352679 96840 353479 96960 6 data_arrays_0_ext_ram_rdata1[22]
port 436 nsew signal input
rlabel metal3 s 352679 98608 353479 98728 6 data_arrays_0_ext_ram_rdata1[23]
port 437 nsew signal input
rlabel metal3 s 352679 100376 353479 100496 6 data_arrays_0_ext_ram_rdata1[24]
port 438 nsew signal input
rlabel metal3 s 352679 102144 353479 102264 6 data_arrays_0_ext_ram_rdata1[25]
port 439 nsew signal input
rlabel metal3 s 352679 103912 353479 104032 6 data_arrays_0_ext_ram_rdata1[26]
port 440 nsew signal input
rlabel metal3 s 352679 105680 353479 105800 6 data_arrays_0_ext_ram_rdata1[27]
port 441 nsew signal input
rlabel metal3 s 352679 107448 353479 107568 6 data_arrays_0_ext_ram_rdata1[28]
port 442 nsew signal input
rlabel metal3 s 352679 109216 353479 109336 6 data_arrays_0_ext_ram_rdata1[29]
port 443 nsew signal input
rlabel metal3 s 352679 61208 353479 61328 6 data_arrays_0_ext_ram_rdata1[2]
port 444 nsew signal input
rlabel metal3 s 352679 110984 353479 111104 6 data_arrays_0_ext_ram_rdata1[30]
port 445 nsew signal input
rlabel metal3 s 352679 112752 353479 112872 6 data_arrays_0_ext_ram_rdata1[31]
port 446 nsew signal input
rlabel metal3 s 352679 62976 353479 63096 6 data_arrays_0_ext_ram_rdata1[3]
port 447 nsew signal input
rlabel metal3 s 352679 64744 353479 64864 6 data_arrays_0_ext_ram_rdata1[4]
port 448 nsew signal input
rlabel metal3 s 352679 66512 353479 66632 6 data_arrays_0_ext_ram_rdata1[5]
port 449 nsew signal input
rlabel metal3 s 352679 68280 353479 68400 6 data_arrays_0_ext_ram_rdata1[6]
port 450 nsew signal input
rlabel metal3 s 352679 70048 353479 70168 6 data_arrays_0_ext_ram_rdata1[7]
port 451 nsew signal input
rlabel metal3 s 352679 71952 353479 72072 6 data_arrays_0_ext_ram_rdata1[8]
port 452 nsew signal input
rlabel metal3 s 352679 73720 353479 73840 6 data_arrays_0_ext_ram_rdata1[9]
port 453 nsew signal input
rlabel metal3 s 352679 114520 353479 114640 6 data_arrays_0_ext_ram_rdata2[0]
port 454 nsew signal input
rlabel metal3 s 352679 132336 353479 132456 6 data_arrays_0_ext_ram_rdata2[10]
port 455 nsew signal input
rlabel metal3 s 352679 134104 353479 134224 6 data_arrays_0_ext_ram_rdata2[11]
port 456 nsew signal input
rlabel metal3 s 352679 135872 353479 135992 6 data_arrays_0_ext_ram_rdata2[12]
port 457 nsew signal input
rlabel metal3 s 352679 137640 353479 137760 6 data_arrays_0_ext_ram_rdata2[13]
port 458 nsew signal input
rlabel metal3 s 352679 139408 353479 139528 6 data_arrays_0_ext_ram_rdata2[14]
port 459 nsew signal input
rlabel metal3 s 352679 141176 353479 141296 6 data_arrays_0_ext_ram_rdata2[15]
port 460 nsew signal input
rlabel metal3 s 352679 143080 353479 143200 6 data_arrays_0_ext_ram_rdata2[16]
port 461 nsew signal input
rlabel metal3 s 352679 144848 353479 144968 6 data_arrays_0_ext_ram_rdata2[17]
port 462 nsew signal input
rlabel metal3 s 352679 146616 353479 146736 6 data_arrays_0_ext_ram_rdata2[18]
port 463 nsew signal input
rlabel metal3 s 352679 148384 353479 148504 6 data_arrays_0_ext_ram_rdata2[19]
port 464 nsew signal input
rlabel metal3 s 352679 116288 353479 116408 6 data_arrays_0_ext_ram_rdata2[1]
port 465 nsew signal input
rlabel metal3 s 352679 150152 353479 150272 6 data_arrays_0_ext_ram_rdata2[20]
port 466 nsew signal input
rlabel metal3 s 352679 151920 353479 152040 6 data_arrays_0_ext_ram_rdata2[21]
port 467 nsew signal input
rlabel metal3 s 352679 153688 353479 153808 6 data_arrays_0_ext_ram_rdata2[22]
port 468 nsew signal input
rlabel metal3 s 352679 155456 353479 155576 6 data_arrays_0_ext_ram_rdata2[23]
port 469 nsew signal input
rlabel metal3 s 352679 157224 353479 157344 6 data_arrays_0_ext_ram_rdata2[24]
port 470 nsew signal input
rlabel metal3 s 352679 158992 353479 159112 6 data_arrays_0_ext_ram_rdata2[25]
port 471 nsew signal input
rlabel metal3 s 352679 160760 353479 160880 6 data_arrays_0_ext_ram_rdata2[26]
port 472 nsew signal input
rlabel metal3 s 352679 162528 353479 162648 6 data_arrays_0_ext_ram_rdata2[27]
port 473 nsew signal input
rlabel metal3 s 352679 164296 353479 164416 6 data_arrays_0_ext_ram_rdata2[28]
port 474 nsew signal input
rlabel metal3 s 352679 166064 353479 166184 6 data_arrays_0_ext_ram_rdata2[29]
port 475 nsew signal input
rlabel metal3 s 352679 118056 353479 118176 6 data_arrays_0_ext_ram_rdata2[2]
port 476 nsew signal input
rlabel metal3 s 352679 167968 353479 168088 6 data_arrays_0_ext_ram_rdata2[30]
port 477 nsew signal input
rlabel metal3 s 352679 169736 353479 169856 6 data_arrays_0_ext_ram_rdata2[31]
port 478 nsew signal input
rlabel metal3 s 352679 119960 353479 120080 6 data_arrays_0_ext_ram_rdata2[3]
port 479 nsew signal input
rlabel metal3 s 352679 121728 353479 121848 6 data_arrays_0_ext_ram_rdata2[4]
port 480 nsew signal input
rlabel metal3 s 352679 123496 353479 123616 6 data_arrays_0_ext_ram_rdata2[5]
port 481 nsew signal input
rlabel metal3 s 352679 125264 353479 125384 6 data_arrays_0_ext_ram_rdata2[6]
port 482 nsew signal input
rlabel metal3 s 352679 127032 353479 127152 6 data_arrays_0_ext_ram_rdata2[7]
port 483 nsew signal input
rlabel metal3 s 352679 128800 353479 128920 6 data_arrays_0_ext_ram_rdata2[8]
port 484 nsew signal input
rlabel metal3 s 352679 130568 353479 130688 6 data_arrays_0_ext_ram_rdata2[9]
port 485 nsew signal input
rlabel metal3 s 352679 171504 353479 171624 6 data_arrays_0_ext_ram_rdata3[0]
port 486 nsew signal input
rlabel metal3 s 352679 189184 353479 189304 6 data_arrays_0_ext_ram_rdata3[10]
port 487 nsew signal input
rlabel metal3 s 352679 191088 353479 191208 6 data_arrays_0_ext_ram_rdata3[11]
port 488 nsew signal input
rlabel metal3 s 352679 192856 353479 192976 6 data_arrays_0_ext_ram_rdata3[12]
port 489 nsew signal input
rlabel metal3 s 352679 194624 353479 194744 6 data_arrays_0_ext_ram_rdata3[13]
port 490 nsew signal input
rlabel metal3 s 352679 196392 353479 196512 6 data_arrays_0_ext_ram_rdata3[14]
port 491 nsew signal input
rlabel metal3 s 352679 198160 353479 198280 6 data_arrays_0_ext_ram_rdata3[15]
port 492 nsew signal input
rlabel metal3 s 352679 199928 353479 200048 6 data_arrays_0_ext_ram_rdata3[16]
port 493 nsew signal input
rlabel metal3 s 352679 201696 353479 201816 6 data_arrays_0_ext_ram_rdata3[17]
port 494 nsew signal input
rlabel metal3 s 352679 203464 353479 203584 6 data_arrays_0_ext_ram_rdata3[18]
port 495 nsew signal input
rlabel metal3 s 352679 205232 353479 205352 6 data_arrays_0_ext_ram_rdata3[19]
port 496 nsew signal input
rlabel metal3 s 352679 173272 353479 173392 6 data_arrays_0_ext_ram_rdata3[1]
port 497 nsew signal input
rlabel metal3 s 352679 207000 353479 207120 6 data_arrays_0_ext_ram_rdata3[20]
port 498 nsew signal input
rlabel metal3 s 352679 208768 353479 208888 6 data_arrays_0_ext_ram_rdata3[21]
port 499 nsew signal input
rlabel metal3 s 352679 210536 353479 210656 6 data_arrays_0_ext_ram_rdata3[22]
port 500 nsew signal input
rlabel metal3 s 352679 212304 353479 212424 6 data_arrays_0_ext_ram_rdata3[23]
port 501 nsew signal input
rlabel metal3 s 352679 214208 353479 214328 6 data_arrays_0_ext_ram_rdata3[24]
port 502 nsew signal input
rlabel metal3 s 352679 215976 353479 216096 6 data_arrays_0_ext_ram_rdata3[25]
port 503 nsew signal input
rlabel metal3 s 352679 217744 353479 217864 6 data_arrays_0_ext_ram_rdata3[26]
port 504 nsew signal input
rlabel metal3 s 352679 219512 353479 219632 6 data_arrays_0_ext_ram_rdata3[27]
port 505 nsew signal input
rlabel metal3 s 352679 221280 353479 221400 6 data_arrays_0_ext_ram_rdata3[28]
port 506 nsew signal input
rlabel metal3 s 352679 223048 353479 223168 6 data_arrays_0_ext_ram_rdata3[29]
port 507 nsew signal input
rlabel metal3 s 352679 175040 353479 175160 6 data_arrays_0_ext_ram_rdata3[2]
port 508 nsew signal input
rlabel metal3 s 352679 224816 353479 224936 6 data_arrays_0_ext_ram_rdata3[30]
port 509 nsew signal input
rlabel metal3 s 352679 226584 353479 226704 6 data_arrays_0_ext_ram_rdata3[31]
port 510 nsew signal input
rlabel metal3 s 352679 176808 353479 176928 6 data_arrays_0_ext_ram_rdata3[3]
port 511 nsew signal input
rlabel metal3 s 352679 178576 353479 178696 6 data_arrays_0_ext_ram_rdata3[4]
port 512 nsew signal input
rlabel metal3 s 352679 180344 353479 180464 6 data_arrays_0_ext_ram_rdata3[5]
port 513 nsew signal input
rlabel metal3 s 352679 182112 353479 182232 6 data_arrays_0_ext_ram_rdata3[6]
port 514 nsew signal input
rlabel metal3 s 352679 183880 353479 184000 6 data_arrays_0_ext_ram_rdata3[7]
port 515 nsew signal input
rlabel metal3 s 352679 185648 353479 185768 6 data_arrays_0_ext_ram_rdata3[8]
port 516 nsew signal input
rlabel metal3 s 352679 187416 353479 187536 6 data_arrays_0_ext_ram_rdata3[9]
port 517 nsew signal input
rlabel metal3 s 352679 246168 353479 246288 6 data_arrays_0_ext_ram_wdata[0]
port 518 nsew signal output
rlabel metal3 s 352679 263984 353479 264104 6 data_arrays_0_ext_ram_wdata[10]
port 519 nsew signal output
rlabel metal3 s 352679 265752 353479 265872 6 data_arrays_0_ext_ram_wdata[11]
port 520 nsew signal output
rlabel metal3 s 352679 267520 353479 267640 6 data_arrays_0_ext_ram_wdata[12]
port 521 nsew signal output
rlabel metal3 s 352679 269288 353479 269408 6 data_arrays_0_ext_ram_wdata[13]
port 522 nsew signal output
rlabel metal3 s 352679 271056 353479 271176 6 data_arrays_0_ext_ram_wdata[14]
port 523 nsew signal output
rlabel metal3 s 352679 272824 353479 272944 6 data_arrays_0_ext_ram_wdata[15]
port 524 nsew signal output
rlabel metal3 s 352679 274592 353479 274712 6 data_arrays_0_ext_ram_wdata[16]
port 525 nsew signal output
rlabel metal3 s 352679 276360 353479 276480 6 data_arrays_0_ext_ram_wdata[17]
port 526 nsew signal output
rlabel metal3 s 352679 278128 353479 278248 6 data_arrays_0_ext_ram_wdata[18]
port 527 nsew signal output
rlabel metal3 s 352679 279896 353479 280016 6 data_arrays_0_ext_ram_wdata[19]
port 528 nsew signal output
rlabel metal3 s 352679 247936 353479 248056 6 data_arrays_0_ext_ram_wdata[1]
port 529 nsew signal output
rlabel metal3 s 352679 281664 353479 281784 6 data_arrays_0_ext_ram_wdata[20]
port 530 nsew signal output
rlabel metal3 s 352679 283432 353479 283552 6 data_arrays_0_ext_ram_wdata[21]
port 531 nsew signal output
rlabel metal3 s 352679 285336 353479 285456 6 data_arrays_0_ext_ram_wdata[22]
port 532 nsew signal output
rlabel metal3 s 352679 287104 353479 287224 6 data_arrays_0_ext_ram_wdata[23]
port 533 nsew signal output
rlabel metal3 s 352679 288872 353479 288992 6 data_arrays_0_ext_ram_wdata[24]
port 534 nsew signal output
rlabel metal3 s 352679 290640 353479 290760 6 data_arrays_0_ext_ram_wdata[25]
port 535 nsew signal output
rlabel metal3 s 352679 292408 353479 292528 6 data_arrays_0_ext_ram_wdata[26]
port 536 nsew signal output
rlabel metal3 s 352679 294176 353479 294296 6 data_arrays_0_ext_ram_wdata[27]
port 537 nsew signal output
rlabel metal3 s 352679 295944 353479 296064 6 data_arrays_0_ext_ram_wdata[28]
port 538 nsew signal output
rlabel metal3 s 352679 297712 353479 297832 6 data_arrays_0_ext_ram_wdata[29]
port 539 nsew signal output
rlabel metal3 s 352679 249704 353479 249824 6 data_arrays_0_ext_ram_wdata[2]
port 540 nsew signal output
rlabel metal3 s 352679 299480 353479 299600 6 data_arrays_0_ext_ram_wdata[30]
port 541 nsew signal output
rlabel metal3 s 352679 301248 353479 301368 6 data_arrays_0_ext_ram_wdata[31]
port 542 nsew signal output
rlabel metal3 s 352679 251472 353479 251592 6 data_arrays_0_ext_ram_wdata[3]
port 543 nsew signal output
rlabel metal3 s 352679 253240 353479 253360 6 data_arrays_0_ext_ram_wdata[4]
port 544 nsew signal output
rlabel metal3 s 352679 255008 353479 255128 6 data_arrays_0_ext_ram_wdata[5]
port 545 nsew signal output
rlabel metal3 s 352679 256776 353479 256896 6 data_arrays_0_ext_ram_wdata[6]
port 546 nsew signal output
rlabel metal3 s 352679 258544 353479 258664 6 data_arrays_0_ext_ram_wdata[7]
port 547 nsew signal output
rlabel metal3 s 352679 260312 353479 260432 6 data_arrays_0_ext_ram_wdata[8]
port 548 nsew signal output
rlabel metal3 s 352679 262216 353479 262336 6 data_arrays_0_ext_ram_wdata[9]
port 549 nsew signal output
rlabel metal3 s 352679 324368 353479 324488 6 data_arrays_0_ext_ram_web
port 550 nsew signal output
rlabel metal3 s 352679 303016 353479 303136 6 data_arrays_0_ext_ram_wmask[0]
port 551 nsew signal output
rlabel metal3 s 352679 304784 353479 304904 6 data_arrays_0_ext_ram_wmask[1]
port 552 nsew signal output
rlabel metal3 s 352679 306552 353479 306672 6 data_arrays_0_ext_ram_wmask[2]
port 553 nsew signal output
rlabel metal3 s 352679 308320 353479 308440 6 data_arrays_0_ext_ram_wmask[3]
port 554 nsew signal output
rlabel metal2 s 1490 354823 1546 355623 6 io_in[0]
port 555 nsew signal input
rlabel metal2 s 94502 354823 94558 355623 6 io_in[10]
port 556 nsew signal input
rlabel metal2 s 103794 354823 103850 355623 6 io_in[11]
port 557 nsew signal input
rlabel metal2 s 113086 354823 113142 355623 6 io_in[12]
port 558 nsew signal input
rlabel metal2 s 122378 354823 122434 355623 6 io_in[13]
port 559 nsew signal input
rlabel metal2 s 131670 354823 131726 355623 6 io_in[14]
port 560 nsew signal input
rlabel metal2 s 140962 354823 141018 355623 6 io_in[15]
port 561 nsew signal input
rlabel metal2 s 150254 354823 150310 355623 6 io_in[16]
port 562 nsew signal input
rlabel metal2 s 159546 354823 159602 355623 6 io_in[17]
port 563 nsew signal input
rlabel metal2 s 168838 354823 168894 355623 6 io_in[18]
port 564 nsew signal input
rlabel metal2 s 178222 354823 178278 355623 6 io_in[19]
port 565 nsew signal input
rlabel metal2 s 10782 354823 10838 355623 6 io_in[1]
port 566 nsew signal input
rlabel metal2 s 187514 354823 187570 355623 6 io_in[20]
port 567 nsew signal input
rlabel metal2 s 196806 354823 196862 355623 6 io_in[21]
port 568 nsew signal input
rlabel metal2 s 206098 354823 206154 355623 6 io_in[22]
port 569 nsew signal input
rlabel metal2 s 215390 354823 215446 355623 6 io_in[23]
port 570 nsew signal input
rlabel metal2 s 224682 354823 224738 355623 6 io_in[24]
port 571 nsew signal input
rlabel metal2 s 233974 354823 234030 355623 6 io_in[25]
port 572 nsew signal input
rlabel metal2 s 243266 354823 243322 355623 6 io_in[26]
port 573 nsew signal input
rlabel metal2 s 252558 354823 252614 355623 6 io_in[27]
port 574 nsew signal input
rlabel metal2 s 261850 354823 261906 355623 6 io_in[28]
port 575 nsew signal input
rlabel metal2 s 271234 354823 271290 355623 6 io_in[29]
port 576 nsew signal input
rlabel metal2 s 20074 354823 20130 355623 6 io_in[2]
port 577 nsew signal input
rlabel metal2 s 280526 354823 280582 355623 6 io_in[30]
port 578 nsew signal input
rlabel metal2 s 289818 354823 289874 355623 6 io_in[31]
port 579 nsew signal input
rlabel metal2 s 299110 354823 299166 355623 6 io_in[32]
port 580 nsew signal input
rlabel metal2 s 308402 354823 308458 355623 6 io_in[33]
port 581 nsew signal input
rlabel metal2 s 317694 354823 317750 355623 6 io_in[34]
port 582 nsew signal input
rlabel metal2 s 326986 354823 327042 355623 6 io_in[35]
port 583 nsew signal input
rlabel metal2 s 336278 354823 336334 355623 6 io_in[36]
port 584 nsew signal input
rlabel metal2 s 345570 354823 345626 355623 6 io_in[37]
port 585 nsew signal input
rlabel metal2 s 29366 354823 29422 355623 6 io_in[3]
port 586 nsew signal input
rlabel metal2 s 38658 354823 38714 355623 6 io_in[4]
port 587 nsew signal input
rlabel metal2 s 47950 354823 48006 355623 6 io_in[5]
port 588 nsew signal input
rlabel metal2 s 57242 354823 57298 355623 6 io_in[6]
port 589 nsew signal input
rlabel metal2 s 66534 354823 66590 355623 6 io_in[7]
port 590 nsew signal input
rlabel metal2 s 75826 354823 75882 355623 6 io_in[8]
port 591 nsew signal input
rlabel metal2 s 85118 354823 85174 355623 6 io_in[9]
port 592 nsew signal input
rlabel metal2 s 4526 354823 4582 355623 6 io_oeb[0]
port 593 nsew signal output
rlabel metal2 s 97538 354823 97594 355623 6 io_oeb[10]
port 594 nsew signal output
rlabel metal2 s 106830 354823 106886 355623 6 io_oeb[11]
port 595 nsew signal output
rlabel metal2 s 116122 354823 116178 355623 6 io_oeb[12]
port 596 nsew signal output
rlabel metal2 s 125506 354823 125562 355623 6 io_oeb[13]
port 597 nsew signal output
rlabel metal2 s 134798 354823 134854 355623 6 io_oeb[14]
port 598 nsew signal output
rlabel metal2 s 144090 354823 144146 355623 6 io_oeb[15]
port 599 nsew signal output
rlabel metal2 s 153382 354823 153438 355623 6 io_oeb[16]
port 600 nsew signal output
rlabel metal2 s 162674 354823 162730 355623 6 io_oeb[17]
port 601 nsew signal output
rlabel metal2 s 171966 354823 172022 355623 6 io_oeb[18]
port 602 nsew signal output
rlabel metal2 s 181258 354823 181314 355623 6 io_oeb[19]
port 603 nsew signal output
rlabel metal2 s 13818 354823 13874 355623 6 io_oeb[1]
port 604 nsew signal output
rlabel metal2 s 190550 354823 190606 355623 6 io_oeb[20]
port 605 nsew signal output
rlabel metal2 s 199842 354823 199898 355623 6 io_oeb[21]
port 606 nsew signal output
rlabel metal2 s 209226 354823 209282 355623 6 io_oeb[22]
port 607 nsew signal output
rlabel metal2 s 218518 354823 218574 355623 6 io_oeb[23]
port 608 nsew signal output
rlabel metal2 s 227810 354823 227866 355623 6 io_oeb[24]
port 609 nsew signal output
rlabel metal2 s 237102 354823 237158 355623 6 io_oeb[25]
port 610 nsew signal output
rlabel metal2 s 246394 354823 246450 355623 6 io_oeb[26]
port 611 nsew signal output
rlabel metal2 s 255686 354823 255742 355623 6 io_oeb[27]
port 612 nsew signal output
rlabel metal2 s 264978 354823 265034 355623 6 io_oeb[28]
port 613 nsew signal output
rlabel metal2 s 274270 354823 274326 355623 6 io_oeb[29]
port 614 nsew signal output
rlabel metal2 s 23110 354823 23166 355623 6 io_oeb[2]
port 615 nsew signal output
rlabel metal2 s 283562 354823 283618 355623 6 io_oeb[30]
port 616 nsew signal output
rlabel metal2 s 292854 354823 292910 355623 6 io_oeb[31]
port 617 nsew signal output
rlabel metal2 s 302238 354823 302294 355623 6 io_oeb[32]
port 618 nsew signal output
rlabel metal2 s 311530 354823 311586 355623 6 io_oeb[33]
port 619 nsew signal output
rlabel metal2 s 320822 354823 320878 355623 6 io_oeb[34]
port 620 nsew signal output
rlabel metal2 s 330114 354823 330170 355623 6 io_oeb[35]
port 621 nsew signal output
rlabel metal2 s 339406 354823 339462 355623 6 io_oeb[36]
port 622 nsew signal output
rlabel metal2 s 348698 354823 348754 355623 6 io_oeb[37]
port 623 nsew signal output
rlabel metal2 s 32494 354823 32550 355623 6 io_oeb[3]
port 624 nsew signal output
rlabel metal2 s 41786 354823 41842 355623 6 io_oeb[4]
port 625 nsew signal output
rlabel metal2 s 51078 354823 51134 355623 6 io_oeb[5]
port 626 nsew signal output
rlabel metal2 s 60370 354823 60426 355623 6 io_oeb[6]
port 627 nsew signal output
rlabel metal2 s 69662 354823 69718 355623 6 io_oeb[7]
port 628 nsew signal output
rlabel metal2 s 78954 354823 79010 355623 6 io_oeb[8]
port 629 nsew signal output
rlabel metal2 s 88246 354823 88302 355623 6 io_oeb[9]
port 630 nsew signal output
rlabel metal2 s 7654 354823 7710 355623 6 io_out[0]
port 631 nsew signal output
rlabel metal2 s 100666 354823 100722 355623 6 io_out[10]
port 632 nsew signal output
rlabel metal2 s 109958 354823 110014 355623 6 io_out[11]
port 633 nsew signal output
rlabel metal2 s 119250 354823 119306 355623 6 io_out[12]
port 634 nsew signal output
rlabel metal2 s 128542 354823 128598 355623 6 io_out[13]
port 635 nsew signal output
rlabel metal2 s 137834 354823 137890 355623 6 io_out[14]
port 636 nsew signal output
rlabel metal2 s 147126 354823 147182 355623 6 io_out[15]
port 637 nsew signal output
rlabel metal2 s 156510 354823 156566 355623 6 io_out[16]
port 638 nsew signal output
rlabel metal2 s 165802 354823 165858 355623 6 io_out[17]
port 639 nsew signal output
rlabel metal2 s 175094 354823 175150 355623 6 io_out[18]
port 640 nsew signal output
rlabel metal2 s 184386 354823 184442 355623 6 io_out[19]
port 641 nsew signal output
rlabel metal2 s 16946 354823 17002 355623 6 io_out[1]
port 642 nsew signal output
rlabel metal2 s 193678 354823 193734 355623 6 io_out[20]
port 643 nsew signal output
rlabel metal2 s 202970 354823 203026 355623 6 io_out[21]
port 644 nsew signal output
rlabel metal2 s 212262 354823 212318 355623 6 io_out[22]
port 645 nsew signal output
rlabel metal2 s 221554 354823 221610 355623 6 io_out[23]
port 646 nsew signal output
rlabel metal2 s 230846 354823 230902 355623 6 io_out[24]
port 647 nsew signal output
rlabel metal2 s 240230 354823 240286 355623 6 io_out[25]
port 648 nsew signal output
rlabel metal2 s 249522 354823 249578 355623 6 io_out[26]
port 649 nsew signal output
rlabel metal2 s 258814 354823 258870 355623 6 io_out[27]
port 650 nsew signal output
rlabel metal2 s 268106 354823 268162 355623 6 io_out[28]
port 651 nsew signal output
rlabel metal2 s 277398 354823 277454 355623 6 io_out[29]
port 652 nsew signal output
rlabel metal2 s 26238 354823 26294 355623 6 io_out[2]
port 653 nsew signal output
rlabel metal2 s 286690 354823 286746 355623 6 io_out[30]
port 654 nsew signal output
rlabel metal2 s 295982 354823 296038 355623 6 io_out[31]
port 655 nsew signal output
rlabel metal2 s 305274 354823 305330 355623 6 io_out[32]
port 656 nsew signal output
rlabel metal2 s 314566 354823 314622 355623 6 io_out[33]
port 657 nsew signal output
rlabel metal2 s 323858 354823 323914 355623 6 io_out[34]
port 658 nsew signal output
rlabel metal2 s 333242 354823 333298 355623 6 io_out[35]
port 659 nsew signal output
rlabel metal2 s 342534 354823 342590 355623 6 io_out[36]
port 660 nsew signal output
rlabel metal2 s 351826 354823 351882 355623 6 io_out[37]
port 661 nsew signal output
rlabel metal2 s 35530 354823 35586 355623 6 io_out[3]
port 662 nsew signal output
rlabel metal2 s 44822 354823 44878 355623 6 io_out[4]
port 663 nsew signal output
rlabel metal2 s 54114 354823 54170 355623 6 io_out[5]
port 664 nsew signal output
rlabel metal2 s 63498 354823 63554 355623 6 io_out[6]
port 665 nsew signal output
rlabel metal2 s 72790 354823 72846 355623 6 io_out[7]
port 666 nsew signal output
rlabel metal2 s 82082 354823 82138 355623 6 io_out[8]
port 667 nsew signal output
rlabel metal2 s 91374 354823 91430 355623 6 io_out[9]
port 668 nsew signal output
rlabel metal2 s 351550 0 351606 800 6 irq[0]
port 669 nsew signal output
rlabel metal2 s 352286 0 352342 800 6 irq[1]
port 670 nsew signal output
rlabel metal2 s 353022 0 353078 800 6 irq[2]
port 671 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 la_data_in[0]
port 672 nsew signal input
rlabel metal2 s 291382 0 291438 800 6 la_data_in[100]
port 673 nsew signal input
rlabel metal2 s 293498 0 293554 800 6 la_data_in[101]
port 674 nsew signal input
rlabel metal2 s 295614 0 295670 800 6 la_data_in[102]
port 675 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_data_in[103]
port 676 nsew signal input
rlabel metal2 s 299938 0 299994 800 6 la_data_in[104]
port 677 nsew signal input
rlabel metal2 s 302054 0 302110 800 6 la_data_in[105]
port 678 nsew signal input
rlabel metal2 s 304262 0 304318 800 6 la_data_in[106]
port 679 nsew signal input
rlabel metal2 s 306378 0 306434 800 6 la_data_in[107]
port 680 nsew signal input
rlabel metal2 s 308586 0 308642 800 6 la_data_in[108]
port 681 nsew signal input
rlabel metal2 s 310702 0 310758 800 6 la_data_in[109]
port 682 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[10]
port 683 nsew signal input
rlabel metal2 s 312818 0 312874 800 6 la_data_in[110]
port 684 nsew signal input
rlabel metal2 s 315026 0 315082 800 6 la_data_in[111]
port 685 nsew signal input
rlabel metal2 s 317142 0 317198 800 6 la_data_in[112]
port 686 nsew signal input
rlabel metal2 s 319258 0 319314 800 6 la_data_in[113]
port 687 nsew signal input
rlabel metal2 s 321466 0 321522 800 6 la_data_in[114]
port 688 nsew signal input
rlabel metal2 s 323582 0 323638 800 6 la_data_in[115]
port 689 nsew signal input
rlabel metal2 s 325790 0 325846 800 6 la_data_in[116]
port 690 nsew signal input
rlabel metal2 s 327906 0 327962 800 6 la_data_in[117]
port 691 nsew signal input
rlabel metal2 s 330022 0 330078 800 6 la_data_in[118]
port 692 nsew signal input
rlabel metal2 s 332230 0 332286 800 6 la_data_in[119]
port 693 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[11]
port 694 nsew signal input
rlabel metal2 s 334346 0 334402 800 6 la_data_in[120]
port 695 nsew signal input
rlabel metal2 s 336462 0 336518 800 6 la_data_in[121]
port 696 nsew signal input
rlabel metal2 s 338670 0 338726 800 6 la_data_in[122]
port 697 nsew signal input
rlabel metal2 s 340786 0 340842 800 6 la_data_in[123]
port 698 nsew signal input
rlabel metal2 s 342994 0 343050 800 6 la_data_in[124]
port 699 nsew signal input
rlabel metal2 s 345110 0 345166 800 6 la_data_in[125]
port 700 nsew signal input
rlabel metal2 s 347226 0 347282 800 6 la_data_in[126]
port 701 nsew signal input
rlabel metal2 s 349434 0 349490 800 6 la_data_in[127]
port 702 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[12]
port 703 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[13]
port 704 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_data_in[14]
port 705 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[15]
port 706 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[16]
port 707 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[17]
port 708 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[18]
port 709 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[19]
port 710 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[1]
port 711 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[20]
port 712 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[21]
port 713 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_data_in[22]
port 714 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_data_in[23]
port 715 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_data_in[24]
port 716 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[25]
port 717 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_data_in[26]
port 718 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[27]
port 719 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_data_in[28]
port 720 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_data_in[29]
port 721 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[2]
port 722 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[30]
port 723 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_data_in[31]
port 724 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[32]
port 725 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_data_in[33]
port 726 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[34]
port 727 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_data_in[35]
port 728 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[36]
port 729 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_data_in[37]
port 730 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[38]
port 731 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 la_data_in[39]
port 732 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[3]
port 733 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_data_in[40]
port 734 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_data_in[41]
port 735 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_data_in[42]
port 736 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[43]
port 737 nsew signal input
rlabel metal2 s 170862 0 170918 800 6 la_data_in[44]
port 738 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 la_data_in[45]
port 739 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[46]
port 740 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_data_in[47]
port 741 nsew signal input
rlabel metal2 s 179510 0 179566 800 6 la_data_in[48]
port 742 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 la_data_in[49]
port 743 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[4]
port 744 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_data_in[50]
port 745 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_data_in[51]
port 746 nsew signal input
rlabel metal2 s 188066 0 188122 800 6 la_data_in[52]
port 747 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[53]
port 748 nsew signal input
rlabel metal2 s 192390 0 192446 800 6 la_data_in[54]
port 749 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_data_in[55]
port 750 nsew signal input
rlabel metal2 s 196714 0 196770 800 6 la_data_in[56]
port 751 nsew signal input
rlabel metal2 s 198830 0 198886 800 6 la_data_in[57]
port 752 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_data_in[58]
port 753 nsew signal input
rlabel metal2 s 203154 0 203210 800 6 la_data_in[59]
port 754 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[5]
port 755 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_data_in[60]
port 756 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_data_in[61]
port 757 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_data_in[62]
port 758 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_data_in[63]
port 759 nsew signal input
rlabel metal2 s 213918 0 213974 800 6 la_data_in[64]
port 760 nsew signal input
rlabel metal2 s 216034 0 216090 800 6 la_data_in[65]
port 761 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_data_in[66]
port 762 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_data_in[67]
port 763 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_data_in[68]
port 764 nsew signal input
rlabel metal2 s 224682 0 224738 800 6 la_data_in[69]
port 765 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[6]
port 766 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_data_in[70]
port 767 nsew signal input
rlabel metal2 s 229006 0 229062 800 6 la_data_in[71]
port 768 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_data_in[72]
port 769 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_data_in[73]
port 770 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_data_in[74]
port 771 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_data_in[75]
port 772 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_data_in[76]
port 773 nsew signal input
rlabel metal2 s 241886 0 241942 800 6 la_data_in[77]
port 774 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 la_data_in[78]
port 775 nsew signal input
rlabel metal2 s 246210 0 246266 800 6 la_data_in[79]
port 776 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_data_in[7]
port 777 nsew signal input
rlabel metal2 s 248326 0 248382 800 6 la_data_in[80]
port 778 nsew signal input
rlabel metal2 s 250442 0 250498 800 6 la_data_in[81]
port 779 nsew signal input
rlabel metal2 s 252650 0 252706 800 6 la_data_in[82]
port 780 nsew signal input
rlabel metal2 s 254766 0 254822 800 6 la_data_in[83]
port 781 nsew signal input
rlabel metal2 s 256882 0 256938 800 6 la_data_in[84]
port 782 nsew signal input
rlabel metal2 s 259090 0 259146 800 6 la_data_in[85]
port 783 nsew signal input
rlabel metal2 s 261206 0 261262 800 6 la_data_in[86]
port 784 nsew signal input
rlabel metal2 s 263414 0 263470 800 6 la_data_in[87]
port 785 nsew signal input
rlabel metal2 s 265530 0 265586 800 6 la_data_in[88]
port 786 nsew signal input
rlabel metal2 s 267646 0 267702 800 6 la_data_in[89]
port 787 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[8]
port 788 nsew signal input
rlabel metal2 s 269854 0 269910 800 6 la_data_in[90]
port 789 nsew signal input
rlabel metal2 s 271970 0 272026 800 6 la_data_in[91]
port 790 nsew signal input
rlabel metal2 s 274086 0 274142 800 6 la_data_in[92]
port 791 nsew signal input
rlabel metal2 s 276294 0 276350 800 6 la_data_in[93]
port 792 nsew signal input
rlabel metal2 s 278410 0 278466 800 6 la_data_in[94]
port 793 nsew signal input
rlabel metal2 s 280618 0 280674 800 6 la_data_in[95]
port 794 nsew signal input
rlabel metal2 s 282734 0 282790 800 6 la_data_in[96]
port 795 nsew signal input
rlabel metal2 s 284850 0 284906 800 6 la_data_in[97]
port 796 nsew signal input
rlabel metal2 s 287058 0 287114 800 6 la_data_in[98]
port 797 nsew signal input
rlabel metal2 s 289174 0 289230 800 6 la_data_in[99]
port 798 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[9]
port 799 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_out[0]
port 800 nsew signal output
rlabel metal2 s 292026 0 292082 800 6 la_data_out[100]
port 801 nsew signal output
rlabel metal2 s 294234 0 294290 800 6 la_data_out[101]
port 802 nsew signal output
rlabel metal2 s 296350 0 296406 800 6 la_data_out[102]
port 803 nsew signal output
rlabel metal2 s 298466 0 298522 800 6 la_data_out[103]
port 804 nsew signal output
rlabel metal2 s 300674 0 300730 800 6 la_data_out[104]
port 805 nsew signal output
rlabel metal2 s 302790 0 302846 800 6 la_data_out[105]
port 806 nsew signal output
rlabel metal2 s 304998 0 305054 800 6 la_data_out[106]
port 807 nsew signal output
rlabel metal2 s 307114 0 307170 800 6 la_data_out[107]
port 808 nsew signal output
rlabel metal2 s 309230 0 309286 800 6 la_data_out[108]
port 809 nsew signal output
rlabel metal2 s 311438 0 311494 800 6 la_data_out[109]
port 810 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[10]
port 811 nsew signal output
rlabel metal2 s 313554 0 313610 800 6 la_data_out[110]
port 812 nsew signal output
rlabel metal2 s 315670 0 315726 800 6 la_data_out[111]
port 813 nsew signal output
rlabel metal2 s 317878 0 317934 800 6 la_data_out[112]
port 814 nsew signal output
rlabel metal2 s 319994 0 320050 800 6 la_data_out[113]
port 815 nsew signal output
rlabel metal2 s 322202 0 322258 800 6 la_data_out[114]
port 816 nsew signal output
rlabel metal2 s 324318 0 324374 800 6 la_data_out[115]
port 817 nsew signal output
rlabel metal2 s 326434 0 326490 800 6 la_data_out[116]
port 818 nsew signal output
rlabel metal2 s 328642 0 328698 800 6 la_data_out[117]
port 819 nsew signal output
rlabel metal2 s 330758 0 330814 800 6 la_data_out[118]
port 820 nsew signal output
rlabel metal2 s 332966 0 333022 800 6 la_data_out[119]
port 821 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[11]
port 822 nsew signal output
rlabel metal2 s 335082 0 335138 800 6 la_data_out[120]
port 823 nsew signal output
rlabel metal2 s 337198 0 337254 800 6 la_data_out[121]
port 824 nsew signal output
rlabel metal2 s 339406 0 339462 800 6 la_data_out[122]
port 825 nsew signal output
rlabel metal2 s 341522 0 341578 800 6 la_data_out[123]
port 826 nsew signal output
rlabel metal2 s 343638 0 343694 800 6 la_data_out[124]
port 827 nsew signal output
rlabel metal2 s 345846 0 345902 800 6 la_data_out[125]
port 828 nsew signal output
rlabel metal2 s 347962 0 348018 800 6 la_data_out[126]
port 829 nsew signal output
rlabel metal2 s 350170 0 350226 800 6 la_data_out[127]
port 830 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[12]
port 831 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[13]
port 832 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[14]
port 833 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[15]
port 834 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 la_data_out[16]
port 835 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 la_data_out[17]
port 836 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 la_data_out[18]
port 837 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[19]
port 838 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[1]
port 839 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 la_data_out[20]
port 840 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[21]
port 841 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 la_data_out[22]
port 842 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[23]
port 843 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 la_data_out[24]
port 844 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[25]
port 845 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[26]
port 846 nsew signal output
rlabel metal2 s 135074 0 135130 800 6 la_data_out[27]
port 847 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[28]
port 848 nsew signal output
rlabel metal2 s 139306 0 139362 800 6 la_data_out[29]
port 849 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[2]
port 850 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[30]
port 851 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[31]
port 852 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[32]
port 853 nsew signal output
rlabel metal2 s 147954 0 148010 800 6 la_data_out[33]
port 854 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[34]
port 855 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[35]
port 856 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[36]
port 857 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[37]
port 858 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 la_data_out[38]
port 859 nsew signal output
rlabel metal2 s 160834 0 160890 800 6 la_data_out[39]
port 860 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[3]
port 861 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 la_data_out[40]
port 862 nsew signal output
rlabel metal2 s 165158 0 165214 800 6 la_data_out[41]
port 863 nsew signal output
rlabel metal2 s 167274 0 167330 800 6 la_data_out[42]
port 864 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[43]
port 865 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 la_data_out[44]
port 866 nsew signal output
rlabel metal2 s 173714 0 173770 800 6 la_data_out[45]
port 867 nsew signal output
rlabel metal2 s 175922 0 175978 800 6 la_data_out[46]
port 868 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 la_data_out[47]
port 869 nsew signal output
rlabel metal2 s 180246 0 180302 800 6 la_data_out[48]
port 870 nsew signal output
rlabel metal2 s 182362 0 182418 800 6 la_data_out[49]
port 871 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[4]
port 872 nsew signal output
rlabel metal2 s 184478 0 184534 800 6 la_data_out[50]
port 873 nsew signal output
rlabel metal2 s 186686 0 186742 800 6 la_data_out[51]
port 874 nsew signal output
rlabel metal2 s 188802 0 188858 800 6 la_data_out[52]
port 875 nsew signal output
rlabel metal2 s 190918 0 190974 800 6 la_data_out[53]
port 876 nsew signal output
rlabel metal2 s 193126 0 193182 800 6 la_data_out[54]
port 877 nsew signal output
rlabel metal2 s 195242 0 195298 800 6 la_data_out[55]
port 878 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 la_data_out[56]
port 879 nsew signal output
rlabel metal2 s 199566 0 199622 800 6 la_data_out[57]
port 880 nsew signal output
rlabel metal2 s 201682 0 201738 800 6 la_data_out[58]
port 881 nsew signal output
rlabel metal2 s 203890 0 203946 800 6 la_data_out[59]
port 882 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[5]
port 883 nsew signal output
rlabel metal2 s 206006 0 206062 800 6 la_data_out[60]
port 884 nsew signal output
rlabel metal2 s 208214 0 208270 800 6 la_data_out[61]
port 885 nsew signal output
rlabel metal2 s 210330 0 210386 800 6 la_data_out[62]
port 886 nsew signal output
rlabel metal2 s 212446 0 212502 800 6 la_data_out[63]
port 887 nsew signal output
rlabel metal2 s 214654 0 214710 800 6 la_data_out[64]
port 888 nsew signal output
rlabel metal2 s 216770 0 216826 800 6 la_data_out[65]
port 889 nsew signal output
rlabel metal2 s 218886 0 218942 800 6 la_data_out[66]
port 890 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 la_data_out[67]
port 891 nsew signal output
rlabel metal2 s 223210 0 223266 800 6 la_data_out[68]
port 892 nsew signal output
rlabel metal2 s 225418 0 225474 800 6 la_data_out[69]
port 893 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[6]
port 894 nsew signal output
rlabel metal2 s 227534 0 227590 800 6 la_data_out[70]
port 895 nsew signal output
rlabel metal2 s 229650 0 229706 800 6 la_data_out[71]
port 896 nsew signal output
rlabel metal2 s 231858 0 231914 800 6 la_data_out[72]
port 897 nsew signal output
rlabel metal2 s 233974 0 234030 800 6 la_data_out[73]
port 898 nsew signal output
rlabel metal2 s 236090 0 236146 800 6 la_data_out[74]
port 899 nsew signal output
rlabel metal2 s 238298 0 238354 800 6 la_data_out[75]
port 900 nsew signal output
rlabel metal2 s 240414 0 240470 800 6 la_data_out[76]
port 901 nsew signal output
rlabel metal2 s 242622 0 242678 800 6 la_data_out[77]
port 902 nsew signal output
rlabel metal2 s 244738 0 244794 800 6 la_data_out[78]
port 903 nsew signal output
rlabel metal2 s 246854 0 246910 800 6 la_data_out[79]
port 904 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[7]
port 905 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 la_data_out[80]
port 906 nsew signal output
rlabel metal2 s 251178 0 251234 800 6 la_data_out[81]
port 907 nsew signal output
rlabel metal2 s 253294 0 253350 800 6 la_data_out[82]
port 908 nsew signal output
rlabel metal2 s 255502 0 255558 800 6 la_data_out[83]
port 909 nsew signal output
rlabel metal2 s 257618 0 257674 800 6 la_data_out[84]
port 910 nsew signal output
rlabel metal2 s 259826 0 259882 800 6 la_data_out[85]
port 911 nsew signal output
rlabel metal2 s 261942 0 261998 800 6 la_data_out[86]
port 912 nsew signal output
rlabel metal2 s 264058 0 264114 800 6 la_data_out[87]
port 913 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[88]
port 914 nsew signal output
rlabel metal2 s 268382 0 268438 800 6 la_data_out[89]
port 915 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 la_data_out[8]
port 916 nsew signal output
rlabel metal2 s 270590 0 270646 800 6 la_data_out[90]
port 917 nsew signal output
rlabel metal2 s 272706 0 272762 800 6 la_data_out[91]
port 918 nsew signal output
rlabel metal2 s 274822 0 274878 800 6 la_data_out[92]
port 919 nsew signal output
rlabel metal2 s 277030 0 277086 800 6 la_data_out[93]
port 920 nsew signal output
rlabel metal2 s 279146 0 279202 800 6 la_data_out[94]
port 921 nsew signal output
rlabel metal2 s 281262 0 281318 800 6 la_data_out[95]
port 922 nsew signal output
rlabel metal2 s 283470 0 283526 800 6 la_data_out[96]
port 923 nsew signal output
rlabel metal2 s 285586 0 285642 800 6 la_data_out[97]
port 924 nsew signal output
rlabel metal2 s 287794 0 287850 800 6 la_data_out[98]
port 925 nsew signal output
rlabel metal2 s 289910 0 289966 800 6 la_data_out[99]
port 926 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[9]
port 927 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_oenb[0]
port 928 nsew signal input
rlabel metal2 s 292762 0 292818 800 6 la_oenb[100]
port 929 nsew signal input
rlabel metal2 s 294878 0 294934 800 6 la_oenb[101]
port 930 nsew signal input
rlabel metal2 s 297086 0 297142 800 6 la_oenb[102]
port 931 nsew signal input
rlabel metal2 s 299202 0 299258 800 6 la_oenb[103]
port 932 nsew signal input
rlabel metal2 s 301410 0 301466 800 6 la_oenb[104]
port 933 nsew signal input
rlabel metal2 s 303526 0 303582 800 6 la_oenb[105]
port 934 nsew signal input
rlabel metal2 s 305642 0 305698 800 6 la_oenb[106]
port 935 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 la_oenb[107]
port 936 nsew signal input
rlabel metal2 s 309966 0 310022 800 6 la_oenb[108]
port 937 nsew signal input
rlabel metal2 s 312174 0 312230 800 6 la_oenb[109]
port 938 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[10]
port 939 nsew signal input
rlabel metal2 s 314290 0 314346 800 6 la_oenb[110]
port 940 nsew signal input
rlabel metal2 s 316406 0 316462 800 6 la_oenb[111]
port 941 nsew signal input
rlabel metal2 s 318614 0 318670 800 6 la_oenb[112]
port 942 nsew signal input
rlabel metal2 s 320730 0 320786 800 6 la_oenb[113]
port 943 nsew signal input
rlabel metal2 s 322846 0 322902 800 6 la_oenb[114]
port 944 nsew signal input
rlabel metal2 s 325054 0 325110 800 6 la_oenb[115]
port 945 nsew signal input
rlabel metal2 s 327170 0 327226 800 6 la_oenb[116]
port 946 nsew signal input
rlabel metal2 s 329378 0 329434 800 6 la_oenb[117]
port 947 nsew signal input
rlabel metal2 s 331494 0 331550 800 6 la_oenb[118]
port 948 nsew signal input
rlabel metal2 s 333610 0 333666 800 6 la_oenb[119]
port 949 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[11]
port 950 nsew signal input
rlabel metal2 s 335818 0 335874 800 6 la_oenb[120]
port 951 nsew signal input
rlabel metal2 s 337934 0 337990 800 6 la_oenb[121]
port 952 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 la_oenb[122]
port 953 nsew signal input
rlabel metal2 s 342258 0 342314 800 6 la_oenb[123]
port 954 nsew signal input
rlabel metal2 s 344374 0 344430 800 6 la_oenb[124]
port 955 nsew signal input
rlabel metal2 s 346582 0 346638 800 6 la_oenb[125]
port 956 nsew signal input
rlabel metal2 s 348698 0 348754 800 6 la_oenb[126]
port 957 nsew signal input
rlabel metal2 s 350814 0 350870 800 6 la_oenb[127]
port 958 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_oenb[12]
port 959 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_oenb[13]
port 960 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_oenb[14]
port 961 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_oenb[15]
port 962 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_oenb[16]
port 963 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_oenb[17]
port 964 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[18]
port 965 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_oenb[19]
port 966 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[1]
port 967 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[20]
port 968 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_oenb[21]
port 969 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_oenb[22]
port 970 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_oenb[23]
port 971 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_oenb[24]
port 972 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[25]
port 973 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[26]
port 974 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_oenb[27]
port 975 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[28]
port 976 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_oenb[29]
port 977 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[2]
port 978 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[30]
port 979 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_oenb[31]
port 980 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_oenb[32]
port 981 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_oenb[33]
port 982 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_oenb[34]
port 983 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[35]
port 984 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oenb[36]
port 985 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 la_oenb[37]
port 986 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_oenb[38]
port 987 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_oenb[39]
port 988 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oenb[3]
port 989 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_oenb[40]
port 990 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oenb[41]
port 991 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_oenb[42]
port 992 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_oenb[43]
port 993 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 la_oenb[44]
port 994 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 la_oenb[45]
port 995 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 la_oenb[46]
port 996 nsew signal input
rlabel metal2 s 178774 0 178830 800 6 la_oenb[47]
port 997 nsew signal input
rlabel metal2 s 180890 0 180946 800 6 la_oenb[48]
port 998 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_oenb[49]
port 999 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[4]
port 1000 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_oenb[50]
port 1001 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_oenb[51]
port 1002 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_oenb[52]
port 1003 nsew signal input
rlabel metal2 s 191654 0 191710 800 6 la_oenb[53]
port 1004 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_oenb[54]
port 1005 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_oenb[55]
port 1006 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_oenb[56]
port 1007 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_oenb[57]
port 1008 nsew signal input
rlabel metal2 s 202418 0 202474 800 6 la_oenb[58]
port 1009 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_oenb[59]
port 1010 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[5]
port 1011 nsew signal input
rlabel metal2 s 206742 0 206798 800 6 la_oenb[60]
port 1012 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 la_oenb[61]
port 1013 nsew signal input
rlabel metal2 s 211066 0 211122 800 6 la_oenb[62]
port 1014 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_oenb[63]
port 1015 nsew signal input
rlabel metal2 s 215298 0 215354 800 6 la_oenb[64]
port 1016 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_oenb[65]
port 1017 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 la_oenb[66]
port 1018 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 la_oenb[67]
port 1019 nsew signal input
rlabel metal2 s 223946 0 224002 800 6 la_oenb[68]
port 1020 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 la_oenb[69]
port 1021 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_oenb[6]
port 1022 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_oenb[70]
port 1023 nsew signal input
rlabel metal2 s 230386 0 230442 800 6 la_oenb[71]
port 1024 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_oenb[72]
port 1025 nsew signal input
rlabel metal2 s 234710 0 234766 800 6 la_oenb[73]
port 1026 nsew signal input
rlabel metal2 s 236826 0 236882 800 6 la_oenb[74]
port 1027 nsew signal input
rlabel metal2 s 239034 0 239090 800 6 la_oenb[75]
port 1028 nsew signal input
rlabel metal2 s 241150 0 241206 800 6 la_oenb[76]
port 1029 nsew signal input
rlabel metal2 s 243266 0 243322 800 6 la_oenb[77]
port 1030 nsew signal input
rlabel metal2 s 245474 0 245530 800 6 la_oenb[78]
port 1031 nsew signal input
rlabel metal2 s 247590 0 247646 800 6 la_oenb[79]
port 1032 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[7]
port 1033 nsew signal input
rlabel metal2 s 249798 0 249854 800 6 la_oenb[80]
port 1034 nsew signal input
rlabel metal2 s 251914 0 251970 800 6 la_oenb[81]
port 1035 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_oenb[82]
port 1036 nsew signal input
rlabel metal2 s 256238 0 256294 800 6 la_oenb[83]
port 1037 nsew signal input
rlabel metal2 s 258354 0 258410 800 6 la_oenb[84]
port 1038 nsew signal input
rlabel metal2 s 260470 0 260526 800 6 la_oenb[85]
port 1039 nsew signal input
rlabel metal2 s 262678 0 262734 800 6 la_oenb[86]
port 1040 nsew signal input
rlabel metal2 s 264794 0 264850 800 6 la_oenb[87]
port 1041 nsew signal input
rlabel metal2 s 267002 0 267058 800 6 la_oenb[88]
port 1042 nsew signal input
rlabel metal2 s 269118 0 269174 800 6 la_oenb[89]
port 1043 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[8]
port 1044 nsew signal input
rlabel metal2 s 271234 0 271290 800 6 la_oenb[90]
port 1045 nsew signal input
rlabel metal2 s 273442 0 273498 800 6 la_oenb[91]
port 1046 nsew signal input
rlabel metal2 s 275558 0 275614 800 6 la_oenb[92]
port 1047 nsew signal input
rlabel metal2 s 277674 0 277730 800 6 la_oenb[93]
port 1048 nsew signal input
rlabel metal2 s 279882 0 279938 800 6 la_oenb[94]
port 1049 nsew signal input
rlabel metal2 s 281998 0 282054 800 6 la_oenb[95]
port 1050 nsew signal input
rlabel metal2 s 284206 0 284262 800 6 la_oenb[96]
port 1051 nsew signal input
rlabel metal2 s 286322 0 286378 800 6 la_oenb[97]
port 1052 nsew signal input
rlabel metal2 s 288438 0 288494 800 6 la_oenb[98]
port 1053 nsew signal input
rlabel metal2 s 290646 0 290702 800 6 la_oenb[99]
port 1054 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[9]
port 1055 nsew signal input
rlabel metal3 s 0 327632 800 327752 6 tag_array_ext_ram_addr1[0]
port 1056 nsew signal output
rlabel metal3 s 0 328448 800 328568 6 tag_array_ext_ram_addr1[1]
port 1057 nsew signal output
rlabel metal3 s 0 329128 800 329248 6 tag_array_ext_ram_addr1[2]
port 1058 nsew signal output
rlabel metal3 s 0 329808 800 329928 6 tag_array_ext_ram_addr1[3]
port 1059 nsew signal output
rlabel metal3 s 0 330488 800 330608 6 tag_array_ext_ram_addr1[4]
port 1060 nsew signal output
rlabel metal3 s 0 331168 800 331288 6 tag_array_ext_ram_addr1[5]
port 1061 nsew signal output
rlabel metal3 s 0 331848 800 331968 6 tag_array_ext_ram_addr1[6]
port 1062 nsew signal output
rlabel metal3 s 0 332664 800 332784 6 tag_array_ext_ram_addr1[7]
port 1063 nsew signal output
rlabel metal3 s 0 272008 800 272128 6 tag_array_ext_ram_addr[0]
port 1064 nsew signal output
rlabel metal3 s 0 272688 800 272808 6 tag_array_ext_ram_addr[1]
port 1065 nsew signal output
rlabel metal3 s 0 273504 800 273624 6 tag_array_ext_ram_addr[2]
port 1066 nsew signal output
rlabel metal3 s 0 274184 800 274304 6 tag_array_ext_ram_addr[3]
port 1067 nsew signal output
rlabel metal3 s 0 274864 800 274984 6 tag_array_ext_ram_addr[4]
port 1068 nsew signal output
rlabel metal3 s 0 275544 800 275664 6 tag_array_ext_ram_addr[5]
port 1069 nsew signal output
rlabel metal3 s 0 276224 800 276344 6 tag_array_ext_ram_addr[6]
port 1070 nsew signal output
rlabel metal3 s 0 277040 800 277160 6 tag_array_ext_ram_addr[7]
port 1071 nsew signal output
rlabel metal3 s 0 277720 800 277840 6 tag_array_ext_ram_clk
port 1072 nsew signal output
rlabel metal3 s 0 324912 800 325032 6 tag_array_ext_ram_csb
port 1073 nsew signal output
rlabel metal3 s 0 326272 800 326392 6 tag_array_ext_ram_csb1[0]
port 1074 nsew signal output
rlabel metal3 s 0 326952 800 327072 6 tag_array_ext_ram_csb1[1]
port 1075 nsew signal output
rlabel metal3 s 0 249568 800 249688 6 tag_array_ext_ram_rdata0[0]
port 1076 nsew signal input
rlabel metal3 s 0 256504 800 256624 6 tag_array_ext_ram_rdata0[10]
port 1077 nsew signal input
rlabel metal3 s 0 257320 800 257440 6 tag_array_ext_ram_rdata0[11]
port 1078 nsew signal input
rlabel metal3 s 0 258000 800 258120 6 tag_array_ext_ram_rdata0[12]
port 1079 nsew signal input
rlabel metal3 s 0 258680 800 258800 6 tag_array_ext_ram_rdata0[13]
port 1080 nsew signal input
rlabel metal3 s 0 259360 800 259480 6 tag_array_ext_ram_rdata0[14]
port 1081 nsew signal input
rlabel metal3 s 0 260040 800 260160 6 tag_array_ext_ram_rdata0[15]
port 1082 nsew signal input
rlabel metal3 s 0 260720 800 260840 6 tag_array_ext_ram_rdata0[16]
port 1083 nsew signal input
rlabel metal3 s 0 261536 800 261656 6 tag_array_ext_ram_rdata0[17]
port 1084 nsew signal input
rlabel metal3 s 0 262216 800 262336 6 tag_array_ext_ram_rdata0[18]
port 1085 nsew signal input
rlabel metal3 s 0 262896 800 263016 6 tag_array_ext_ram_rdata0[19]
port 1086 nsew signal input
rlabel metal3 s 0 250248 800 250368 6 tag_array_ext_ram_rdata0[1]
port 1087 nsew signal input
rlabel metal3 s 0 263576 800 263696 6 tag_array_ext_ram_rdata0[20]
port 1088 nsew signal input
rlabel metal3 s 0 264256 800 264376 6 tag_array_ext_ram_rdata0[21]
port 1089 nsew signal input
rlabel metal3 s 0 265072 800 265192 6 tag_array_ext_ram_rdata0[22]
port 1090 nsew signal input
rlabel metal3 s 0 265752 800 265872 6 tag_array_ext_ram_rdata0[23]
port 1091 nsew signal input
rlabel metal3 s 0 266432 800 266552 6 tag_array_ext_ram_rdata0[24]
port 1092 nsew signal input
rlabel metal3 s 0 267112 800 267232 6 tag_array_ext_ram_rdata0[25]
port 1093 nsew signal input
rlabel metal3 s 0 267792 800 267912 6 tag_array_ext_ram_rdata0[26]
port 1094 nsew signal input
rlabel metal3 s 0 268472 800 268592 6 tag_array_ext_ram_rdata0[27]
port 1095 nsew signal input
rlabel metal3 s 0 269288 800 269408 6 tag_array_ext_ram_rdata0[28]
port 1096 nsew signal input
rlabel metal3 s 0 269968 800 270088 6 tag_array_ext_ram_rdata0[29]
port 1097 nsew signal input
rlabel metal3 s 0 250928 800 251048 6 tag_array_ext_ram_rdata0[2]
port 1098 nsew signal input
rlabel metal3 s 0 270648 800 270768 6 tag_array_ext_ram_rdata0[30]
port 1099 nsew signal input
rlabel metal3 s 0 271328 800 271448 6 tag_array_ext_ram_rdata0[31]
port 1100 nsew signal input
rlabel metal3 s 0 251608 800 251728 6 tag_array_ext_ram_rdata0[3]
port 1101 nsew signal input
rlabel metal3 s 0 252288 800 252408 6 tag_array_ext_ram_rdata0[4]
port 1102 nsew signal input
rlabel metal3 s 0 252968 800 253088 6 tag_array_ext_ram_rdata0[5]
port 1103 nsew signal input
rlabel metal3 s 0 253784 800 253904 6 tag_array_ext_ram_rdata0[6]
port 1104 nsew signal input
rlabel metal3 s 0 254464 800 254584 6 tag_array_ext_ram_rdata0[7]
port 1105 nsew signal input
rlabel metal3 s 0 255144 800 255264 6 tag_array_ext_ram_rdata0[8]
port 1106 nsew signal input
rlabel metal3 s 0 255824 800 255944 6 tag_array_ext_ram_rdata0[9]
port 1107 nsew signal input
rlabel metal3 s 0 333344 800 333464 6 tag_array_ext_ram_rdata1[0]
port 1108 nsew signal input
rlabel metal3 s 0 340416 800 340536 6 tag_array_ext_ram_rdata1[10]
port 1109 nsew signal input
rlabel metal3 s 0 341096 800 341216 6 tag_array_ext_ram_rdata1[11]
port 1110 nsew signal input
rlabel metal3 s 0 341776 800 341896 6 tag_array_ext_ram_rdata1[12]
port 1111 nsew signal input
rlabel metal3 s 0 342456 800 342576 6 tag_array_ext_ram_rdata1[13]
port 1112 nsew signal input
rlabel metal3 s 0 343136 800 343256 6 tag_array_ext_ram_rdata1[14]
port 1113 nsew signal input
rlabel metal3 s 0 343816 800 343936 6 tag_array_ext_ram_rdata1[15]
port 1114 nsew signal input
rlabel metal3 s 0 344632 800 344752 6 tag_array_ext_ram_rdata1[16]
port 1115 nsew signal input
rlabel metal3 s 0 345312 800 345432 6 tag_array_ext_ram_rdata1[17]
port 1116 nsew signal input
rlabel metal3 s 0 345992 800 346112 6 tag_array_ext_ram_rdata1[18]
port 1117 nsew signal input
rlabel metal3 s 0 346672 800 346792 6 tag_array_ext_ram_rdata1[19]
port 1118 nsew signal input
rlabel metal3 s 0 334024 800 334144 6 tag_array_ext_ram_rdata1[1]
port 1119 nsew signal input
rlabel metal3 s 0 347352 800 347472 6 tag_array_ext_ram_rdata1[20]
port 1120 nsew signal input
rlabel metal3 s 0 348168 800 348288 6 tag_array_ext_ram_rdata1[21]
port 1121 nsew signal input
rlabel metal3 s 0 348848 800 348968 6 tag_array_ext_ram_rdata1[22]
port 1122 nsew signal input
rlabel metal3 s 0 349528 800 349648 6 tag_array_ext_ram_rdata1[23]
port 1123 nsew signal input
rlabel metal3 s 0 350208 800 350328 6 tag_array_ext_ram_rdata1[24]
port 1124 nsew signal input
rlabel metal3 s 0 350888 800 351008 6 tag_array_ext_ram_rdata1[25]
port 1125 nsew signal input
rlabel metal3 s 0 351568 800 351688 6 tag_array_ext_ram_rdata1[26]
port 1126 nsew signal input
rlabel metal3 s 0 352384 800 352504 6 tag_array_ext_ram_rdata1[27]
port 1127 nsew signal input
rlabel metal3 s 0 353064 800 353184 6 tag_array_ext_ram_rdata1[28]
port 1128 nsew signal input
rlabel metal3 s 0 353744 800 353864 6 tag_array_ext_ram_rdata1[29]
port 1129 nsew signal input
rlabel metal3 s 0 334704 800 334824 6 tag_array_ext_ram_rdata1[2]
port 1130 nsew signal input
rlabel metal3 s 0 354424 800 354544 6 tag_array_ext_ram_rdata1[30]
port 1131 nsew signal input
rlabel metal3 s 0 355104 800 355224 6 tag_array_ext_ram_rdata1[31]
port 1132 nsew signal input
rlabel metal3 s 0 335384 800 335504 6 tag_array_ext_ram_rdata1[3]
port 1133 nsew signal input
rlabel metal3 s 0 336200 800 336320 6 tag_array_ext_ram_rdata1[4]
port 1134 nsew signal input
rlabel metal3 s 0 336880 800 337000 6 tag_array_ext_ram_rdata1[5]
port 1135 nsew signal input
rlabel metal3 s 0 337560 800 337680 6 tag_array_ext_ram_rdata1[6]
port 1136 nsew signal input
rlabel metal3 s 0 338240 800 338360 6 tag_array_ext_ram_rdata1[7]
port 1137 nsew signal input
rlabel metal3 s 0 338920 800 339040 6 tag_array_ext_ram_rdata1[8]
port 1138 nsew signal input
rlabel metal3 s 0 339600 800 339720 6 tag_array_ext_ram_rdata1[9]
port 1139 nsew signal input
rlabel metal3 s 0 278400 800 278520 6 tag_array_ext_ram_wdata[0]
port 1140 nsew signal output
rlabel metal3 s 0 285472 800 285592 6 tag_array_ext_ram_wdata[10]
port 1141 nsew signal output
rlabel metal3 s 0 286152 800 286272 6 tag_array_ext_ram_wdata[11]
port 1142 nsew signal output
rlabel metal3 s 0 286832 800 286952 6 tag_array_ext_ram_wdata[12]
port 1143 nsew signal output
rlabel metal3 s 0 287512 800 287632 6 tag_array_ext_ram_wdata[13]
port 1144 nsew signal output
rlabel metal3 s 0 288192 800 288312 6 tag_array_ext_ram_wdata[14]
port 1145 nsew signal output
rlabel metal3 s 0 289008 800 289128 6 tag_array_ext_ram_wdata[15]
port 1146 nsew signal output
rlabel metal3 s 0 289688 800 289808 6 tag_array_ext_ram_wdata[16]
port 1147 nsew signal output
rlabel metal3 s 0 290368 800 290488 6 tag_array_ext_ram_wdata[17]
port 1148 nsew signal output
rlabel metal3 s 0 291048 800 291168 6 tag_array_ext_ram_wdata[18]
port 1149 nsew signal output
rlabel metal3 s 0 291728 800 291848 6 tag_array_ext_ram_wdata[19]
port 1150 nsew signal output
rlabel metal3 s 0 279080 800 279200 6 tag_array_ext_ram_wdata[1]
port 1151 nsew signal output
rlabel metal3 s 0 292408 800 292528 6 tag_array_ext_ram_wdata[20]
port 1152 nsew signal output
rlabel metal3 s 0 293224 800 293344 6 tag_array_ext_ram_wdata[21]
port 1153 nsew signal output
rlabel metal3 s 0 293904 800 294024 6 tag_array_ext_ram_wdata[22]
port 1154 nsew signal output
rlabel metal3 s 0 294584 800 294704 6 tag_array_ext_ram_wdata[23]
port 1155 nsew signal output
rlabel metal3 s 0 295264 800 295384 6 tag_array_ext_ram_wdata[24]
port 1156 nsew signal output
rlabel metal3 s 0 295944 800 296064 6 tag_array_ext_ram_wdata[25]
port 1157 nsew signal output
rlabel metal3 s 0 296760 800 296880 6 tag_array_ext_ram_wdata[26]
port 1158 nsew signal output
rlabel metal3 s 0 297440 800 297560 6 tag_array_ext_ram_wdata[27]
port 1159 nsew signal output
rlabel metal3 s 0 298120 800 298240 6 tag_array_ext_ram_wdata[28]
port 1160 nsew signal output
rlabel metal3 s 0 298800 800 298920 6 tag_array_ext_ram_wdata[29]
port 1161 nsew signal output
rlabel metal3 s 0 279760 800 279880 6 tag_array_ext_ram_wdata[2]
port 1162 nsew signal output
rlabel metal3 s 0 299480 800 299600 6 tag_array_ext_ram_wdata[30]
port 1163 nsew signal output
rlabel metal3 s 0 300160 800 300280 6 tag_array_ext_ram_wdata[31]
port 1164 nsew signal output
rlabel metal3 s 0 300976 800 301096 6 tag_array_ext_ram_wdata[32]
port 1165 nsew signal output
rlabel metal3 s 0 301656 800 301776 6 tag_array_ext_ram_wdata[33]
port 1166 nsew signal output
rlabel metal3 s 0 302336 800 302456 6 tag_array_ext_ram_wdata[34]
port 1167 nsew signal output
rlabel metal3 s 0 303016 800 303136 6 tag_array_ext_ram_wdata[35]
port 1168 nsew signal output
rlabel metal3 s 0 303696 800 303816 6 tag_array_ext_ram_wdata[36]
port 1169 nsew signal output
rlabel metal3 s 0 304376 800 304496 6 tag_array_ext_ram_wdata[37]
port 1170 nsew signal output
rlabel metal3 s 0 305192 800 305312 6 tag_array_ext_ram_wdata[38]
port 1171 nsew signal output
rlabel metal3 s 0 305872 800 305992 6 tag_array_ext_ram_wdata[39]
port 1172 nsew signal output
rlabel metal3 s 0 280440 800 280560 6 tag_array_ext_ram_wdata[3]
port 1173 nsew signal output
rlabel metal3 s 0 306552 800 306672 6 tag_array_ext_ram_wdata[40]
port 1174 nsew signal output
rlabel metal3 s 0 307232 800 307352 6 tag_array_ext_ram_wdata[41]
port 1175 nsew signal output
rlabel metal3 s 0 307912 800 308032 6 tag_array_ext_ram_wdata[42]
port 1176 nsew signal output
rlabel metal3 s 0 308728 800 308848 6 tag_array_ext_ram_wdata[43]
port 1177 nsew signal output
rlabel metal3 s 0 309408 800 309528 6 tag_array_ext_ram_wdata[44]
port 1178 nsew signal output
rlabel metal3 s 0 310088 800 310208 6 tag_array_ext_ram_wdata[45]
port 1179 nsew signal output
rlabel metal3 s 0 310768 800 310888 6 tag_array_ext_ram_wdata[46]
port 1180 nsew signal output
rlabel metal3 s 0 311448 800 311568 6 tag_array_ext_ram_wdata[47]
port 1181 nsew signal output
rlabel metal3 s 0 312128 800 312248 6 tag_array_ext_ram_wdata[48]
port 1182 nsew signal output
rlabel metal3 s 0 312944 800 313064 6 tag_array_ext_ram_wdata[49]
port 1183 nsew signal output
rlabel metal3 s 0 281256 800 281376 6 tag_array_ext_ram_wdata[4]
port 1184 nsew signal output
rlabel metal3 s 0 313624 800 313744 6 tag_array_ext_ram_wdata[50]
port 1185 nsew signal output
rlabel metal3 s 0 314304 800 314424 6 tag_array_ext_ram_wdata[51]
port 1186 nsew signal output
rlabel metal3 s 0 314984 800 315104 6 tag_array_ext_ram_wdata[52]
port 1187 nsew signal output
rlabel metal3 s 0 315664 800 315784 6 tag_array_ext_ram_wdata[53]
port 1188 nsew signal output
rlabel metal3 s 0 316480 800 316600 6 tag_array_ext_ram_wdata[54]
port 1189 nsew signal output
rlabel metal3 s 0 317160 800 317280 6 tag_array_ext_ram_wdata[55]
port 1190 nsew signal output
rlabel metal3 s 0 317840 800 317960 6 tag_array_ext_ram_wdata[56]
port 1191 nsew signal output
rlabel metal3 s 0 318520 800 318640 6 tag_array_ext_ram_wdata[57]
port 1192 nsew signal output
rlabel metal3 s 0 319200 800 319320 6 tag_array_ext_ram_wdata[58]
port 1193 nsew signal output
rlabel metal3 s 0 319880 800 320000 6 tag_array_ext_ram_wdata[59]
port 1194 nsew signal output
rlabel metal3 s 0 281936 800 282056 6 tag_array_ext_ram_wdata[5]
port 1195 nsew signal output
rlabel metal3 s 0 320696 800 320816 6 tag_array_ext_ram_wdata[60]
port 1196 nsew signal output
rlabel metal3 s 0 321376 800 321496 6 tag_array_ext_ram_wdata[61]
port 1197 nsew signal output
rlabel metal3 s 0 322056 800 322176 6 tag_array_ext_ram_wdata[62]
port 1198 nsew signal output
rlabel metal3 s 0 322736 800 322856 6 tag_array_ext_ram_wdata[63]
port 1199 nsew signal output
rlabel metal3 s 0 282616 800 282736 6 tag_array_ext_ram_wdata[6]
port 1200 nsew signal output
rlabel metal3 s 0 283296 800 283416 6 tag_array_ext_ram_wdata[7]
port 1201 nsew signal output
rlabel metal3 s 0 283976 800 284096 6 tag_array_ext_ram_wdata[8]
port 1202 nsew signal output
rlabel metal3 s 0 284792 800 284912 6 tag_array_ext_ram_wdata[9]
port 1203 nsew signal output
rlabel metal3 s 0 325592 800 325712 6 tag_array_ext_ram_web
port 1204 nsew signal output
rlabel metal3 s 0 323416 800 323536 6 tag_array_ext_ram_wmask[0]
port 1205 nsew signal output
rlabel metal3 s 0 324096 800 324216 6 tag_array_ext_ram_wmask[1]
port 1206 nsew signal output
rlabel metal4 s 4208 2128 4528 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 34928 2128 35248 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 65648 2128 65968 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 96368 2128 96688 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 127088 2128 127408 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 157808 2128 158128 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 188528 2128 188848 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 219248 2128 219568 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 249968 2128 250288 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 280688 2128 281008 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 311408 2128 311728 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 342128 2128 342448 353104 6 vccd1
port 1207 nsew power input
rlabel metal4 s 19568 2128 19888 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 50288 2128 50608 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 81008 2128 81328 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 111728 2128 112048 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 142448 2128 142768 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 173168 2128 173488 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 203888 2128 204208 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 234608 2128 234928 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 265328 2128 265648 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 296048 2128 296368 353104 6 vssd1
port 1208 nsew ground input
rlabel metal4 s 326768 2128 327088 353104 6 vssd1
port 1208 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 1209 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 1210 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_ack_o
port 1211 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[0]
port 1212 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[10]
port 1213 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[11]
port 1214 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[12]
port 1215 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_adr_i[13]
port 1216 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_adr_i[14]
port 1217 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_adr_i[15]
port 1218 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_adr_i[16]
port 1219 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 wbs_adr_i[17]
port 1220 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_adr_i[18]
port 1221 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[19]
port 1222 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[1]
port 1223 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[20]
port 1224 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 wbs_adr_i[21]
port 1225 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 wbs_adr_i[22]
port 1226 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_adr_i[23]
port 1227 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 wbs_adr_i[24]
port 1228 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[25]
port 1229 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 wbs_adr_i[26]
port 1230 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 wbs_adr_i[27]
port 1231 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 wbs_adr_i[28]
port 1232 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 wbs_adr_i[29]
port 1233 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[2]
port 1234 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 wbs_adr_i[30]
port 1235 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_adr_i[31]
port 1236 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_adr_i[3]
port 1237 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[4]
port 1238 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_adr_i[5]
port 1239 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[6]
port 1240 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[7]
port 1241 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[8]
port 1242 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[9]
port 1243 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_cyc_i
port 1244 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_i[0]
port 1245 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_i[10]
port 1246 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[11]
port 1247 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[12]
port 1248 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[13]
port 1249 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[14]
port 1250 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_i[15]
port 1251 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[16]
port 1252 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_i[17]
port 1253 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_i[18]
port 1254 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_i[19]
port 1255 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[1]
port 1256 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[20]
port 1257 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 wbs_dat_i[21]
port 1258 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_i[22]
port 1259 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_i[23]
port 1260 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_i[24]
port 1261 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_i[25]
port 1262 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_i[26]
port 1263 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 wbs_dat_i[27]
port 1264 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_i[28]
port 1265 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 wbs_dat_i[29]
port 1266 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[2]
port 1267 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 wbs_dat_i[30]
port 1268 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 wbs_dat_i[31]
port 1269 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[3]
port 1270 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[4]
port 1271 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[5]
port 1272 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[6]
port 1273 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[7]
port 1274 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[8]
port 1275 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[9]
port 1276 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_o[0]
port 1277 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[10]
port 1278 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_o[11]
port 1279 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_o[12]
port 1280 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[13]
port 1281 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_o[14]
port 1282 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[15]
port 1283 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_o[16]
port 1284 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_o[17]
port 1285 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[18]
port 1286 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_o[19]
port 1287 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[1]
port 1288 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_o[20]
port 1289 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_o[21]
port 1290 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 wbs_dat_o[22]
port 1291 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_o[23]
port 1292 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[24]
port 1293 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 wbs_dat_o[25]
port 1294 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_o[26]
port 1295 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 wbs_dat_o[27]
port 1296 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 wbs_dat_o[28]
port 1297 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 wbs_dat_o[29]
port 1298 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[2]
port 1299 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_o[30]
port 1300 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_o[31]
port 1301 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[3]
port 1302 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[4]
port 1303 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[5]
port 1304 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_o[6]
port 1305 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[7]
port 1306 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[8]
port 1307 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[9]
port 1308 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_sel_i[0]
port 1309 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_sel_i[1]
port 1310 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_sel_i[2]
port 1311 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_sel_i[3]
port 1312 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_stb_i
port 1313 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_we_i
port 1314 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 353479 355623
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 306684690
string GDS_FILE /home/shc/Development/efabless/marmot_asic/openlane/marmot/runs/marmot/results/finishing/Marmot.magic.gds
string GDS_START 2048228
<< end >>

