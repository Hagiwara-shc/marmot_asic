// xip.hex
case (address)
  11'h000: out <= 32'h08002137;
  11'h001: out <= 32'hff010113;
  11'h002: out <= 32'h006f2cf5;
  11'h003: out <= 32'hf5930000;
  11'h004: out <= 32'h07330ff5;
  11'h005: out <= 32'h87aa00c5;
  11'h006: out <= 32'h00c05763;
  11'h007: out <= 32'h8fa30785;
  11'h008: out <= 32'h1de3feb7;
  11'h009: out <= 32'h8082fef7;
  11'h00a: out <= 32'h00c05c63;
  11'h00b: out <= 32'h87aa962a;
  11'h00c: out <= 32'h0005c703;
  11'h00d: out <= 32'h05850785;
  11'h00e: out <= 32'hfee78fa3;
  11'h00f: out <= 32'hfef61ae3;
  11'h010: out <= 32'h55638082;
  11'h011: out <= 32'h962e02c0;
  11'h012: out <= 32'h0163a019;
  11'h013: out <= 32'h478302b6;
  11'h014: out <= 32'hc7030005;
  11'h015: out <= 32'h05050005;
  11'h016: out <= 32'h88e30585;
  11'h017: out <= 32'h3533fee7;
  11'h018: out <= 32'h053300f7;
  11'h019: out <= 32'h890940a0;
  11'h01a: out <= 32'h8082157d;
  11'h01b: out <= 32'h80824501;
  11'h01c: out <= 32'h00054783;
  11'h01d: out <= 32'h4501872a;
  11'h01e: out <= 32'h0505cb81;
  11'h01f: out <= 32'h00a707b3;
  11'h020: out <= 32'h0007c783;
  11'h021: out <= 32'h8082fbfd;
  11'h022: out <= 32'hc7838082;
  11'h023: out <= 32'h00230005;
  11'h024: out <= 32'hc78300f5;
  11'h025: out <= 32'hcb990005;
  11'h026: out <= 32'hc70387aa;
  11'h027: out <= 32'h05850015;
  11'h028: out <= 32'h80230785;
  11'h029: out <= 32'hc70300e7;
  11'h02a: out <= 32'hfb650005;
  11'h02b: out <= 32'ha0198082;
  11'h02c: out <= 32'h00e79d63;
  11'h02d: out <= 32'h00054783;
  11'h02e: out <= 32'h0005c703;
  11'h02f: out <= 32'h05850505;
  11'h030: out <= 32'h00e7e6b3;
  11'h031: out <= 32'h4501f6f5;
  11'h032: out <= 32'h35338082;
  11'h033: out <= 32'h053300f7;
  11'h034: out <= 32'h890940a0;
  11'h035: out <= 32'h8082157d;
  11'h036: out <= 32'h083387aa;
  11'h037: out <= 32'hc70300c5;
  11'h038: out <= 32'h06b30007;
  11'h039: out <= 32'heb1940f8;
  11'h03a: out <= 32'h0005c703;
  11'h03b: out <= 32'h9532c70d;
  11'h03c: out <= 32'h25338d1d;
  11'h03d: out <= 32'h053300a0;
  11'h03e: out <= 32'h808240a0;
  11'h03f: out <= 32'h00d05d63;
  11'h040: out <= 32'h0005c683;
  11'h041: out <= 32'h05850785;
  11'h042: out <= 32'hfce68be3;
  11'h043: out <= 32'he6e34505;
  11'h044: out <= 32'h557dfee6;
  11'h045: out <= 32'h45018082;
  11'h046: out <= 32'h11418082;
  11'h047: out <= 32'hc606c422;
  11'h048: out <= 32'h842a47a9;
  11'h049: out <= 32'h00f50863;
  11'h04a: out <= 32'h442285a2;
  11'h04b: out <= 32'h450140b2;
  11'h04c: out <= 32'ha2490141;
  11'h04d: out <= 32'h450145b5;
  11'h04e: out <= 32'h85a22ab5;
  11'h04f: out <= 32'h40b24422;
  11'h050: out <= 32'h01414501;
  11'h051: out <= 32'h1141aa85;
  11'h052: out <= 32'hc4224501;
  11'h053: out <= 32'h2a71c606;
  11'h054: out <= 32'h442947b5;
  11'h055: out <= 32'h00f50363;
  11'h056: out <= 32'h8522842a;
  11'h057: out <= 32'h40b23f7d;
  11'h058: out <= 32'h44228522;
  11'h059: out <= 32'h80820141;
  11'h05a: out <= 32'hc4221141;
  11'h05b: out <= 32'h842ac606;
  11'h05c: out <= 32'h00054503;
  11'h05d: out <= 32'h0405c511;
  11'h05e: out <= 32'h4503374d;
  11'h05f: out <= 32'hfd650004;
  11'h060: out <= 32'h442240b2;
  11'h061: out <= 32'h01414501;
  11'h062: out <= 32'h11418082;
  11'h063: out <= 32'hc226c422;
  11'h064: out <= 32'hc606c04a;
  11'h065: out <= 32'h842a4929;
  11'h066: out <= 32'h37754481;
  11'h067: out <= 32'h01250c63;
  11'h068: out <= 32'h00a40023;
  11'h069: out <= 32'h00148793;
  11'h06a: out <= 32'hc5190405;
  11'h06b: out <= 32'h3f6184be;
  11'h06c: out <= 32'hff2518e3;
  11'h06d: out <= 32'h00040023;
  11'h06e: out <= 32'h442240b2;
  11'h06f: out <= 32'h85264902;
  11'h070: out <= 32'h01414492;
  11'h071: out <= 32'h11018082;
  11'h072: out <= 32'hcc22ce06;
  11'h073: out <= 32'h00010623;
  11'h074: out <= 32'he191ed05;
  11'h075: out <= 32'h07934585;
  11'h076: out <= 32'h071300b1;
  11'h077: out <= 32'hc5910300;
  11'h078: out <= 32'h00e78023;
  11'h079: out <= 32'h17fd15fd;
  11'h07a: out <= 32'hc503fde5;
  11'h07b: out <= 32'h84130017;
  11'h07c: out <= 32'hc5110017;
  11'h07d: out <= 32'h37150405;
  11'h07e: out <= 32'h00044503;
  11'h07f: out <= 32'h40f2fd65;
  11'h080: out <= 32'h45014462;
  11'h081: out <= 32'h80826105;
  11'h082: out <= 32'h6841872a;
  11'h083: out <= 32'h00f77793;
  11'h084: out <= 32'h37880813;
  11'h085: out <= 32'hc50397c2;
  11'h086: out <= 32'h04130007;
  11'h087: out <= 32'h079300b1;
  11'h088: out <= 32'h80a3fff4;
  11'h089: out <= 32'h831100a7;
  11'h08a: out <= 32'h15fdcd99;
  11'h08b: out <= 32'h843ed75d;
  11'h08c: out <= 32'h00f77793;
  11'h08d: out <= 32'hc50397c2;
  11'h08e: out <= 32'h83110007;
  11'h08f: out <= 32'hfff40793;
  11'h090: out <= 32'h00a780a3;
  11'h091: out <= 32'h7693f1fd;
  11'h092: out <= 32'h96c200f7;
  11'h093: out <= 32'hfff78613;
  11'h094: out <= 32'hc503d34d;
  11'h095: out <= 32'h83110006;
  11'h096: out <= 32'h8023843e;
  11'h097: out <= 32'h769300a7;
  11'h098: out <= 32'h87b200f7;
  11'h099: out <= 32'h861396c2;
  11'h09a: out <= 32'hd741fff7;
  11'h09b: out <= 32'h1793b7dd;
  11'h09c: out <= 32'h65410025;
  11'h09d: out <= 32'h36050513;
  11'h09e: out <= 32'h4118953e;
  11'h09f: out <= 32'hc71c4785;
  11'h0a0: out <= 32'h8a63c75c;
  11'h0a1: out <= 32'h079300f5;
  11'h0a2: out <= 32'hcf1c3630;
  11'h0a3: out <= 32'hdfe3435c;
  11'h0a4: out <= 32'h4501fe07;
  11'h0a5: out <= 32'h47bd8082;
  11'h0a6: out <= 32'hbfcdcf1c;
  11'h0a7: out <= 32'h00251793;
  11'h0a8: out <= 32'h05136541;
  11'h0a9: out <= 32'h953e3605;
  11'h0aa: out <= 32'h4388411c;
  11'h0ab: out <= 32'hfff54513;
  11'h0ac: out <= 32'h8082817d;
  11'h0ad: out <= 32'h00251793;
  11'h0ae: out <= 32'h05136541;
  11'h0af: out <= 32'h953e3605;
  11'h0b0: out <= 32'h431c4118;
  11'h0b1: out <= 32'hfe07cfe3;
  11'h0b2: out <= 32'h4501c30c;
  11'h0b3: out <= 32'h17938082;
  11'h0b4: out <= 32'h65410025;
  11'h0b5: out <= 32'h36050513;
  11'h0b6: out <= 32'h411c953e;
  11'h0b7: out <= 32'hc51343dc;
  11'h0b8: out <= 32'h8023fff7;
  11'h0b9: out <= 32'h817d00f5;
  11'h0ba: out <= 32'h17938082;
  11'h0bb: out <= 32'h65410025;
  11'h0bc: out <= 32'h36050513;
  11'h0bd: out <= 32'h411c953e;
  11'h0be: out <= 32'h4fe343c8;
  11'h0bf: out <= 32'h7513fe05;
  11'h0c0: out <= 32'h80820ff5;
  11'h0c1: out <= 32'h08000537;
  11'h0c2: out <= 32'h080007b7;
  11'h0c3: out <= 32'h00478793;
  11'h0c4: out <= 32'h00050613;
  11'h0c5: out <= 32'h114165c1;
  11'h0c6: out <= 32'h40c78633;
  11'h0c7: out <= 32'h38c58593;
  11'h0c8: out <= 32'h00050513;
  11'h0c9: out <= 32'h3309c606;
  11'h0ca: out <= 32'h08000537;
  11'h0cb: out <= 32'h080007b7;
  11'h0cc: out <= 32'h00478793;
  11'h0cd: out <= 32'h00450613;
  11'h0ce: out <= 32'h40c78633;
  11'h0cf: out <= 32'h05134581;
  11'h0d0: out <= 32'h31f10045;
  11'h0d1: out <= 32'h080007b7;
  11'h0d2: out <= 32'h0007a583;
  11'h0d3: out <= 32'h37054501;
  11'h0d4: out <= 32'h202007b7;
  11'h0d5: out <= 32'h40b29782;
  11'h0d6: out <= 32'h01414501;
  11'h0d7: out <= 32'h00008082;
  11'h0d8: out <= 32'h10013000;
  11'h0d9: out <= 32'h10023000;
  11'h0da: out <= 32'h10033000;
  11'h0db: out <= 32'h10043000;
  11'h0dc: out <= 32'h10053000;
  11'h0dd: out <= 32'h10063000;
  11'h0de: out <= 32'h33323130;
  11'h0df: out <= 32'h37363534;
  11'h0e0: out <= 32'h62613938;
  11'h0e1: out <= 32'h66656463;
  11'h0e2: out <= 32'h00000000;
  11'h0e3: out <= 32'h00000001;
  default: out <= 32'hdeadbeef;
endcase
