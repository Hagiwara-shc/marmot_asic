// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module marmot
(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // IRQ
    output [2:0] irq
);

    wire clk;
    wire rst;

    // Assuming LA probes [65:64] are for controlling the count clk & reset  
    assign clk = (~la_oenb[64]) ? la_data_in[64]: wb_clk_i;
    assign rst = (~la_oenb[65]) ? la_data_in[65]: wb_rst_i;

 MarmotCaravelChip MarmotCaravelChip (
  .wb_clk_i(clk),
  .wb_rst_i(rst),
  .wbs_stb_i(wbs_stb_i),
  .wbs_cyc_i(wbs_cyc_i),
  .wbs_we_i(wbs_we_i),
  .wbs_sel_i_0(wbs_sel_i[0]),
  .wbs_sel_i_1(wbs_sel_i[1]),
  .wbs_sel_i_2(wbs_sel_i[2]),
  .wbs_sel_i_3(wbs_sel_i[3]),
  .wbs_dat_i_0(wbs_dat_i[0]),
  .wbs_dat_i_1(wbs_dat_i[1]),
  .wbs_dat_i_2(wbs_dat_i[2]),
  .wbs_dat_i_3(wbs_dat_i[3]),
  .wbs_dat_i_4(wbs_dat_i[4]),
  .wbs_dat_i_5(wbs_dat_i[5]),
  .wbs_dat_i_6(wbs_dat_i[6]),
  .wbs_dat_i_7(wbs_dat_i[7]),
  .wbs_dat_i_8(wbs_dat_i[8]),
  .wbs_dat_i_9(wbs_dat_i[9]),
  .wbs_dat_i_10(wbs_dat_i[10]),
  .wbs_dat_i_11(wbs_dat_i[11]),
  .wbs_dat_i_12(wbs_dat_i[12]),
  .wbs_dat_i_13(wbs_dat_i[13]),
  .wbs_dat_i_14(wbs_dat_i[14]),
  .wbs_dat_i_15(wbs_dat_i[15]),
  .wbs_dat_i_16(wbs_dat_i[16]),
  .wbs_dat_i_17(wbs_dat_i[17]),
  .wbs_dat_i_18(wbs_dat_i[18]),
  .wbs_dat_i_19(wbs_dat_i[19]),
  .wbs_dat_i_20(wbs_dat_i[20]),
  .wbs_dat_i_21(wbs_dat_i[21]),
  .wbs_dat_i_22(wbs_dat_i[22]),
  .wbs_dat_i_23(wbs_dat_i[23]),
  .wbs_dat_i_24(wbs_dat_i[24]),
  .wbs_dat_i_25(wbs_dat_i[25]),
  .wbs_dat_i_26(wbs_dat_i[26]),
  .wbs_dat_i_27(wbs_dat_i[27]),
  .wbs_dat_i_28(wbs_dat_i[28]),
  .wbs_dat_i_29(wbs_dat_i[29]),
  .wbs_dat_i_30(wbs_dat_i[30]),
  .wbs_dat_i_31(wbs_dat_i[31]),
  .wbs_ack_o(wbs_ack_o),
  .wbs_dat_o_0(wbs_dat_o[0]),
  .wbs_dat_o_1(wbs_dat_o[1]),
  .wbs_dat_o_2(wbs_dat_o[2]),
  .wbs_dat_o_3(wbs_dat_o[3]),
  .wbs_dat_o_4(wbs_dat_o[4]),
  .wbs_dat_o_5(wbs_dat_o[5]),
  .wbs_dat_o_6(wbs_dat_o[6]),
  .wbs_dat_o_7(wbs_dat_o[7]),
  .wbs_dat_o_8(wbs_dat_o[8]),
  .wbs_dat_o_9(wbs_dat_o[9]),
  .wbs_dat_o_10(wbs_dat_o[10]),
  .wbs_dat_o_11(wbs_dat_o[11]),
  .wbs_dat_o_12(wbs_dat_o[12]),
  .wbs_dat_o_13(wbs_dat_o[13]),
  .wbs_dat_o_14(wbs_dat_o[14]),
  .wbs_dat_o_15(wbs_dat_o[15]),
  .wbs_dat_o_16(wbs_dat_o[16]),
  .wbs_dat_o_17(wbs_dat_o[17]),
  .wbs_dat_o_18(wbs_dat_o[18]),
  .wbs_dat_o_19(wbs_dat_o[19]),
  .wbs_dat_o_20(wbs_dat_o[20]),
  .wbs_dat_o_21(wbs_dat_o[21]),
  .wbs_dat_o_22(wbs_dat_o[22]),
  .wbs_dat_o_23(wbs_dat_o[23]),
  .wbs_dat_o_24(wbs_dat_o[24]),
  .wbs_dat_o_25(wbs_dat_o[25]),
  .wbs_dat_o_26(wbs_dat_o[26]),
  .wbs_dat_o_27(wbs_dat_o[27]),
  .wbs_dat_o_28(wbs_dat_o[28]),
  .wbs_dat_o_29(wbs_dat_o[29]),
  .wbs_dat_o_30(wbs_dat_o[30]),
  .wbs_dat_o_31(wbs_dat_o[31]),
  .la_data_in_0(la_data_in[0]),
  .la_data_in_1(la_data_in[1]),
  .la_data_in_2(la_data_in[2]),
  .la_data_in_3(la_data_in[3]),
  .la_data_in_4(la_data_in[4]),
  .la_data_in_5(la_data_in[5]),
  .la_data_in_6(la_data_in[6]),
  .la_data_in_7(la_data_in[7]),
  .la_data_in_8(la_data_in[8]),
  .la_data_in_9(la_data_in[9]),
  .la_data_in_10(la_data_in[10]),
  .la_data_in_11(la_data_in[11]),
  .la_data_in_12(la_data_in[12]),
  .la_data_in_13(la_data_in[13]),
  .la_data_in_14(la_data_in[14]),
  .la_data_in_15(la_data_in[15]),
  .la_data_in_16(la_data_in[16]),
  .la_data_in_17(la_data_in[17]),
  .la_data_in_18(la_data_in[18]),
  .la_data_in_19(la_data_in[19]),
  .la_data_in_20(la_data_in[20]),
  .la_data_in_21(la_data_in[21]),
  .la_data_in_22(la_data_in[22]),
  .la_data_in_23(la_data_in[23]),
  .la_data_in_24(la_data_in[24]),
  .la_data_in_25(la_data_in[25]),
  .la_data_in_26(la_data_in[26]),
  .la_data_in_27(la_data_in[27]),
  .la_data_in_28(la_data_in[28]),
  .la_data_in_29(la_data_in[29]),
  .la_data_in_30(la_data_in[30]),
  .la_data_in_31(la_data_in[31]),
  .la_data_in_32(la_data_in[32]),
  .la_data_in_33(la_data_in[33]),
  .la_data_in_34(la_data_in[34]),
  .la_data_in_35(la_data_in[35]),
  .la_data_in_36(la_data_in[36]),
  .la_data_in_37(la_data_in[37]),
  .la_data_in_38(la_data_in[38]),
  .la_data_in_39(la_data_in[39]),
  .la_data_in_40(la_data_in[40]),
  .la_data_in_41(la_data_in[41]),
  .la_data_in_42(la_data_in[42]),
  .la_data_in_43(la_data_in[43]),
  .la_data_in_44(la_data_in[44]),
  .la_data_in_45(la_data_in[45]),
  .la_data_in_46(la_data_in[46]),
  .la_data_in_47(la_data_in[47]),
  .la_data_in_48(la_data_in[48]),
  .la_data_in_49(la_data_in[49]),
  .la_data_in_50(la_data_in[50]),
  .la_data_in_51(la_data_in[51]),
  .la_data_in_52(la_data_in[52]),
  .la_data_in_53(la_data_in[53]),
  .la_data_in_54(la_data_in[54]),
  .la_data_in_55(la_data_in[55]),
  .la_data_in_56(la_data_in[56]),
  .la_data_in_57(la_data_in[57]),
  .la_data_in_58(la_data_in[58]),
  .la_data_in_59(la_data_in[59]),
  .la_data_in_60(la_data_in[60]),
  .la_data_in_61(la_data_in[61]),
  .la_data_in_62(la_data_in[62]),
  .la_data_in_63(la_data_in[63]),
  .la_data_in_64(la_data_in[64]),
  .la_data_in_65(la_data_in[65]),
  .la_data_in_66(la_data_in[66]),
  .la_data_in_67(la_data_in[67]),
  .la_data_in_68(la_data_in[68]),
  .la_data_in_69(la_data_in[69]),
  .la_data_in_70(la_data_in[70]),
  .la_data_in_71(la_data_in[71]),
  .la_data_in_72(la_data_in[72]),
  .la_data_in_73(la_data_in[73]),
  .la_data_in_74(la_data_in[74]),
  .la_data_in_75(la_data_in[75]),
  .la_data_in_76(la_data_in[76]),
  .la_data_in_77(la_data_in[77]),
  .la_data_in_78(la_data_in[78]),
  .la_data_in_79(la_data_in[79]),
  .la_data_in_80(la_data_in[80]),
  .la_data_in_81(la_data_in[81]),
  .la_data_in_82(la_data_in[82]),
  .la_data_in_83(la_data_in[83]),
  .la_data_in_84(la_data_in[84]),
  .la_data_in_85(la_data_in[85]),
  .la_data_in_86(la_data_in[86]),
  .la_data_in_87(la_data_in[87]),
  .la_data_in_88(la_data_in[88]),
  .la_data_in_89(la_data_in[89]),
  .la_data_in_90(la_data_in[90]),
  .la_data_in_91(la_data_in[91]),
  .la_data_in_92(la_data_in[92]),
  .la_data_in_93(la_data_in[93]),
  .la_data_in_94(la_data_in[94]),
  .la_data_in_95(la_data_in[95]),
  .la_data_in_96(la_data_in[96]),
  .la_data_in_97(la_data_in[97]),
  .la_data_in_98(la_data_in[98]),
  .la_data_in_99(la_data_in[99]),
  .la_data_in_100(la_data_in[100]),
  .la_data_in_101(la_data_in[101]),
  .la_data_in_102(la_data_in[102]),
  .la_data_in_103(la_data_in[103]),
  .la_data_in_104(la_data_in[104]),
  .la_data_in_105(la_data_in[105]),
  .la_data_in_106(la_data_in[106]),
  .la_data_in_107(la_data_in[107]),
  .la_data_in_108(la_data_in[108]),
  .la_data_in_109(la_data_in[109]),
  .la_data_in_110(la_data_in[110]),
  .la_data_in_111(la_data_in[111]),
  .la_data_in_112(la_data_in[112]),
  .la_data_in_113(la_data_in[113]),
  .la_data_in_114(la_data_in[114]),
  .la_data_in_115(la_data_in[115]),
  .la_data_in_116(la_data_in[116]),
  .la_data_in_117(la_data_in[117]),
  .la_data_in_118(la_data_in[118]),
  .la_data_in_119(la_data_in[119]),
  .la_data_in_120(la_data_in[120]),
  .la_data_in_121(la_data_in[121]),
  .la_data_in_122(la_data_in[122]),
  .la_data_in_123(la_data_in[123]),
  .la_data_in_124(la_data_in[124]),
  .la_data_in_125(la_data_in[125]),
  .la_data_in_126(la_data_in[126]),
  .la_data_in_127(la_data_in[127]),
  .la_data_out_0(la_data_out[0]),
  .la_data_out_1(la_data_out[1]),
  .la_data_out_2(la_data_out[2]),
  .la_data_out_3(la_data_out[3]),
  .la_data_out_4(la_data_out[4]),
  .la_data_out_5(la_data_out[5]),
  .la_data_out_6(la_data_out[6]),
  .la_data_out_7(la_data_out[7]),
  .la_data_out_8(la_data_out[8]),
  .la_data_out_9(la_data_out[9]),
  .la_data_out_10(la_data_out[10]),
  .la_data_out_11(la_data_out[11]),
  .la_data_out_12(la_data_out[12]),
  .la_data_out_13(la_data_out[13]),
  .la_data_out_14(la_data_out[14]),
  .la_data_out_15(la_data_out[15]),
  .la_data_out_16(la_data_out[16]),
  .la_data_out_17(la_data_out[17]),
  .la_data_out_18(la_data_out[18]),
  .la_data_out_19(la_data_out[19]),
  .la_data_out_20(la_data_out[20]),
  .la_data_out_21(la_data_out[21]),
  .la_data_out_22(la_data_out[22]),
  .la_data_out_23(la_data_out[23]),
  .la_data_out_24(la_data_out[24]),
  .la_data_out_25(la_data_out[25]),
  .la_data_out_26(la_data_out[26]),
  .la_data_out_27(la_data_out[27]),
  .la_data_out_28(la_data_out[28]),
  .la_data_out_29(la_data_out[29]),
  .la_data_out_30(la_data_out[30]),
  .la_data_out_31(la_data_out[31]),
  .la_data_out_32(la_data_out[32]),
  .la_data_out_33(la_data_out[33]),
  .la_data_out_34(la_data_out[34]),
  .la_data_out_35(la_data_out[35]),
  .la_data_out_36(la_data_out[36]),
  .la_data_out_37(la_data_out[37]),
  .la_data_out_38(la_data_out[38]),
  .la_data_out_39(la_data_out[39]),
  .la_data_out_40(la_data_out[40]),
  .la_data_out_41(la_data_out[41]),
  .la_data_out_42(la_data_out[42]),
  .la_data_out_43(la_data_out[43]),
  .la_data_out_44(la_data_out[44]),
  .la_data_out_45(la_data_out[45]),
  .la_data_out_46(la_data_out[46]),
  .la_data_out_47(la_data_out[47]),
  .la_data_out_48(la_data_out[48]),
  .la_data_out_49(la_data_out[49]),
  .la_data_out_50(la_data_out[50]),
  .la_data_out_51(la_data_out[51]),
  .la_data_out_52(la_data_out[52]),
  .la_data_out_53(la_data_out[53]),
  .la_data_out_54(la_data_out[54]),
  .la_data_out_55(la_data_out[55]),
  .la_data_out_56(la_data_out[56]),
  .la_data_out_57(la_data_out[57]),
  .la_data_out_58(la_data_out[58]),
  .la_data_out_59(la_data_out[59]),
  .la_data_out_60(la_data_out[60]),
  .la_data_out_61(la_data_out[61]),
  .la_data_out_62(la_data_out[62]),
  .la_data_out_63(la_data_out[63]),
  .la_data_out_64(la_data_out[64]),
  .la_data_out_65(la_data_out[65]),
  .la_data_out_66(la_data_out[66]),
  .la_data_out_67(la_data_out[67]),
  .la_data_out_68(la_data_out[68]),
  .la_data_out_69(la_data_out[69]),
  .la_data_out_70(la_data_out[70]),
  .la_data_out_71(la_data_out[71]),
  .la_data_out_72(la_data_out[72]),
  .la_data_out_73(la_data_out[73]),
  .la_data_out_74(la_data_out[74]),
  .la_data_out_75(la_data_out[75]),
  .la_data_out_76(la_data_out[76]),
  .la_data_out_77(la_data_out[77]),
  .la_data_out_78(la_data_out[78]),
  .la_data_out_79(la_data_out[79]),
  .la_data_out_80(la_data_out[80]),
  .la_data_out_81(la_data_out[81]),
  .la_data_out_82(la_data_out[82]),
  .la_data_out_83(la_data_out[83]),
  .la_data_out_84(la_data_out[84]),
  .la_data_out_85(la_data_out[85]),
  .la_data_out_86(la_data_out[86]),
  .la_data_out_87(la_data_out[87]),
  .la_data_out_88(la_data_out[88]),
  .la_data_out_89(la_data_out[89]),
  .la_data_out_90(la_data_out[90]),
  .la_data_out_91(la_data_out[91]),
  .la_data_out_92(la_data_out[92]),
  .la_data_out_93(la_data_out[93]),
  .la_data_out_94(la_data_out[94]),
  .la_data_out_95(la_data_out[95]),
  .la_data_out_96(la_data_out[96]),
  .la_data_out_97(la_data_out[97]),
  .la_data_out_98(la_data_out[98]),
  .la_data_out_99(la_data_out[99]),
  .la_data_out_100(la_data_out[100]),
  .la_data_out_101(la_data_out[101]),
  .la_data_out_102(la_data_out[102]),
  .la_data_out_103(la_data_out[103]),
  .la_data_out_104(la_data_out[104]),
  .la_data_out_105(la_data_out[105]),
  .la_data_out_106(la_data_out[106]),
  .la_data_out_107(la_data_out[107]),
  .la_data_out_108(la_data_out[108]),
  .la_data_out_109(la_data_out[109]),
  .la_data_out_110(la_data_out[110]),
  .la_data_out_111(la_data_out[111]),
  .la_data_out_112(la_data_out[112]),
  .la_data_out_113(la_data_out[113]),
  .la_data_out_114(la_data_out[114]),
  .la_data_out_115(la_data_out[115]),
  .la_data_out_116(la_data_out[116]),
  .la_data_out_117(la_data_out[117]),
  .la_data_out_118(la_data_out[118]),
  .la_data_out_119(la_data_out[119]),
  .la_data_out_120(la_data_out[120]),
  .la_data_out_121(la_data_out[121]),
  .la_data_out_122(la_data_out[122]),
  .la_data_out_123(la_data_out[123]),
  .la_data_out_124(la_data_out[124]),
  .la_data_out_125(la_data_out[125]),
  .la_data_out_126(la_data_out[126]),
  .la_data_out_127(la_data_out[127]),
  .la_oenb_0(la_oenb[0]),
  .la_oenb_1(la_oenb[1]),
  .la_oenb_2(la_oenb[2]),
  .la_oenb_3(la_oenb[3]),
  .la_oenb_4(la_oenb[4]),
  .la_oenb_5(la_oenb[5]),
  .la_oenb_6(la_oenb[6]),
  .la_oenb_7(la_oenb[7]),
  .la_oenb_8(la_oenb[8]),
  .la_oenb_9(la_oenb[9]),
  .la_oenb_10(la_oenb[10]),
  .la_oenb_11(la_oenb[11]),
  .la_oenb_12(la_oenb[12]),
  .la_oenb_13(la_oenb[13]),
  .la_oenb_14(la_oenb[14]),
  .la_oenb_15(la_oenb[15]),
  .la_oenb_16(la_oenb[16]),
  .la_oenb_17(la_oenb[17]),
  .la_oenb_18(la_oenb[18]),
  .la_oenb_19(la_oenb[19]),
  .la_oenb_20(la_oenb[20]),
  .la_oenb_21(la_oenb[21]),
  .la_oenb_22(la_oenb[22]),
  .la_oenb_23(la_oenb[23]),
  .la_oenb_24(la_oenb[24]),
  .la_oenb_25(la_oenb[25]),
  .la_oenb_26(la_oenb[26]),
  .la_oenb_27(la_oenb[27]),
  .la_oenb_28(la_oenb[28]),
  .la_oenb_29(la_oenb[29]),
  .la_oenb_30(la_oenb[30]),
  .la_oenb_31(la_oenb[31]),
  .la_oenb_32(la_oenb[32]),
  .la_oenb_33(la_oenb[33]),
  .la_oenb_34(la_oenb[34]),
  .la_oenb_35(la_oenb[35]),
  .la_oenb_36(la_oenb[36]),
  .la_oenb_37(la_oenb[37]),
  .la_oenb_38(la_oenb[38]),
  .la_oenb_39(la_oenb[39]),
  .la_oenb_40(la_oenb[40]),
  .la_oenb_41(la_oenb[41]),
  .la_oenb_42(la_oenb[42]),
  .la_oenb_43(la_oenb[43]),
  .la_oenb_44(la_oenb[44]),
  .la_oenb_45(la_oenb[45]),
  .la_oenb_46(la_oenb[46]),
  .la_oenb_47(la_oenb[47]),
  .la_oenb_48(la_oenb[48]),
  .la_oenb_49(la_oenb[49]),
  .la_oenb_50(la_oenb[50]),
  .la_oenb_51(la_oenb[51]),
  .la_oenb_52(la_oenb[52]),
  .la_oenb_53(la_oenb[53]),
  .la_oenb_54(la_oenb[54]),
  .la_oenb_55(la_oenb[55]),
  .la_oenb_56(la_oenb[56]),
  .la_oenb_57(la_oenb[57]),
  .la_oenb_58(la_oenb[58]),
  .la_oenb_59(la_oenb[59]),
  .la_oenb_60(la_oenb[60]),
  .la_oenb_61(la_oenb[61]),
  .la_oenb_62(la_oenb[62]),
  .la_oenb_63(la_oenb[63]),
  .la_oenb_64(la_oenb[64]),
  .la_oenb_65(la_oenb[65]),
  .la_oenb_66(la_oenb[66]),
  .la_oenb_67(la_oenb[67]),
  .la_oenb_68(la_oenb[68]),
  .la_oenb_69(la_oenb[69]),
  .la_oenb_70(la_oenb[70]),
  .la_oenb_71(la_oenb[71]),
  .la_oenb_72(la_oenb[72]),
  .la_oenb_73(la_oenb[73]),
  .la_oenb_74(la_oenb[74]),
  .la_oenb_75(la_oenb[75]),
  .la_oenb_76(la_oenb[76]),
  .la_oenb_77(la_oenb[77]),
  .la_oenb_78(la_oenb[78]),
  .la_oenb_79(la_oenb[79]),
  .la_oenb_80(la_oenb[80]),
  .la_oenb_81(la_oenb[81]),
  .la_oenb_82(la_oenb[82]),
  .la_oenb_83(la_oenb[83]),
  .la_oenb_84(la_oenb[84]),
  .la_oenb_85(la_oenb[85]),
  .la_oenb_86(la_oenb[86]),
  .la_oenb_87(la_oenb[87]),
  .la_oenb_88(la_oenb[88]),
  .la_oenb_89(la_oenb[89]),
  .la_oenb_90(la_oenb[90]),
  .la_oenb_91(la_oenb[91]),
  .la_oenb_92(la_oenb[92]),
  .la_oenb_93(la_oenb[93]),
  .la_oenb_94(la_oenb[94]),
  .la_oenb_95(la_oenb[95]),
  .la_oenb_96(la_oenb[96]),
  .la_oenb_97(la_oenb[97]),
  .la_oenb_98(la_oenb[98]),
  .la_oenb_99(la_oenb[99]),
  .la_oenb_100(la_oenb[100]),
  .la_oenb_101(la_oenb[101]),
  .la_oenb_102(la_oenb[102]),
  .la_oenb_103(la_oenb[103]),
  .la_oenb_104(la_oenb[104]),
  .la_oenb_105(la_oenb[105]),
  .la_oenb_106(la_oenb[106]),
  .la_oenb_107(la_oenb[107]),
  .la_oenb_108(la_oenb[108]),
  .la_oenb_109(la_oenb[109]),
  .la_oenb_110(la_oenb[110]),
  .la_oenb_111(la_oenb[111]),
  .la_oenb_112(la_oenb[112]),
  .la_oenb_113(la_oenb[113]),
  .la_oenb_114(la_oenb[114]),
  .la_oenb_115(la_oenb[115]),
  .la_oenb_116(la_oenb[116]),
  .la_oenb_117(la_oenb[117]),
  .la_oenb_118(la_oenb[118]),
  .la_oenb_119(la_oenb[119]),
  .la_oenb_120(la_oenb[120]),
  .la_oenb_121(la_oenb[121]),
  .la_oenb_122(la_oenb[122]),
  .la_oenb_123(la_oenb[123]),
  .la_oenb_124(la_oenb[124]),
  .la_oenb_125(la_oenb[125]),
  .la_oenb_126(la_oenb[126]),
  .la_oenb_127(la_oenb[127]),
  .io_in_0(io_in[0]),
  .io_in_1(io_in[1]),
  .io_in_2(io_in[2]),
  .io_in_3(io_in[3]),
  .io_in_4(io_in[4]),
  .io_in_5(io_in[5]),
  .io_in_6(io_in[6]),
  .io_in_7(io_in[7]),
  .io_in_8(io_in[8]),
  .io_in_9(io_in[9]),
  .io_in_10(io_in[10]),
  .io_in_11(io_in[11]),
  .io_in_12(io_in[12]),
  .io_in_13(io_in[13]),
  .io_in_14(io_in[14]),
  .io_in_15(io_in[15]),
  .io_in_16(io_in[16]),
  .io_in_17(io_in[17]),
  .io_in_18(io_in[18]),
  .io_in_19(io_in[19]),
  .io_in_20(io_in[20]),
  .io_in_21(io_in[21]),
  .io_in_22(io_in[22]),
  .io_in_23(io_in[23]),
  .io_in_24(io_in[24]),
  .io_in_25(io_in[25]),
  .io_in_26(io_in[26]),
  .io_in_27(io_in[27]),
  .io_in_28(io_in[28]),
  .io_in_29(io_in[29]),
  .io_in_30(io_in[30]),
  .io_in_31(io_in[31]),
  .io_in_32(io_in[32]),
  .io_in_33(io_in[33]),
  .io_in_34(io_in[34]),
  .io_in_35(io_in[35]),
  .io_in_36(io_in[36]),
  .io_in_37(io_in[37]),
  .io_out_0(io_out[0]),
  .io_out_1(io_out[1]),
  .io_out_2(io_out[2]),
  .io_out_3(io_out[3]),
  .io_out_4(io_out[4]),
  .io_out_5(io_out[5]),
  .io_out_6(io_out[6]),
  .io_out_7(io_out[7]),
  .io_out_8(io_out[8]),
  .io_out_9(io_out[9]),
  .io_out_10(io_out[10]),
  .io_out_11(io_out[11]),
  .io_out_12(io_out[12]),
  .io_out_13(io_out[13]),
  .io_out_14(io_out[14]),
  .io_out_15(io_out[15]),
  .io_out_16(io_out[16]),
  .io_out_17(io_out[17]),
  .io_out_18(io_out[18]),
  .io_out_19(io_out[19]),
  .io_out_20(io_out[20]),
  .io_out_21(io_out[21]),
  .io_out_22(io_out[22]),
  .io_out_23(io_out[23]),
  .io_out_24(io_out[24]),
  .io_out_25(io_out[25]),
  .io_out_26(io_out[26]),
  .io_out_27(io_out[27]),
  .io_out_28(io_out[28]),
  .io_out_29(io_out[29]),
  .io_out_30(io_out[30]),
  .io_out_31(io_out[31]),
  .io_out_32(io_out[32]),
  .io_out_33(io_out[33]),
  .io_out_34(io_out[34]),
  .io_out_35(io_out[35]),
  .io_out_36(io_out[36]),
  .io_out_37(io_out[37]),
  .io_oeb_0(io_oeb[0]),
  .io_oeb_1(io_oeb[1]),
  .io_oeb_2(io_oeb[2]),
  .io_oeb_3(io_oeb[3]),
  .io_oeb_4(io_oeb[4]),
  .io_oeb_5(io_oeb[5]),
  .io_oeb_6(io_oeb[6]),
  .io_oeb_7(io_oeb[7]),
  .io_oeb_8(io_oeb[8]),
  .io_oeb_9(io_oeb[9]),
  .io_oeb_10(io_oeb[10]),
  .io_oeb_11(io_oeb[11]),
  .io_oeb_12(io_oeb[12]),
  .io_oeb_13(io_oeb[13]),
  .io_oeb_14(io_oeb[14]),
  .io_oeb_15(io_oeb[15]),
  .io_oeb_16(io_oeb[16]),
  .io_oeb_17(io_oeb[17]),
  .io_oeb_18(io_oeb[18]),
  .io_oeb_19(io_oeb[19]),
  .io_oeb_20(io_oeb[20]),
  .io_oeb_21(io_oeb[21]),
  .io_oeb_22(io_oeb[22]),
  .io_oeb_23(io_oeb[23]),
  .io_oeb_24(io_oeb[24]),
  .io_oeb_25(io_oeb[25]),
  .io_oeb_26(io_oeb[26]),
  .io_oeb_27(io_oeb[27]),
  .io_oeb_28(io_oeb[28]),
  .io_oeb_29(io_oeb[29]),
  .io_oeb_30(io_oeb[30]),
  .io_oeb_31(io_oeb[31]),
  .io_oeb_32(io_oeb[32]),
  .io_oeb_33(io_oeb[33]),
  .io_oeb_34(io_oeb[34]),
  .io_oeb_35(io_oeb[35]),
  .io_oeb_36(io_oeb[36]),
  .io_oeb_37(io_oeb[37]),
  .irq_0(irq[0]),
  .irq_1(irq[1]),
  .irq_2(irq[2])
 );

endmodule

