// /home/shc/Research/RISC-V/freedom/builds/marmotcaravel/xip.hex
case (address)
  11'h000: out <= 32'hf1402573;
  11'h001: out <= 32'h00000597;
  11'h002: out <= 32'h01058593;
  11'h003: out <= 32'h200002b7;
  11'h004: out <= 32'h00028067;
  11'h005: out <= 32'hedfe0dd0;
  11'h006: out <= 32'h1a0f0000;
  11'h007: out <= 32'h38000000;
  11'h008: out <= 32'h940d0000;
  11'h009: out <= 32'h28000000;
  11'h00a: out <= 32'h11000000;
  11'h00b: out <= 32'h10000000;
  11'h00c: out <= 32'h00000000;
  11'h00d: out <= 32'h86010000;
  11'h00e: out <= 32'h5c0d0000;
  11'h00f: out <= 32'h00000000;
  11'h010: out <= 32'h00000000;
  11'h011: out <= 32'h00000000;
  11'h012: out <= 32'h00000000;
  11'h013: out <= 32'h01000000;
  11'h014: out <= 32'h00000000;
  11'h015: out <= 32'h03000000;
  11'h016: out <= 32'h04000000;
  11'h017: out <= 32'h00000000;
  11'h018: out <= 32'h01000000;
  11'h019: out <= 32'h03000000;
  11'h01a: out <= 32'h04000000;
  11'h01b: out <= 32'h0f000000;
  11'h01c: out <= 32'h01000000;
  11'h01d: out <= 32'h03000000;
  11'h01e: out <= 32'h21000000;
  11'h01f: out <= 32'h1b000000;
  11'h020: out <= 32'h65657266;
  11'h021: out <= 32'h70696863;
  11'h022: out <= 32'h6f722c73;
  11'h023: out <= 32'h74656b63;
  11'h024: out <= 32'h70696863;
  11'h025: out <= 32'h6b6e752d;
  11'h026: out <= 32'h6e776f6e;
  11'h027: out <= 32'h7665642d;
  11'h028: out <= 32'h00000000;
  11'h029: out <= 32'h03000000;
  11'h02a: out <= 32'h1d000000;
  11'h02b: out <= 32'h26000000;
  11'h02c: out <= 32'h65657266;
  11'h02d: out <= 32'h70696863;
  11'h02e: out <= 32'h6f722c73;
  11'h02f: out <= 32'h74656b63;
  11'h030: out <= 32'h70696863;
  11'h031: out <= 32'h6b6e752d;
  11'h032: out <= 32'h6e776f6e;
  11'h033: out <= 32'h00000000;
  11'h034: out <= 32'h01000000;
  11'h035: out <= 32'h61696c61;
  11'h036: out <= 32'h00736573;
  11'h037: out <= 32'h03000000;
  11'h038: out <= 32'h15000000;
  11'h039: out <= 32'h2c000000;
  11'h03a: out <= 32'h636f732f;
  11'h03b: out <= 32'h7265732f;
  11'h03c: out <= 32'h406c6169;
  11'h03d: out <= 32'h31303031;
  11'h03e: out <= 32'h30303033;
  11'h03f: out <= 32'h00000000;
  11'h040: out <= 32'h03000000;
  11'h041: out <= 32'h15000000;
  11'h042: out <= 32'h34000000;
  11'h043: out <= 32'h636f732f;
  11'h044: out <= 32'h7265732f;
  11'h045: out <= 32'h406c6169;
  11'h046: out <= 32'h32303031;
  11'h047: out <= 32'h30303033;
  11'h048: out <= 32'h00000000;
  11'h049: out <= 32'h03000000;
  11'h04a: out <= 32'h15000000;
  11'h04b: out <= 32'h3c000000;
  11'h04c: out <= 32'h636f732f;
  11'h04d: out <= 32'h7265732f;
  11'h04e: out <= 32'h406c6169;
  11'h04f: out <= 32'h33303031;
  11'h050: out <= 32'h30303033;
  11'h051: out <= 32'h00000000;
  11'h052: out <= 32'h03000000;
  11'h053: out <= 32'h15000000;
  11'h054: out <= 32'h44000000;
  11'h055: out <= 32'h636f732f;
  11'h056: out <= 32'h7265732f;
  11'h057: out <= 32'h406c6169;
  11'h058: out <= 32'h34303031;
  11'h059: out <= 32'h30303033;
  11'h05a: out <= 32'h00000000;
  11'h05b: out <= 32'h03000000;
  11'h05c: out <= 32'h15000000;
  11'h05d: out <= 32'h4c000000;
  11'h05e: out <= 32'h636f732f;
  11'h05f: out <= 32'h7265732f;
  11'h060: out <= 32'h406c6169;
  11'h061: out <= 32'h35303031;
  11'h062: out <= 32'h30303033;
  11'h063: out <= 32'h00000000;
  11'h064: out <= 32'h02000000;
  11'h065: out <= 32'h01000000;
  11'h066: out <= 32'h73757063;
  11'h067: out <= 32'h00000000;
  11'h068: out <= 32'h03000000;
  11'h069: out <= 32'h04000000;
  11'h06a: out <= 32'h00000000;
  11'h06b: out <= 32'h01000000;
  11'h06c: out <= 32'h03000000;
  11'h06d: out <= 32'h04000000;
  11'h06e: out <= 32'h0f000000;
  11'h06f: out <= 32'h00000000;
  11'h070: out <= 32'h01000000;
  11'h071: out <= 32'h40757063;
  11'h072: out <= 32'h00000030;
  11'h073: out <= 32'h03000000;
  11'h074: out <= 32'h04000000;
  11'h075: out <= 32'h54000000;
  11'h076: out <= 32'h00000000;
  11'h077: out <= 32'h03000000;
  11'h078: out <= 32'h15000000;
  11'h079: out <= 32'h1b000000;
  11'h07a: out <= 32'h69666973;
  11'h07b: out <= 32'h722c6576;
  11'h07c: out <= 32'h656b636f;
  11'h07d: out <= 32'h72003074;
  11'h07e: out <= 32'h76637369;
  11'h07f: out <= 32'h00000000;
  11'h080: out <= 32'h03000000;
  11'h081: out <= 32'h04000000;
  11'h082: out <= 32'h64000000;
  11'h083: out <= 32'h00757063;
  11'h084: out <= 32'h03000000;
  11'h085: out <= 32'h04000000;
  11'h086: out <= 32'h70000000;
  11'h087: out <= 32'h40000000;
  11'h088: out <= 32'h03000000;
  11'h089: out <= 32'h04000000;
  11'h08a: out <= 32'h83000000;
  11'h08b: out <= 32'h80000000;
  11'h08c: out <= 32'h03000000;
  11'h08d: out <= 32'h04000000;
  11'h08e: out <= 32'h90000000;
  11'h08f: out <= 32'h00400000;
  11'h090: out <= 32'h03000000;
  11'h091: out <= 32'h04000000;
  11'h092: out <= 32'h9d000000;
  11'h093: out <= 32'h00000000;
  11'h094: out <= 32'h03000000;
  11'h095: out <= 32'h09000000;
  11'h096: out <= 32'ha1000000;
  11'h097: out <= 32'h32337672;
  11'h098: out <= 32'h63616d69;
  11'h099: out <= 32'h00000000;
  11'h09a: out <= 32'h03000000;
  11'h09b: out <= 32'h04000000;
  11'h09c: out <= 32'hab000000;
  11'h09d: out <= 32'h01000000;
  11'h09e: out <= 32'h03000000;
  11'h09f: out <= 32'h04000000;
  11'h0a0: out <= 32'hb7000000;
  11'h0a1: out <= 32'h02000000;
  11'h0a2: out <= 32'h03000000;
  11'h0a3: out <= 32'h05000000;
  11'h0a4: out <= 32'hc3000000;
  11'h0a5: out <= 32'h79616b6f;
  11'h0a6: out <= 32'h00000000;
  11'h0a7: out <= 32'h03000000;
  11'h0a8: out <= 32'h04000000;
  11'h0a9: out <= 32'hca000000;
  11'h0aa: out <= 32'h00800000;
  11'h0ab: out <= 32'h01000000;
  11'h0ac: out <= 32'h65746e69;
  11'h0ad: out <= 32'h70757272;
  11'h0ae: out <= 32'h6f632d74;
  11'h0af: out <= 32'h6f72746e;
  11'h0b0: out <= 32'h72656c6c;
  11'h0b1: out <= 32'h00000000;
  11'h0b2: out <= 32'h03000000;
  11'h0b3: out <= 32'h04000000;
  11'h0b4: out <= 32'hdd000000;
  11'h0b5: out <= 32'h01000000;
  11'h0b6: out <= 32'h03000000;
  11'h0b7: out <= 32'h0f000000;
  11'h0b8: out <= 32'h1b000000;
  11'h0b9: out <= 32'h63736972;
  11'h0ba: out <= 32'h70632c76;
  11'h0bb: out <= 32'h6e692d75;
  11'h0bc: out <= 32'h00006374;
  11'h0bd: out <= 32'h03000000;
  11'h0be: out <= 32'h00000000;
  11'h0bf: out <= 32'hee000000;
  11'h0c0: out <= 32'h03000000;
  11'h0c1: out <= 32'h04000000;
  11'h0c2: out <= 32'h03010000;
  11'h0c3: out <= 32'h04000000;
  11'h0c4: out <= 32'h02000000;
  11'h0c5: out <= 32'h02000000;
  11'h0c6: out <= 32'h02000000;
  11'h0c7: out <= 32'h01000000;
  11'h0c8: out <= 32'h00636f73;
  11'h0c9: out <= 32'h03000000;
  11'h0ca: out <= 32'h04000000;
  11'h0cb: out <= 32'h00000000;
  11'h0cc: out <= 32'h01000000;
  11'h0cd: out <= 32'h03000000;
  11'h0ce: out <= 32'h04000000;
  11'h0cf: out <= 32'h0f000000;
  11'h0d0: out <= 32'h01000000;
  11'h0d1: out <= 32'h03000000;
  11'h0d2: out <= 32'h2c000000;
  11'h0d3: out <= 32'h1b000000;
  11'h0d4: out <= 32'h65657266;
  11'h0d5: out <= 32'h70696863;
  11'h0d6: out <= 32'h6f722c73;
  11'h0d7: out <= 32'h74656b63;
  11'h0d8: out <= 32'h70696863;
  11'h0d9: out <= 32'h6b6e752d;
  11'h0da: out <= 32'h6e776f6e;
  11'h0db: out <= 32'h636f732d;
  11'h0dc: out <= 32'h6d697300;
  11'h0dd: out <= 32'h2d656c70;
  11'h0de: out <= 32'h00737562;
  11'h0df: out <= 32'h03000000;
  11'h0e0: out <= 32'h00000000;
  11'h0e1: out <= 32'h0b010000;
  11'h0e2: out <= 32'h01000000;
  11'h0e3: out <= 32'h406e6f61;
  11'h0e4: out <= 32'h30303031;
  11'h0e5: out <= 32'h30303030;
  11'h0e6: out <= 32'h00000000;
  11'h0e7: out <= 32'h03000000;
  11'h0e8: out <= 32'h0c000000;
  11'h0e9: out <= 32'h1b000000;
  11'h0ea: out <= 32'h69666973;
  11'h0eb: out <= 32'h612c6576;
  11'h0ec: out <= 32'h00306e6f;
  11'h0ed: out <= 32'h03000000;
  11'h0ee: out <= 32'h04000000;
  11'h0ef: out <= 32'h12010000;
  11'h0f0: out <= 32'h03000000;
  11'h0f1: out <= 32'h03000000;
  11'h0f2: out <= 32'h08000000;
  11'h0f3: out <= 32'h23010000;
  11'h0f4: out <= 32'h01000000;
  11'h0f5: out <= 32'h02000000;
  11'h0f6: out <= 32'h03000000;
  11'h0f7: out <= 32'h08000000;
  11'h0f8: out <= 32'h9d000000;
  11'h0f9: out <= 32'h00000010;
  11'h0fa: out <= 32'h00100000;
  11'h0fb: out <= 32'h03000000;
  11'h0fc: out <= 32'h08000000;
  11'h0fd: out <= 32'h2e010000;
  11'h0fe: out <= 32'h746e6f63;
  11'h0ff: out <= 32'h006c6f72;
  11'h100: out <= 32'h02000000;
  11'h101: out <= 32'h01000000;
  11'h102: out <= 32'h6e696c63;
  11'h103: out <= 32'h30324074;
  11'h104: out <= 32'h30303030;
  11'h105: out <= 32'h00000030;
  11'h106: out <= 32'h03000000;
  11'h107: out <= 32'h0d000000;
  11'h108: out <= 32'h1b000000;
  11'h109: out <= 32'h63736972;
  11'h10a: out <= 32'h6c632c76;
  11'h10b: out <= 32'h30746e69;
  11'h10c: out <= 32'h00000000;
  11'h10d: out <= 32'h03000000;
  11'h10e: out <= 32'h10000000;
  11'h10f: out <= 32'h38010000;
  11'h110: out <= 32'h04000000;
  11'h111: out <= 32'h03000000;
  11'h112: out <= 32'h04000000;
  11'h113: out <= 32'h07000000;
  11'h114: out <= 32'h03000000;
  11'h115: out <= 32'h08000000;
  11'h116: out <= 32'h9d000000;
  11'h117: out <= 32'h00000002;
  11'h118: out <= 32'h00000100;
  11'h119: out <= 32'h03000000;
  11'h11a: out <= 32'h08000000;
  11'h11b: out <= 32'h2e010000;
  11'h11c: out <= 32'h746e6f63;
  11'h11d: out <= 32'h006c6f72;
  11'h11e: out <= 32'h02000000;
  11'h11f: out <= 32'h01000000;
  11'h120: out <= 32'h75626564;
  11'h121: out <= 32'h6f632d67;
  11'h122: out <= 32'h6f72746e;
  11'h123: out <= 32'h72656c6c;
  11'h124: out <= 32'h00003040;
  11'h125: out <= 32'h03000000;
  11'h126: out <= 32'h21000000;
  11'h127: out <= 32'h1b000000;
  11'h128: out <= 32'h69666973;
  11'h129: out <= 32'h642c6576;
  11'h12a: out <= 32'h67756265;
  11'h12b: out <= 32'h3331302d;
  11'h12c: out <= 32'h73697200;
  11'h12d: out <= 32'h642c7663;
  11'h12e: out <= 32'h67756265;
  11'h12f: out <= 32'h3331302d;
  11'h130: out <= 32'h00000000;
  11'h131: out <= 32'h03000000;
  11'h132: out <= 32'h08000000;
  11'h133: out <= 32'h38010000;
  11'h134: out <= 32'h04000000;
  11'h135: out <= 32'hffff0000;
  11'h136: out <= 32'h03000000;
  11'h137: out <= 32'h08000000;
  11'h138: out <= 32'h9d000000;
  11'h139: out <= 32'h00000000;
  11'h13a: out <= 32'h00100000;
  11'h13b: out <= 32'h03000000;
  11'h13c: out <= 32'h08000000;
  11'h13d: out <= 32'h2e010000;
  11'h13e: out <= 32'h746e6f63;
  11'h13f: out <= 32'h006c6f72;
  11'h140: out <= 32'h02000000;
  11'h141: out <= 32'h01000000;
  11'h142: out <= 32'h6d697464;
  11'h143: out <= 32'h30303840;
  11'h144: out <= 32'h30303030;
  11'h145: out <= 32'h00000030;
  11'h146: out <= 32'h03000000;
  11'h147: out <= 32'h0d000000;
  11'h148: out <= 32'h1b000000;
  11'h149: out <= 32'h69666973;
  11'h14a: out <= 32'h642c6576;
  11'h14b: out <= 32'h306d6974;
  11'h14c: out <= 32'h00000000;
  11'h14d: out <= 32'h03000000;
  11'h14e: out <= 32'h08000000;
  11'h14f: out <= 32'h9d000000;
  11'h150: out <= 32'h00000080;
  11'h151: out <= 32'h00400000;
  11'h152: out <= 32'h03000000;
  11'h153: out <= 32'h04000000;
  11'h154: out <= 32'h2e010000;
  11'h155: out <= 32'h006d656d;
  11'h156: out <= 32'h03000000;
  11'h157: out <= 32'h04000000;
  11'h158: out <= 32'h03010000;
  11'h159: out <= 32'h01000000;
  11'h15a: out <= 32'h02000000;
  11'h15b: out <= 32'h01000000;
  11'h15c: out <= 32'h6f727265;
  11'h15d: out <= 32'h65642d72;
  11'h15e: out <= 32'h65636976;
  11'h15f: out <= 32'h30303340;
  11'h160: out <= 32'h00000030;
  11'h161: out <= 32'h03000000;
  11'h162: out <= 32'h0e000000;
  11'h163: out <= 32'h1b000000;
  11'h164: out <= 32'h69666973;
  11'h165: out <= 32'h652c6576;
  11'h166: out <= 32'h726f7272;
  11'h167: out <= 32'h00000030;
  11'h168: out <= 32'h03000000;
  11'h169: out <= 32'h08000000;
  11'h16a: out <= 32'h9d000000;
  11'h16b: out <= 32'h00300000;
  11'h16c: out <= 32'h00100000;
  11'h16d: out <= 32'h02000000;
  11'h16e: out <= 32'h01000000;
  11'h16f: out <= 32'h6f697067;
  11'h170: out <= 32'h30303140;
  11'h171: out <= 32'h30303231;
  11'h172: out <= 32'h00000030;
  11'h173: out <= 32'h03000000;
  11'h174: out <= 32'h04000000;
  11'h175: out <= 32'h4c010000;
  11'h176: out <= 32'h02000000;
  11'h177: out <= 32'h03000000;
  11'h178: out <= 32'h04000000;
  11'h179: out <= 32'hdd000000;
  11'h17a: out <= 32'h02000000;
  11'h17b: out <= 32'h03000000;
  11'h17c: out <= 32'h0d000000;
  11'h17d: out <= 32'h1b000000;
  11'h17e: out <= 32'h69666973;
  11'h17f: out <= 32'h672c6576;
  11'h180: out <= 32'h306f6970;
  11'h181: out <= 32'h00000000;
  11'h182: out <= 32'h03000000;
  11'h183: out <= 32'h00000000;
  11'h184: out <= 32'h58010000;
  11'h185: out <= 32'h03000000;
  11'h186: out <= 32'h00000000;
  11'h187: out <= 32'hee000000;
  11'h188: out <= 32'h03000000;
  11'h189: out <= 32'h04000000;
  11'h18a: out <= 32'h12010000;
  11'h18b: out <= 32'h03000000;
  11'h18c: out <= 32'h03000000;
  11'h18d: out <= 32'h80000000;
  11'h18e: out <= 32'h23010000;
  11'h18f: out <= 32'h0b000000;
  11'h190: out <= 32'h0c000000;
  11'h191: out <= 32'h0d000000;
  11'h192: out <= 32'h0e000000;
  11'h193: out <= 32'h0f000000;
  11'h194: out <= 32'h10000000;
  11'h195: out <= 32'h11000000;
  11'h196: out <= 32'h12000000;
  11'h197: out <= 32'h13000000;
  11'h198: out <= 32'h14000000;
  11'h199: out <= 32'h15000000;
  11'h19a: out <= 32'h16000000;
  11'h19b: out <= 32'h17000000;
  11'h19c: out <= 32'h18000000;
  11'h19d: out <= 32'h19000000;
  11'h19e: out <= 32'h1a000000;
  11'h19f: out <= 32'h1b000000;
  11'h1a0: out <= 32'h1c000000;
  11'h1a1: out <= 32'h1d000000;
  11'h1a2: out <= 32'h1e000000;
  11'h1a3: out <= 32'h1f000000;
  11'h1a4: out <= 32'h20000000;
  11'h1a5: out <= 32'h21000000;
  11'h1a6: out <= 32'h22000000;
  11'h1a7: out <= 32'h23000000;
  11'h1a8: out <= 32'h24000000;
  11'h1a9: out <= 32'h25000000;
  11'h1aa: out <= 32'h26000000;
  11'h1ab: out <= 32'h27000000;
  11'h1ac: out <= 32'h28000000;
  11'h1ad: out <= 32'h29000000;
  11'h1ae: out <= 32'h2a000000;
  11'h1af: out <= 32'h03000000;
  11'h1b0: out <= 32'h08000000;
  11'h1b1: out <= 32'h9d000000;
  11'h1b2: out <= 32'h00200110;
  11'h1b3: out <= 32'h00100000;
  11'h1b4: out <= 32'h03000000;
  11'h1b5: out <= 32'h08000000;
  11'h1b6: out <= 32'h2e010000;
  11'h1b7: out <= 32'h746e6f63;
  11'h1b8: out <= 32'h006c6f72;
  11'h1b9: out <= 32'h02000000;
  11'h1ba: out <= 32'h01000000;
  11'h1bb: out <= 32'h40633269;
  11'h1bc: out <= 32'h31303031;
  11'h1bd: out <= 32'h30303036;
  11'h1be: out <= 32'h00000000;
  11'h1bf: out <= 32'h03000000;
  11'h1c0: out <= 32'h0c000000;
  11'h1c1: out <= 32'h1b000000;
  11'h1c2: out <= 32'h69666973;
  11'h1c3: out <= 32'h692c6576;
  11'h1c4: out <= 32'h00306332;
  11'h1c5: out <= 32'h03000000;
  11'h1c6: out <= 32'h04000000;
  11'h1c7: out <= 32'h12010000;
  11'h1c8: out <= 32'h03000000;
  11'h1c9: out <= 32'h03000000;
  11'h1ca: out <= 32'h04000000;
  11'h1cb: out <= 32'h23010000;
  11'h1cc: out <= 32'h2b000000;
  11'h1cd: out <= 32'h03000000;
  11'h1ce: out <= 32'h08000000;
  11'h1cf: out <= 32'h9d000000;
  11'h1d0: out <= 32'h00600110;
  11'h1d1: out <= 32'h00100000;
  11'h1d2: out <= 32'h03000000;
  11'h1d3: out <= 32'h08000000;
  11'h1d4: out <= 32'h2e010000;
  11'h1d5: out <= 32'h746e6f63;
  11'h1d6: out <= 32'h006c6f72;
  11'h1d7: out <= 32'h02000000;
  11'h1d8: out <= 32'h01000000;
  11'h1d9: out <= 32'h40633269;
  11'h1da: out <= 32'h32303031;
  11'h1db: out <= 32'h30303036;
  11'h1dc: out <= 32'h00000000;
  11'h1dd: out <= 32'h03000000;
  11'h1de: out <= 32'h0c000000;
  11'h1df: out <= 32'h1b000000;
  11'h1e0: out <= 32'h69666973;
  11'h1e1: out <= 32'h692c6576;
  11'h1e2: out <= 32'h00306332;
  11'h1e3: out <= 32'h03000000;
  11'h1e4: out <= 32'h04000000;
  11'h1e5: out <= 32'h12010000;
  11'h1e6: out <= 32'h03000000;
  11'h1e7: out <= 32'h03000000;
  11'h1e8: out <= 32'h04000000;
  11'h1e9: out <= 32'h23010000;
  11'h1ea: out <= 32'h2c000000;
  11'h1eb: out <= 32'h03000000;
  11'h1ec: out <= 32'h08000000;
  11'h1ed: out <= 32'h9d000000;
  11'h1ee: out <= 32'h00600210;
  11'h1ef: out <= 32'h00100000;
  11'h1f0: out <= 32'h03000000;
  11'h1f1: out <= 32'h08000000;
  11'h1f2: out <= 32'h2e010000;
  11'h1f3: out <= 32'h746e6f63;
  11'h1f4: out <= 32'h006c6f72;
  11'h1f5: out <= 32'h02000000;
  11'h1f6: out <= 32'h01000000;
  11'h1f7: out <= 32'h65746e69;
  11'h1f8: out <= 32'h70757272;
  11'h1f9: out <= 32'h6f632d74;
  11'h1fa: out <= 32'h6f72746e;
  11'h1fb: out <= 32'h72656c6c;
  11'h1fc: out <= 32'h30306340;
  11'h1fd: out <= 32'h30303030;
  11'h1fe: out <= 32'h00000000;
  11'h1ff: out <= 32'h03000000;
  11'h200: out <= 32'h04000000;
  11'h201: out <= 32'hdd000000;
  11'h202: out <= 32'h01000000;
  11'h203: out <= 32'h03000000;
  11'h204: out <= 32'h0c000000;
  11'h205: out <= 32'h1b000000;
  11'h206: out <= 32'h63736972;
  11'h207: out <= 32'h6c702c76;
  11'h208: out <= 32'h00306369;
  11'h209: out <= 32'h03000000;
  11'h20a: out <= 32'h00000000;
  11'h20b: out <= 32'hee000000;
  11'h20c: out <= 32'h03000000;
  11'h20d: out <= 32'h08000000;
  11'h20e: out <= 32'h38010000;
  11'h20f: out <= 32'h04000000;
  11'h210: out <= 32'h0b000000;
  11'h211: out <= 32'h03000000;
  11'h212: out <= 32'h08000000;
  11'h213: out <= 32'h9d000000;
  11'h214: out <= 32'h0000000c;
  11'h215: out <= 32'h00000004;
  11'h216: out <= 32'h03000000;
  11'h217: out <= 32'h08000000;
  11'h218: out <= 32'h2e010000;
  11'h219: out <= 32'h746e6f63;
  11'h21a: out <= 32'h006c6f72;
  11'h21b: out <= 32'h03000000;
  11'h21c: out <= 32'h04000000;
  11'h21d: out <= 32'h68010000;
  11'h21e: out <= 32'h07000000;
  11'h21f: out <= 32'h03000000;
  11'h220: out <= 32'h04000000;
  11'h221: out <= 32'h7b010000;
  11'h222: out <= 32'h2c000000;
  11'h223: out <= 32'h03000000;
  11'h224: out <= 32'h04000000;
  11'h225: out <= 32'h03010000;
  11'h226: out <= 32'h03000000;
  11'h227: out <= 32'h02000000;
  11'h228: out <= 32'h01000000;
  11'h229: out <= 32'h6d697469;
  11'h22a: out <= 32'h30303840;
  11'h22b: out <= 32'h30303030;
  11'h22c: out <= 32'h00000000;
  11'h22d: out <= 32'h03000000;
  11'h22e: out <= 32'h0d000000;
  11'h22f: out <= 32'h1b000000;
  11'h230: out <= 32'h69666973;
  11'h231: out <= 32'h692c6576;
  11'h232: out <= 32'h306d6974;
  11'h233: out <= 32'h00000000;
  11'h234: out <= 32'h03000000;
  11'h235: out <= 32'h08000000;
  11'h236: out <= 32'h9d000000;
  11'h237: out <= 32'h00000008;
  11'h238: out <= 32'h00400000;
  11'h239: out <= 32'h03000000;
  11'h23a: out <= 32'h04000000;
  11'h23b: out <= 32'h2e010000;
  11'h23c: out <= 32'h006d656d;
  11'h23d: out <= 32'h03000000;
  11'h23e: out <= 32'h04000000;
  11'h23f: out <= 32'h03010000;
  11'h240: out <= 32'h02000000;
  11'h241: out <= 32'h02000000;
  11'h242: out <= 32'h01000000;
  11'h243: out <= 32'h406d6f72;
  11'h244: out <= 32'h30303031;
  11'h245: out <= 32'h00000030;
  11'h246: out <= 32'h03000000;
  11'h247: out <= 32'h10000000;
  11'h248: out <= 32'h1b000000;
  11'h249: out <= 32'h69666973;
  11'h24a: out <= 32'h6d2c6576;
  11'h24b: out <= 32'h726b7361;
  11'h24c: out <= 32'h00306d6f;
  11'h24d: out <= 32'h03000000;
  11'h24e: out <= 32'h08000000;
  11'h24f: out <= 32'h9d000000;
  11'h250: out <= 32'h00000100;
  11'h251: out <= 32'h00200000;
  11'h252: out <= 32'h03000000;
  11'h253: out <= 32'h04000000;
  11'h254: out <= 32'h2e010000;
  11'h255: out <= 32'h006d656d;
  11'h256: out <= 32'h02000000;
  11'h257: out <= 32'h01000000;
  11'h258: out <= 32'h69726573;
  11'h259: out <= 32'h31406c61;
  11'h25a: out <= 32'h33313030;
  11'h25b: out <= 32'h00303030;
  11'h25c: out <= 32'h03000000;
  11'h25d: out <= 32'h0d000000;
  11'h25e: out <= 32'h1b000000;
  11'h25f: out <= 32'h69666973;
  11'h260: out <= 32'h752c6576;
  11'h261: out <= 32'h30747261;
  11'h262: out <= 32'h00000000;
  11'h263: out <= 32'h03000000;
  11'h264: out <= 32'h04000000;
  11'h265: out <= 32'h12010000;
  11'h266: out <= 32'h03000000;
  11'h267: out <= 32'h03000000;
  11'h268: out <= 32'h04000000;
  11'h269: out <= 32'h23010000;
  11'h26a: out <= 32'h03000000;
  11'h26b: out <= 32'h03000000;
  11'h26c: out <= 32'h08000000;
  11'h26d: out <= 32'h9d000000;
  11'h26e: out <= 32'h00300110;
  11'h26f: out <= 32'h00100000;
  11'h270: out <= 32'h03000000;
  11'h271: out <= 32'h08000000;
  11'h272: out <= 32'h2e010000;
  11'h273: out <= 32'h746e6f63;
  11'h274: out <= 32'h006c6f72;
  11'h275: out <= 32'h02000000;
  11'h276: out <= 32'h01000000;
  11'h277: out <= 32'h69726573;
  11'h278: out <= 32'h31406c61;
  11'h279: out <= 32'h33323030;
  11'h27a: out <= 32'h00303030;
  11'h27b: out <= 32'h03000000;
  11'h27c: out <= 32'h0d000000;
  11'h27d: out <= 32'h1b000000;
  11'h27e: out <= 32'h69666973;
  11'h27f: out <= 32'h752c6576;
  11'h280: out <= 32'h30747261;
  11'h281: out <= 32'h00000000;
  11'h282: out <= 32'h03000000;
  11'h283: out <= 32'h04000000;
  11'h284: out <= 32'h12010000;
  11'h285: out <= 32'h03000000;
  11'h286: out <= 32'h03000000;
  11'h287: out <= 32'h04000000;
  11'h288: out <= 32'h23010000;
  11'h289: out <= 32'h04000000;
  11'h28a: out <= 32'h03000000;
  11'h28b: out <= 32'h08000000;
  11'h28c: out <= 32'h9d000000;
  11'h28d: out <= 32'h00300210;
  11'h28e: out <= 32'h00100000;
  11'h28f: out <= 32'h03000000;
  11'h290: out <= 32'h08000000;
  11'h291: out <= 32'h2e010000;
  11'h292: out <= 32'h746e6f63;
  11'h293: out <= 32'h006c6f72;
  11'h294: out <= 32'h02000000;
  11'h295: out <= 32'h01000000;
  11'h296: out <= 32'h69726573;
  11'h297: out <= 32'h31406c61;
  11'h298: out <= 32'h33333030;
  11'h299: out <= 32'h00303030;
  11'h29a: out <= 32'h03000000;
  11'h29b: out <= 32'h0d000000;
  11'h29c: out <= 32'h1b000000;
  11'h29d: out <= 32'h69666973;
  11'h29e: out <= 32'h752c6576;
  11'h29f: out <= 32'h30747261;
  11'h2a0: out <= 32'h00000000;
  11'h2a1: out <= 32'h03000000;
  11'h2a2: out <= 32'h04000000;
  11'h2a3: out <= 32'h12010000;
  11'h2a4: out <= 32'h03000000;
  11'h2a5: out <= 32'h03000000;
  11'h2a6: out <= 32'h04000000;
  11'h2a7: out <= 32'h23010000;
  11'h2a8: out <= 32'h05000000;
  11'h2a9: out <= 32'h03000000;
  11'h2aa: out <= 32'h08000000;
  11'h2ab: out <= 32'h9d000000;
  11'h2ac: out <= 32'h00300310;
  11'h2ad: out <= 32'h00100000;
  11'h2ae: out <= 32'h03000000;
  11'h2af: out <= 32'h08000000;
  11'h2b0: out <= 32'h2e010000;
  11'h2b1: out <= 32'h746e6f63;
  11'h2b2: out <= 32'h006c6f72;
  11'h2b3: out <= 32'h02000000;
  11'h2b4: out <= 32'h01000000;
  11'h2b5: out <= 32'h69726573;
  11'h2b6: out <= 32'h31406c61;
  11'h2b7: out <= 32'h33343030;
  11'h2b8: out <= 32'h00303030;
  11'h2b9: out <= 32'h03000000;
  11'h2ba: out <= 32'h0d000000;
  11'h2bb: out <= 32'h1b000000;
  11'h2bc: out <= 32'h69666973;
  11'h2bd: out <= 32'h752c6576;
  11'h2be: out <= 32'h30747261;
  11'h2bf: out <= 32'h00000000;
  11'h2c0: out <= 32'h03000000;
  11'h2c1: out <= 32'h04000000;
  11'h2c2: out <= 32'h12010000;
  11'h2c3: out <= 32'h03000000;
  11'h2c4: out <= 32'h03000000;
  11'h2c5: out <= 32'h04000000;
  11'h2c6: out <= 32'h23010000;
  11'h2c7: out <= 32'h06000000;
  11'h2c8: out <= 32'h03000000;
  11'h2c9: out <= 32'h08000000;
  11'h2ca: out <= 32'h9d000000;
  11'h2cb: out <= 32'h00300410;
  11'h2cc: out <= 32'h00100000;
  11'h2cd: out <= 32'h03000000;
  11'h2ce: out <= 32'h08000000;
  11'h2cf: out <= 32'h2e010000;
  11'h2d0: out <= 32'h746e6f63;
  11'h2d1: out <= 32'h006c6f72;
  11'h2d2: out <= 32'h02000000;
  11'h2d3: out <= 32'h01000000;
  11'h2d4: out <= 32'h69726573;
  11'h2d5: out <= 32'h31406c61;
  11'h2d6: out <= 32'h33353030;
  11'h2d7: out <= 32'h00303030;
  11'h2d8: out <= 32'h03000000;
  11'h2d9: out <= 32'h0d000000;
  11'h2da: out <= 32'h1b000000;
  11'h2db: out <= 32'h69666973;
  11'h2dc: out <= 32'h752c6576;
  11'h2dd: out <= 32'h30747261;
  11'h2de: out <= 32'h00000000;
  11'h2df: out <= 32'h03000000;
  11'h2e0: out <= 32'h04000000;
  11'h2e1: out <= 32'h12010000;
  11'h2e2: out <= 32'h03000000;
  11'h2e3: out <= 32'h03000000;
  11'h2e4: out <= 32'h04000000;
  11'h2e5: out <= 32'h23010000;
  11'h2e6: out <= 32'h07000000;
  11'h2e7: out <= 32'h03000000;
  11'h2e8: out <= 32'h08000000;
  11'h2e9: out <= 32'h9d000000;
  11'h2ea: out <= 32'h00300510;
  11'h2eb: out <= 32'h00100000;
  11'h2ec: out <= 32'h03000000;
  11'h2ed: out <= 32'h08000000;
  11'h2ee: out <= 32'h2e010000;
  11'h2ef: out <= 32'h746e6f63;
  11'h2f0: out <= 32'h006c6f72;
  11'h2f1: out <= 32'h02000000;
  11'h2f2: out <= 32'h01000000;
  11'h2f3: out <= 32'h40697073;
  11'h2f4: out <= 32'h31303031;
  11'h2f5: out <= 32'h30303034;
  11'h2f6: out <= 32'h00000000;
  11'h2f7: out <= 32'h03000000;
  11'h2f8: out <= 32'h04000000;
  11'h2f9: out <= 32'h00000000;
  11'h2fa: out <= 32'h01000000;
  11'h2fb: out <= 32'h03000000;
  11'h2fc: out <= 32'h04000000;
  11'h2fd: out <= 32'h0f000000;
  11'h2fe: out <= 32'h00000000;
  11'h2ff: out <= 32'h03000000;
  11'h300: out <= 32'h0c000000;
  11'h301: out <= 32'h1b000000;
  11'h302: out <= 32'h69666973;
  11'h303: out <= 32'h732c6576;
  11'h304: out <= 32'h00306970;
  11'h305: out <= 32'h03000000;
  11'h306: out <= 32'h04000000;
  11'h307: out <= 32'h12010000;
  11'h308: out <= 32'h03000000;
  11'h309: out <= 32'h03000000;
  11'h30a: out <= 32'h04000000;
  11'h30b: out <= 32'h23010000;
  11'h30c: out <= 32'h08000000;
  11'h30d: out <= 32'h03000000;
  11'h30e: out <= 32'h10000000;
  11'h30f: out <= 32'h9d000000;
  11'h310: out <= 32'h00400110;
  11'h311: out <= 32'h00100000;
  11'h312: out <= 32'h00000020;
  11'h313: out <= 32'h00000020;
  11'h314: out <= 32'h03000000;
  11'h315: out <= 32'h0c000000;
  11'h316: out <= 32'h2e010000;
  11'h317: out <= 32'h746e6f63;
  11'h318: out <= 32'h006c6f72;
  11'h319: out <= 32'h006d656d;
  11'h31a: out <= 32'h02000000;
  11'h31b: out <= 32'h01000000;
  11'h31c: out <= 32'h40697073;
  11'h31d: out <= 32'h32303031;
  11'h31e: out <= 32'h30303034;
  11'h31f: out <= 32'h00000000;
  11'h320: out <= 32'h03000000;
  11'h321: out <= 32'h04000000;
  11'h322: out <= 32'h00000000;
  11'h323: out <= 32'h01000000;
  11'h324: out <= 32'h03000000;
  11'h325: out <= 32'h04000000;
  11'h326: out <= 32'h0f000000;
  11'h327: out <= 32'h00000000;
  11'h328: out <= 32'h03000000;
  11'h329: out <= 32'h0c000000;
  11'h32a: out <= 32'h1b000000;
  11'h32b: out <= 32'h69666973;
  11'h32c: out <= 32'h732c6576;
  11'h32d: out <= 32'h00306970;
  11'h32e: out <= 32'h03000000;
  11'h32f: out <= 32'h04000000;
  11'h330: out <= 32'h12010000;
  11'h331: out <= 32'h03000000;
  11'h332: out <= 32'h03000000;
  11'h333: out <= 32'h04000000;
  11'h334: out <= 32'h23010000;
  11'h335: out <= 32'h09000000;
  11'h336: out <= 32'h03000000;
  11'h337: out <= 32'h08000000;
  11'h338: out <= 32'h9d000000;
  11'h339: out <= 32'h00400210;
  11'h33a: out <= 32'h00100000;
  11'h33b: out <= 32'h03000000;
  11'h33c: out <= 32'h08000000;
  11'h33d: out <= 32'h2e010000;
  11'h33e: out <= 32'h746e6f63;
  11'h33f: out <= 32'h006c6f72;
  11'h340: out <= 32'h02000000;
  11'h341: out <= 32'h01000000;
  11'h342: out <= 32'h40697073;
  11'h343: out <= 32'h33303031;
  11'h344: out <= 32'h30303034;
  11'h345: out <= 32'h00000000;
  11'h346: out <= 32'h03000000;
  11'h347: out <= 32'h04000000;
  11'h348: out <= 32'h00000000;
  11'h349: out <= 32'h01000000;
  11'h34a: out <= 32'h03000000;
  11'h34b: out <= 32'h04000000;
  11'h34c: out <= 32'h0f000000;
  11'h34d: out <= 32'h00000000;
  11'h34e: out <= 32'h03000000;
  11'h34f: out <= 32'h0c000000;
  11'h350: out <= 32'h1b000000;
  11'h351: out <= 32'h69666973;
  11'h352: out <= 32'h732c6576;
  11'h353: out <= 32'h00306970;
  11'h354: out <= 32'h03000000;
  11'h355: out <= 32'h04000000;
  11'h356: out <= 32'h12010000;
  11'h357: out <= 32'h03000000;
  11'h358: out <= 32'h03000000;
  11'h359: out <= 32'h04000000;
  11'h35a: out <= 32'h23010000;
  11'h35b: out <= 32'h0a000000;
  11'h35c: out <= 32'h03000000;
  11'h35d: out <= 32'h08000000;
  11'h35e: out <= 32'h9d000000;
  11'h35f: out <= 32'h00400310;
  11'h360: out <= 32'h00100000;
  11'h361: out <= 32'h03000000;
  11'h362: out <= 32'h08000000;
  11'h363: out <= 32'h2e010000;
  11'h364: out <= 32'h746e6f63;
  11'h365: out <= 32'h006c6f72;
  11'h366: out <= 32'h02000000;
  11'h367: out <= 32'h02000000;
  11'h368: out <= 32'h02000000;
  11'h369: out <= 32'h09000000;
  11'h36a: out <= 32'h64646123;
  11'h36b: out <= 32'h73736572;
  11'h36c: out <= 32'h6c65632d;
  11'h36d: out <= 32'h2300736c;
  11'h36e: out <= 32'h657a6973;
  11'h36f: out <= 32'h6c65632d;
  11'h370: out <= 32'h6300736c;
  11'h371: out <= 32'h61706d6f;
  11'h372: out <= 32'h6c626974;
  11'h373: out <= 32'h6f6d0065;
  11'h374: out <= 32'h006c6564;
  11'h375: out <= 32'h69726573;
  11'h376: out <= 32'h00306c61;
  11'h377: out <= 32'h69726573;
  11'h378: out <= 32'h00316c61;
  11'h379: out <= 32'h69726573;
  11'h37a: out <= 32'h00326c61;
  11'h37b: out <= 32'h69726573;
  11'h37c: out <= 32'h00336c61;
  11'h37d: out <= 32'h69726573;
  11'h37e: out <= 32'h00346c61;
  11'h37f: out <= 32'h636f6c63;
  11'h380: out <= 32'h72662d6b;
  11'h381: out <= 32'h65757165;
  11'h382: out <= 32'h0079636e;
  11'h383: out <= 32'h69766564;
  11'h384: out <= 32'h745f6563;
  11'h385: out <= 32'h00657079;
  11'h386: out <= 32'h61632d69;
  11'h387: out <= 32'h2d656863;
  11'h388: out <= 32'h636f6c62;
  11'h389: out <= 32'h69732d6b;
  11'h38a: out <= 32'h6900657a;
  11'h38b: out <= 32'h6361632d;
  11'h38c: out <= 32'h732d6568;
  11'h38d: out <= 32'h00737465;
  11'h38e: out <= 32'h61632d69;
  11'h38f: out <= 32'h2d656863;
  11'h390: out <= 32'h657a6973;
  11'h391: out <= 32'h67657200;
  11'h392: out <= 32'h73697200;
  11'h393: out <= 32'h692c7663;
  11'h394: out <= 32'h73006173;
  11'h395: out <= 32'h76696669;
  11'h396: out <= 32'h74642c65;
  11'h397: out <= 32'h73006d69;
  11'h398: out <= 32'h76696669;
  11'h399: out <= 32'h74692c65;
  11'h39a: out <= 32'h73006d69;
  11'h39b: out <= 32'h75746174;
  11'h39c: out <= 32'h69740073;
  11'h39d: out <= 32'h6162656d;
  11'h39e: out <= 32'h662d6573;
  11'h39f: out <= 32'h75716572;
  11'h3a0: out <= 32'h79636e65;
  11'h3a1: out <= 32'h6e692300;
  11'h3a2: out <= 32'h72726574;
  11'h3a3: out <= 32'h2d747075;
  11'h3a4: out <= 32'h6c6c6563;
  11'h3a5: out <= 32'h6e690073;
  11'h3a6: out <= 32'h72726574;
  11'h3a7: out <= 32'h2d747075;
  11'h3a8: out <= 32'h746e6f63;
  11'h3a9: out <= 32'h6c6c6f72;
  11'h3aa: out <= 32'h70007265;
  11'h3ab: out <= 32'h646e6168;
  11'h3ac: out <= 32'h7200656c;
  11'h3ad: out <= 32'h65676e61;
  11'h3ae: out <= 32'h6e690073;
  11'h3af: out <= 32'h72726574;
  11'h3b0: out <= 32'h2d747075;
  11'h3b1: out <= 32'h65726170;
  11'h3b2: out <= 32'h6900746e;
  11'h3b3: out <= 32'h7265746e;
  11'h3b4: out <= 32'h74707572;
  11'h3b5: out <= 32'h65720073;
  11'h3b6: out <= 32'h616e2d67;
  11'h3b7: out <= 32'h0073656d;
  11'h3b8: out <= 32'h65746e69;
  11'h3b9: out <= 32'h70757272;
  11'h3ba: out <= 32'h652d7374;
  11'h3bb: out <= 32'h6e657478;
  11'h3bc: out <= 32'h00646564;
  11'h3bd: out <= 32'h69706723;
  11'h3be: out <= 32'h65632d6f;
  11'h3bf: out <= 32'h00736c6c;
  11'h3c0: out <= 32'h6f697067;
  11'h3c1: out <= 32'h6e6f632d;
  11'h3c2: out <= 32'h6c6f7274;
  11'h3c3: out <= 32'h0072656c;
  11'h3c4: out <= 32'h63736972;
  11'h3c5: out <= 32'h616d2c76;
  11'h3c6: out <= 32'h72702d78;
  11'h3c7: out <= 32'h69726f69;
  11'h3c8: out <= 32'h72007974;
  11'h3c9: out <= 32'h76637369;
  11'h3ca: out <= 32'h65646e2c;
  11'h3cb: out <= 32'h00000076;
  default: out <= 32'hdeadbeef;
endcase
