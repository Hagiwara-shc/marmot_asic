magic
tech sky130A
magscale 1 2
timestamp 1653216700
<< obsli1 >>
rect 201104 62159 555856 416881
<< obsm1 >>
rect 566 960 582438 700732
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 583432 703610
rect 572 536 583432 703464
rect 710 326 1590 536
rect 1814 326 2786 536
rect 3010 326 3982 536
rect 4206 326 5178 536
rect 5402 326 6374 536
rect 6598 326 7570 536
rect 7794 326 8674 536
rect 8898 326 9870 536
rect 10094 326 11066 536
rect 11290 326 12262 536
rect 12486 326 13458 536
rect 13682 326 14654 536
rect 14878 326 15850 536
rect 16074 326 16954 536
rect 17178 326 18150 536
rect 18374 326 19346 536
rect 19570 326 20542 536
rect 20766 326 21738 536
rect 21962 326 22934 536
rect 23158 326 24130 536
rect 24354 326 25234 536
rect 25458 326 26430 536
rect 26654 326 27626 536
rect 27850 326 28822 536
rect 29046 326 30018 536
rect 30242 326 31214 536
rect 31438 326 32318 536
rect 32542 326 33514 536
rect 33738 326 34710 536
rect 34934 326 35906 536
rect 36130 326 37102 536
rect 37326 326 38298 536
rect 38522 326 39494 536
rect 39718 326 40598 536
rect 40822 326 41794 536
rect 42018 326 42990 536
rect 43214 326 44186 536
rect 44410 326 45382 536
rect 45606 326 46578 536
rect 46802 326 47774 536
rect 47998 326 48878 536
rect 49102 326 50074 536
rect 50298 326 51270 536
rect 51494 326 52466 536
rect 52690 326 53662 536
rect 53886 326 54858 536
rect 55082 326 55962 536
rect 56186 326 57158 536
rect 57382 326 58354 536
rect 58578 326 59550 536
rect 59774 326 60746 536
rect 60970 326 61942 536
rect 62166 326 63138 536
rect 63362 326 64242 536
rect 64466 326 65438 536
rect 65662 326 66634 536
rect 66858 326 67830 536
rect 68054 326 69026 536
rect 69250 326 70222 536
rect 70446 326 71418 536
rect 71642 326 72522 536
rect 72746 326 73718 536
rect 73942 326 74914 536
rect 75138 326 76110 536
rect 76334 326 77306 536
rect 77530 326 78502 536
rect 78726 326 79606 536
rect 79830 326 80802 536
rect 81026 326 81998 536
rect 82222 326 83194 536
rect 83418 326 84390 536
rect 84614 326 85586 536
rect 85810 326 86782 536
rect 87006 326 87886 536
rect 88110 326 89082 536
rect 89306 326 90278 536
rect 90502 326 91474 536
rect 91698 326 92670 536
rect 92894 326 93866 536
rect 94090 326 95062 536
rect 95286 326 96166 536
rect 96390 326 97362 536
rect 97586 326 98558 536
rect 98782 326 99754 536
rect 99978 326 100950 536
rect 101174 326 102146 536
rect 102370 326 103250 536
rect 103474 326 104446 536
rect 104670 326 105642 536
rect 105866 326 106838 536
rect 107062 326 108034 536
rect 108258 326 109230 536
rect 109454 326 110426 536
rect 110650 326 111530 536
rect 111754 326 112726 536
rect 112950 326 113922 536
rect 114146 326 115118 536
rect 115342 326 116314 536
rect 116538 326 117510 536
rect 117734 326 118706 536
rect 118930 326 119810 536
rect 120034 326 121006 536
rect 121230 326 122202 536
rect 122426 326 123398 536
rect 123622 326 124594 536
rect 124818 326 125790 536
rect 126014 326 126894 536
rect 127118 326 128090 536
rect 128314 326 129286 536
rect 129510 326 130482 536
rect 130706 326 131678 536
rect 131902 326 132874 536
rect 133098 326 134070 536
rect 134294 326 135174 536
rect 135398 326 136370 536
rect 136594 326 137566 536
rect 137790 326 138762 536
rect 138986 326 139958 536
rect 140182 326 141154 536
rect 141378 326 142350 536
rect 142574 326 143454 536
rect 143678 326 144650 536
rect 144874 326 145846 536
rect 146070 326 147042 536
rect 147266 326 148238 536
rect 148462 326 149434 536
rect 149658 326 150538 536
rect 150762 326 151734 536
rect 151958 326 152930 536
rect 153154 326 154126 536
rect 154350 326 155322 536
rect 155546 326 156518 536
rect 156742 326 157714 536
rect 157938 326 158818 536
rect 159042 326 160014 536
rect 160238 326 161210 536
rect 161434 326 162406 536
rect 162630 326 163602 536
rect 163826 326 164798 536
rect 165022 326 165994 536
rect 166218 326 167098 536
rect 167322 326 168294 536
rect 168518 326 169490 536
rect 169714 326 170686 536
rect 170910 326 171882 536
rect 172106 326 173078 536
rect 173302 326 174182 536
rect 174406 326 175378 536
rect 175602 326 176574 536
rect 176798 326 177770 536
rect 177994 326 178966 536
rect 179190 326 180162 536
rect 180386 326 181358 536
rect 181582 326 182462 536
rect 182686 326 183658 536
rect 183882 326 184854 536
rect 185078 326 186050 536
rect 186274 326 187246 536
rect 187470 326 188442 536
rect 188666 326 189638 536
rect 189862 326 190742 536
rect 190966 326 191938 536
rect 192162 326 193134 536
rect 193358 326 194330 536
rect 194554 326 195526 536
rect 195750 326 196722 536
rect 196946 326 197826 536
rect 198050 326 199022 536
rect 199246 326 200218 536
rect 200442 326 201414 536
rect 201638 326 202610 536
rect 202834 326 203806 536
rect 204030 326 205002 536
rect 205226 326 206106 536
rect 206330 326 207302 536
rect 207526 326 208498 536
rect 208722 326 209694 536
rect 209918 326 210890 536
rect 211114 326 212086 536
rect 212310 326 213282 536
rect 213506 326 214386 536
rect 214610 326 215582 536
rect 215806 326 216778 536
rect 217002 326 217974 536
rect 218198 326 219170 536
rect 219394 326 220366 536
rect 220590 326 221470 536
rect 221694 326 222666 536
rect 222890 326 223862 536
rect 224086 326 225058 536
rect 225282 326 226254 536
rect 226478 326 227450 536
rect 227674 326 228646 536
rect 228870 326 229750 536
rect 229974 326 230946 536
rect 231170 326 232142 536
rect 232366 326 233338 536
rect 233562 326 234534 536
rect 234758 326 235730 536
rect 235954 326 236926 536
rect 237150 326 238030 536
rect 238254 326 239226 536
rect 239450 326 240422 536
rect 240646 326 241618 536
rect 241842 326 242814 536
rect 243038 326 244010 536
rect 244234 326 245114 536
rect 245338 326 246310 536
rect 246534 326 247506 536
rect 247730 326 248702 536
rect 248926 326 249898 536
rect 250122 326 251094 536
rect 251318 326 252290 536
rect 252514 326 253394 536
rect 253618 326 254590 536
rect 254814 326 255786 536
rect 256010 326 256982 536
rect 257206 326 258178 536
rect 258402 326 259374 536
rect 259598 326 260570 536
rect 260794 326 261674 536
rect 261898 326 262870 536
rect 263094 326 264066 536
rect 264290 326 265262 536
rect 265486 326 266458 536
rect 266682 326 267654 536
rect 267878 326 268758 536
rect 268982 326 269954 536
rect 270178 326 271150 536
rect 271374 326 272346 536
rect 272570 326 273542 536
rect 273766 326 274738 536
rect 274962 326 275934 536
rect 276158 326 277038 536
rect 277262 326 278234 536
rect 278458 326 279430 536
rect 279654 326 280626 536
rect 280850 326 281822 536
rect 282046 326 283018 536
rect 283242 326 284214 536
rect 284438 326 285318 536
rect 285542 326 286514 536
rect 286738 326 287710 536
rect 287934 326 288906 536
rect 289130 326 290102 536
rect 290326 326 291298 536
rect 291522 326 292494 536
rect 292718 326 293598 536
rect 293822 326 294794 536
rect 295018 326 295990 536
rect 296214 326 297186 536
rect 297410 326 298382 536
rect 298606 326 299578 536
rect 299802 326 300682 536
rect 300906 326 301878 536
rect 302102 326 303074 536
rect 303298 326 304270 536
rect 304494 326 305466 536
rect 305690 326 306662 536
rect 306886 326 307858 536
rect 308082 326 308962 536
rect 309186 326 310158 536
rect 310382 326 311354 536
rect 311578 326 312550 536
rect 312774 326 313746 536
rect 313970 326 314942 536
rect 315166 326 316138 536
rect 316362 326 317242 536
rect 317466 326 318438 536
rect 318662 326 319634 536
rect 319858 326 320830 536
rect 321054 326 322026 536
rect 322250 326 323222 536
rect 323446 326 324326 536
rect 324550 326 325522 536
rect 325746 326 326718 536
rect 326942 326 327914 536
rect 328138 326 329110 536
rect 329334 326 330306 536
rect 330530 326 331502 536
rect 331726 326 332606 536
rect 332830 326 333802 536
rect 334026 326 334998 536
rect 335222 326 336194 536
rect 336418 326 337390 536
rect 337614 326 338586 536
rect 338810 326 339782 536
rect 340006 326 340886 536
rect 341110 326 342082 536
rect 342306 326 343278 536
rect 343502 326 344474 536
rect 344698 326 345670 536
rect 345894 326 346866 536
rect 347090 326 347970 536
rect 348194 326 349166 536
rect 349390 326 350362 536
rect 350586 326 351558 536
rect 351782 326 352754 536
rect 352978 326 353950 536
rect 354174 326 355146 536
rect 355370 326 356250 536
rect 356474 326 357446 536
rect 357670 326 358642 536
rect 358866 326 359838 536
rect 360062 326 361034 536
rect 361258 326 362230 536
rect 362454 326 363426 536
rect 363650 326 364530 536
rect 364754 326 365726 536
rect 365950 326 366922 536
rect 367146 326 368118 536
rect 368342 326 369314 536
rect 369538 326 370510 536
rect 370734 326 371614 536
rect 371838 326 372810 536
rect 373034 326 374006 536
rect 374230 326 375202 536
rect 375426 326 376398 536
rect 376622 326 377594 536
rect 377818 326 378790 536
rect 379014 326 379894 536
rect 380118 326 381090 536
rect 381314 326 382286 536
rect 382510 326 383482 536
rect 383706 326 384678 536
rect 384902 326 385874 536
rect 386098 326 387070 536
rect 387294 326 388174 536
rect 388398 326 389370 536
rect 389594 326 390566 536
rect 390790 326 391762 536
rect 391986 326 392958 536
rect 393182 326 394154 536
rect 394378 326 395258 536
rect 395482 326 396454 536
rect 396678 326 397650 536
rect 397874 326 398846 536
rect 399070 326 400042 536
rect 400266 326 401238 536
rect 401462 326 402434 536
rect 402658 326 403538 536
rect 403762 326 404734 536
rect 404958 326 405930 536
rect 406154 326 407126 536
rect 407350 326 408322 536
rect 408546 326 409518 536
rect 409742 326 410714 536
rect 410938 326 411818 536
rect 412042 326 413014 536
rect 413238 326 414210 536
rect 414434 326 415406 536
rect 415630 326 416602 536
rect 416826 326 417798 536
rect 418022 326 418902 536
rect 419126 326 420098 536
rect 420322 326 421294 536
rect 421518 326 422490 536
rect 422714 326 423686 536
rect 423910 326 424882 536
rect 425106 326 426078 536
rect 426302 326 427182 536
rect 427406 326 428378 536
rect 428602 326 429574 536
rect 429798 326 430770 536
rect 430994 326 431966 536
rect 432190 326 433162 536
rect 433386 326 434358 536
rect 434582 326 435462 536
rect 435686 326 436658 536
rect 436882 326 437854 536
rect 438078 326 439050 536
rect 439274 326 440246 536
rect 440470 326 441442 536
rect 441666 326 442546 536
rect 442770 326 443742 536
rect 443966 326 444938 536
rect 445162 326 446134 536
rect 446358 326 447330 536
rect 447554 326 448526 536
rect 448750 326 449722 536
rect 449946 326 450826 536
rect 451050 326 452022 536
rect 452246 326 453218 536
rect 453442 326 454414 536
rect 454638 326 455610 536
rect 455834 326 456806 536
rect 457030 326 458002 536
rect 458226 326 459106 536
rect 459330 326 460302 536
rect 460526 326 461498 536
rect 461722 326 462694 536
rect 462918 326 463890 536
rect 464114 326 465086 536
rect 465310 326 466190 536
rect 466414 326 467386 536
rect 467610 326 468582 536
rect 468806 326 469778 536
rect 470002 326 470974 536
rect 471198 326 472170 536
rect 472394 326 473366 536
rect 473590 326 474470 536
rect 474694 326 475666 536
rect 475890 326 476862 536
rect 477086 326 478058 536
rect 478282 326 479254 536
rect 479478 326 480450 536
rect 480674 326 481646 536
rect 481870 326 482750 536
rect 482974 326 483946 536
rect 484170 326 485142 536
rect 485366 326 486338 536
rect 486562 326 487534 536
rect 487758 326 488730 536
rect 488954 326 489834 536
rect 490058 326 491030 536
rect 491254 326 492226 536
rect 492450 326 493422 536
rect 493646 326 494618 536
rect 494842 326 495814 536
rect 496038 326 497010 536
rect 497234 326 498114 536
rect 498338 326 499310 536
rect 499534 326 500506 536
rect 500730 326 501702 536
rect 501926 326 502898 536
rect 503122 326 504094 536
rect 504318 326 505290 536
rect 505514 326 506394 536
rect 506618 326 507590 536
rect 507814 326 508786 536
rect 509010 326 509982 536
rect 510206 326 511178 536
rect 511402 326 512374 536
rect 512598 326 513478 536
rect 513702 326 514674 536
rect 514898 326 515870 536
rect 516094 326 517066 536
rect 517290 326 518262 536
rect 518486 326 519458 536
rect 519682 326 520654 536
rect 520878 326 521758 536
rect 521982 326 522954 536
rect 523178 326 524150 536
rect 524374 326 525346 536
rect 525570 326 526542 536
rect 526766 326 527738 536
rect 527962 326 528934 536
rect 529158 326 530038 536
rect 530262 326 531234 536
rect 531458 326 532430 536
rect 532654 326 533626 536
rect 533850 326 534822 536
rect 535046 326 536018 536
rect 536242 326 537122 536
rect 537346 326 538318 536
rect 538542 326 539514 536
rect 539738 326 540710 536
rect 540934 326 541906 536
rect 542130 326 543102 536
rect 543326 326 544298 536
rect 544522 326 545402 536
rect 545626 326 546598 536
rect 546822 326 547794 536
rect 548018 326 548990 536
rect 549214 326 550186 536
rect 550410 326 551382 536
rect 551606 326 552578 536
rect 552802 326 553682 536
rect 553906 326 554878 536
rect 555102 326 556074 536
rect 556298 326 557270 536
rect 557494 326 558466 536
rect 558690 326 559662 536
rect 559886 326 560766 536
rect 560990 326 561962 536
rect 562186 326 563158 536
rect 563382 326 564354 536
rect 564578 326 565550 536
rect 565774 326 566746 536
rect 566970 326 567942 536
rect 568166 326 569046 536
rect 569270 326 570242 536
rect 570466 326 571438 536
rect 571662 326 572634 536
rect 572858 326 573830 536
rect 574054 326 575026 536
rect 575250 326 576222 536
rect 576446 326 577326 536
rect 577550 326 578522 536
rect 578746 326 579718 536
rect 579942 326 580914 536
rect 581138 326 582110 536
rect 582334 326 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 246 697540 583520 700637
rect 560 697404 583520 697540
rect 560 697140 583440 697404
rect 246 697004 583440 697140
rect 246 684484 583520 697004
rect 560 684084 583520 684484
rect 246 684076 583520 684084
rect 246 683676 583440 684076
rect 246 671428 583520 683676
rect 560 671028 583520 671428
rect 246 670884 583520 671028
rect 246 670484 583440 670884
rect 246 658372 583520 670484
rect 560 657972 583520 658372
rect 246 657556 583520 657972
rect 246 657156 583440 657556
rect 246 645316 583520 657156
rect 560 644916 583520 645316
rect 246 644228 583520 644916
rect 246 643828 583440 644228
rect 246 632260 583520 643828
rect 560 631860 583520 632260
rect 246 631036 583520 631860
rect 246 630636 583440 631036
rect 246 619340 583520 630636
rect 560 618940 583520 619340
rect 246 617708 583520 618940
rect 246 617308 583440 617708
rect 246 606284 583520 617308
rect 560 605884 583520 606284
rect 246 604380 583520 605884
rect 246 603980 583440 604380
rect 246 593228 583520 603980
rect 560 592828 583520 593228
rect 246 591188 583520 592828
rect 246 590788 583440 591188
rect 246 580172 583520 590788
rect 560 579772 583520 580172
rect 246 577860 583520 579772
rect 246 577460 583440 577860
rect 246 567116 583520 577460
rect 560 566716 583520 567116
rect 246 564532 583520 566716
rect 246 564132 583440 564532
rect 246 554060 583520 564132
rect 560 553660 583520 554060
rect 246 551340 583520 553660
rect 246 550940 583440 551340
rect 246 541004 583520 550940
rect 560 540604 583520 541004
rect 246 538012 583520 540604
rect 246 537612 583440 538012
rect 246 528084 583520 537612
rect 560 527684 583520 528084
rect 246 524684 583520 527684
rect 246 524284 583440 524684
rect 246 515028 583520 524284
rect 560 514628 583520 515028
rect 246 511492 583520 514628
rect 246 511092 583440 511492
rect 246 501972 583520 511092
rect 560 501572 583520 501972
rect 246 498164 583520 501572
rect 246 497764 583440 498164
rect 246 488916 583520 497764
rect 560 488516 583520 488916
rect 246 484836 583520 488516
rect 246 484436 583440 484836
rect 246 475860 583520 484436
rect 560 475460 583520 475860
rect 246 471644 583520 475460
rect 246 471244 583440 471644
rect 246 462804 583520 471244
rect 560 462404 583520 462804
rect 246 458316 583520 462404
rect 246 457916 583440 458316
rect 246 449748 583520 457916
rect 560 449348 583520 449748
rect 246 444988 583520 449348
rect 246 444588 583440 444988
rect 246 436828 583520 444588
rect 560 436428 583520 436828
rect 246 431796 583520 436428
rect 246 431396 583440 431796
rect 246 423772 583520 431396
rect 560 423372 583520 423772
rect 246 418468 583520 423372
rect 246 418068 583440 418468
rect 246 410716 583520 418068
rect 560 410316 583520 410716
rect 246 405140 583520 410316
rect 246 404740 583440 405140
rect 246 397660 583520 404740
rect 560 397260 583520 397660
rect 246 391948 583520 397260
rect 246 391548 583440 391948
rect 246 384604 583520 391548
rect 560 384204 583520 384604
rect 246 378620 583520 384204
rect 246 378220 583440 378620
rect 246 371548 583520 378220
rect 560 371148 583520 371548
rect 246 365292 583520 371148
rect 246 364892 583440 365292
rect 246 358628 583520 364892
rect 560 358228 583520 358628
rect 246 352100 583520 358228
rect 246 351700 583440 352100
rect 246 345572 583520 351700
rect 560 345172 583520 345572
rect 246 338772 583520 345172
rect 246 338372 583440 338772
rect 246 332516 583520 338372
rect 560 332116 583520 332516
rect 246 325444 583520 332116
rect 246 325044 583440 325444
rect 246 319460 583520 325044
rect 560 319060 583520 319460
rect 246 312252 583520 319060
rect 246 311852 583440 312252
rect 246 306404 583520 311852
rect 560 306004 583520 306404
rect 246 298924 583520 306004
rect 246 298524 583440 298924
rect 246 293348 583520 298524
rect 560 292948 583520 293348
rect 246 285596 583520 292948
rect 246 285196 583440 285596
rect 246 280292 583520 285196
rect 560 279892 583520 280292
rect 246 272404 583520 279892
rect 246 272004 583440 272404
rect 246 267372 583520 272004
rect 560 266972 583520 267372
rect 246 259076 583520 266972
rect 246 258676 583440 259076
rect 246 254316 583520 258676
rect 560 253916 583520 254316
rect 246 245748 583520 253916
rect 246 245348 583440 245748
rect 246 241260 583520 245348
rect 560 240860 583520 241260
rect 246 232556 583520 240860
rect 246 232156 583440 232556
rect 246 228204 583520 232156
rect 560 227804 583520 228204
rect 246 219228 583520 227804
rect 246 218828 583440 219228
rect 246 215148 583520 218828
rect 560 214748 583520 215148
rect 246 205900 583520 214748
rect 246 205500 583440 205900
rect 246 202092 583520 205500
rect 560 201692 583520 202092
rect 246 192708 583520 201692
rect 246 192308 583440 192708
rect 246 189036 583520 192308
rect 560 188636 583520 189036
rect 246 179380 583520 188636
rect 246 178980 583440 179380
rect 246 176116 583520 178980
rect 560 175716 583520 176116
rect 246 166052 583520 175716
rect 246 165652 583440 166052
rect 246 163060 583520 165652
rect 560 162660 583520 163060
rect 246 152860 583520 162660
rect 246 152460 583440 152860
rect 246 150004 583520 152460
rect 560 149604 583520 150004
rect 246 139532 583520 149604
rect 246 139132 583440 139532
rect 246 136948 583520 139132
rect 560 136548 583520 136948
rect 246 126204 583520 136548
rect 246 125804 583440 126204
rect 246 123892 583520 125804
rect 560 123492 583520 123892
rect 246 113012 583520 123492
rect 246 112612 583440 113012
rect 246 110836 583520 112612
rect 560 110436 583520 110836
rect 246 99684 583520 110436
rect 246 99284 583440 99684
rect 246 97780 583520 99284
rect 560 97380 583520 97780
rect 246 86356 583520 97380
rect 246 85956 583440 86356
rect 246 84860 583520 85956
rect 560 84460 583520 84860
rect 246 73164 583520 84460
rect 246 72764 583440 73164
rect 246 71804 583520 72764
rect 560 71404 583520 71804
rect 246 59836 583520 71404
rect 246 59436 583440 59836
rect 246 58748 583520 59436
rect 560 58348 583520 58748
rect 246 46508 583520 58348
rect 246 46108 583440 46508
rect 246 45692 583520 46108
rect 560 45292 583520 45692
rect 246 33316 583520 45292
rect 246 32916 583440 33316
rect 246 32636 583520 32916
rect 560 32236 583520 32636
rect 246 19988 583520 32236
rect 246 19588 583440 19988
rect 246 19580 583520 19588
rect 560 19180 583520 19580
rect 246 6796 583520 19180
rect 246 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 246 5612 583520 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 9234 -5734 9854 709670
rect 11794 -1894 12414 705830
rect 12954 -7654 13574 711590
rect 15514 -3814 16134 707750
rect 19234 -5734 19854 709670
rect 21794 -1894 22414 705830
rect 22954 -7654 23574 711590
rect 25514 -3814 26134 707750
rect 29234 675308 29854 709670
rect 31794 675308 32414 705830
rect 32954 675308 33574 711590
rect 35514 675308 36134 707750
rect 39234 675308 39854 709670
rect 41794 675308 42414 705830
rect 42954 675308 43574 711590
rect 45514 675308 46134 707750
rect 49234 675308 49854 709670
rect 51794 675308 52414 705830
rect 52954 675308 53574 711590
rect 55514 675308 56134 707750
rect 59234 675308 59854 709670
rect 61794 675308 62414 705830
rect 62954 675308 63574 711590
rect 65514 675308 66134 707750
rect 69234 675308 69854 709670
rect 71794 675308 72414 705830
rect 72954 675308 73574 711590
rect 75514 675308 76134 707750
rect 79234 675308 79854 709670
rect 81794 675308 82414 705830
rect 82954 675308 83574 711590
rect 85514 675308 86134 707750
rect 89234 675308 89854 709670
rect 91794 675308 92414 705830
rect 92954 675308 93574 711590
rect 95514 675308 96134 707750
rect 99234 675308 99854 709670
rect 101794 675308 102414 705830
rect 102954 675308 103574 711590
rect 105514 675308 106134 707750
rect 109234 675308 109854 709670
rect 111794 675308 112414 705830
rect 112954 675308 113574 711590
rect 115514 675308 116134 707750
rect 119234 675308 119854 709670
rect 121794 675308 122414 705830
rect 122954 675308 123574 711590
rect 125514 675308 126134 707750
rect 129234 675308 129854 709670
rect 131794 675308 132414 705830
rect 132954 675308 133574 711590
rect 135514 675308 136134 707750
rect 139234 675308 139854 709670
rect 141794 675308 142414 705830
rect 142954 675308 143574 711590
rect 145514 675308 146134 707750
rect 149234 675308 149854 709670
rect 151794 675308 152414 705830
rect 152954 675308 153574 711590
rect 155514 675308 156134 707750
rect 159234 675308 159854 709670
rect 161794 675308 162414 705830
rect 162954 675308 163574 711590
rect 165514 675308 166134 707750
rect 29234 563308 29854 588000
rect 31794 563308 32414 588000
rect 32954 563308 33574 588000
rect 35514 563308 36134 588000
rect 39234 563308 39854 588000
rect 41794 563308 42414 588000
rect 42954 563308 43574 588000
rect 45514 563308 46134 588000
rect 49234 563308 49854 588000
rect 51794 563308 52414 588000
rect 52954 563308 53574 588000
rect 55514 563308 56134 588000
rect 59234 563308 59854 588000
rect 61794 563308 62414 588000
rect 62954 563308 63574 588000
rect 65514 563308 66134 588000
rect 69234 563308 69854 588000
rect 71794 563308 72414 588000
rect 72954 563308 73574 588000
rect 75514 563308 76134 588000
rect 79234 563308 79854 588000
rect 81794 563308 82414 588000
rect 82954 563308 83574 588000
rect 85514 563308 86134 588000
rect 89234 563308 89854 588000
rect 91794 563308 92414 588000
rect 92954 563308 93574 588000
rect 95514 563308 96134 588000
rect 99234 563308 99854 588000
rect 101794 563308 102414 588000
rect 102954 563308 103574 588000
rect 105514 563308 106134 588000
rect 109234 563308 109854 588000
rect 111794 563308 112414 588000
rect 112954 563308 113574 588000
rect 115514 563308 116134 588000
rect 119234 563308 119854 588000
rect 121794 563308 122414 588000
rect 122954 563308 123574 588000
rect 125514 563308 126134 588000
rect 129234 563308 129854 588000
rect 131794 563308 132414 588000
rect 132954 563308 133574 588000
rect 135514 563308 136134 588000
rect 139234 563308 139854 588000
rect 141794 563308 142414 588000
rect 142954 563308 143574 588000
rect 145514 563308 146134 588000
rect 149234 563308 149854 588000
rect 151794 563308 152414 588000
rect 152954 563308 153574 588000
rect 155514 563308 156134 588000
rect 159234 563308 159854 588000
rect 161794 563308 162414 588000
rect 162954 563308 163574 588000
rect 165514 563308 166134 588000
rect 29234 451308 29854 476000
rect 31794 451308 32414 476000
rect 32954 451308 33574 476000
rect 35514 451308 36134 476000
rect 39234 451308 39854 476000
rect 41794 451308 42414 476000
rect 42954 451308 43574 476000
rect 45514 451308 46134 476000
rect 49234 451308 49854 476000
rect 51794 451308 52414 476000
rect 52954 451308 53574 476000
rect 55514 451308 56134 476000
rect 59234 451308 59854 476000
rect 61794 451308 62414 476000
rect 62954 451308 63574 476000
rect 65514 451308 66134 476000
rect 69234 451308 69854 476000
rect 71794 451308 72414 476000
rect 72954 451308 73574 476000
rect 75514 451308 76134 476000
rect 79234 451308 79854 476000
rect 81794 451308 82414 476000
rect 82954 451308 83574 476000
rect 85514 451308 86134 476000
rect 89234 451308 89854 476000
rect 91794 451308 92414 476000
rect 92954 451308 93574 476000
rect 95514 451308 96134 476000
rect 99234 451308 99854 476000
rect 101794 451308 102414 476000
rect 102954 451308 103574 476000
rect 105514 451308 106134 476000
rect 109234 451308 109854 476000
rect 111794 451308 112414 476000
rect 112954 451308 113574 476000
rect 115514 451308 116134 476000
rect 119234 451308 119854 476000
rect 121794 451308 122414 476000
rect 122954 451308 123574 476000
rect 125514 451308 126134 476000
rect 129234 451308 129854 476000
rect 131794 451308 132414 476000
rect 132954 451308 133574 476000
rect 135514 451308 136134 476000
rect 139234 451308 139854 476000
rect 141794 451308 142414 476000
rect 142954 451308 143574 476000
rect 145514 451308 146134 476000
rect 149234 451308 149854 476000
rect 151794 451308 152414 476000
rect 152954 451308 153574 476000
rect 155514 451308 156134 476000
rect 159234 451308 159854 476000
rect 161794 451308 162414 476000
rect 162954 451308 163574 476000
rect 165514 451308 166134 476000
rect 29234 339308 29854 364000
rect 31794 339308 32414 364000
rect 32954 339308 33574 364000
rect 35514 339308 36134 364000
rect 39234 339308 39854 364000
rect 41794 339308 42414 364000
rect 42954 339308 43574 364000
rect 45514 339308 46134 364000
rect 49234 339308 49854 364000
rect 51794 339308 52414 364000
rect 52954 339308 53574 364000
rect 55514 339308 56134 364000
rect 59234 339308 59854 364000
rect 61794 339308 62414 364000
rect 62954 339308 63574 364000
rect 65514 339308 66134 364000
rect 69234 339308 69854 364000
rect 71794 339308 72414 364000
rect 72954 339308 73574 364000
rect 75514 339308 76134 364000
rect 79234 339308 79854 364000
rect 81794 339308 82414 364000
rect 82954 339308 83574 364000
rect 85514 339308 86134 364000
rect 89234 339308 89854 364000
rect 91794 339308 92414 364000
rect 92954 339308 93574 364000
rect 95514 339308 96134 364000
rect 99234 339308 99854 364000
rect 101794 339308 102414 364000
rect 102954 339308 103574 364000
rect 105514 339308 106134 364000
rect 109234 339308 109854 364000
rect 111794 339308 112414 364000
rect 112954 339308 113574 364000
rect 115514 339308 116134 364000
rect 119234 339308 119854 364000
rect 121794 339308 122414 364000
rect 122954 339308 123574 364000
rect 125514 339308 126134 364000
rect 129234 339308 129854 364000
rect 131794 339308 132414 364000
rect 132954 339308 133574 364000
rect 135514 339308 136134 364000
rect 139234 339308 139854 364000
rect 141794 339308 142414 364000
rect 142954 339308 143574 364000
rect 145514 339308 146134 364000
rect 149234 339308 149854 364000
rect 151794 339308 152414 364000
rect 152954 339308 153574 364000
rect 155514 339308 156134 364000
rect 159234 339308 159854 364000
rect 161794 339308 162414 364000
rect 162954 339308 163574 364000
rect 165514 339308 166134 364000
rect 29234 227308 29854 252000
rect 31794 227308 32414 252000
rect 32954 227308 33574 252000
rect 35514 227308 36134 252000
rect 39234 227308 39854 252000
rect 41794 227308 42414 252000
rect 42954 227308 43574 252000
rect 45514 227308 46134 252000
rect 49234 227308 49854 252000
rect 51794 227308 52414 252000
rect 52954 227308 53574 252000
rect 55514 227308 56134 252000
rect 59234 227308 59854 252000
rect 61794 227308 62414 252000
rect 62954 227308 63574 252000
rect 65514 227308 66134 252000
rect 69234 227308 69854 252000
rect 71794 227308 72414 252000
rect 72954 227308 73574 252000
rect 75514 227308 76134 252000
rect 79234 227308 79854 252000
rect 81794 227308 82414 252000
rect 82954 227308 83574 252000
rect 85514 227308 86134 252000
rect 89234 227308 89854 252000
rect 91794 227308 92414 252000
rect 92954 227308 93574 252000
rect 95514 227308 96134 252000
rect 99234 227308 99854 252000
rect 101794 227308 102414 252000
rect 102954 227308 103574 252000
rect 105514 227308 106134 252000
rect 109234 227308 109854 252000
rect 111794 227308 112414 252000
rect 112954 227308 113574 252000
rect 115514 227308 116134 252000
rect 119234 227308 119854 252000
rect 121794 227308 122414 252000
rect 122954 227308 123574 252000
rect 125514 227308 126134 252000
rect 129234 227308 129854 252000
rect 131794 227308 132414 252000
rect 132954 227308 133574 252000
rect 135514 227308 136134 252000
rect 139234 227308 139854 252000
rect 141794 227308 142414 252000
rect 142954 227308 143574 252000
rect 145514 227308 146134 252000
rect 149234 227308 149854 252000
rect 151794 227308 152414 252000
rect 152954 227308 153574 252000
rect 155514 227308 156134 252000
rect 159234 227308 159854 252000
rect 161794 227308 162414 252000
rect 162954 227308 163574 252000
rect 165514 227308 166134 252000
rect 29234 115308 29854 140000
rect 31794 115308 32414 140000
rect 32954 115308 33574 140000
rect 35514 115308 36134 140000
rect 39234 115308 39854 140000
rect 41794 115308 42414 140000
rect 42954 115308 43574 140000
rect 45514 115308 46134 140000
rect 49234 115308 49854 140000
rect 51794 115308 52414 140000
rect 52954 115308 53574 140000
rect 55514 115308 56134 140000
rect 59234 115308 59854 140000
rect 61794 115308 62414 140000
rect 62954 115308 63574 140000
rect 65514 115308 66134 140000
rect 69234 115308 69854 140000
rect 71794 115308 72414 140000
rect 72954 115308 73574 140000
rect 75514 115308 76134 140000
rect 79234 115308 79854 140000
rect 81794 115308 82414 140000
rect 82954 115308 83574 140000
rect 85514 115308 86134 140000
rect 89234 115308 89854 140000
rect 91794 115308 92414 140000
rect 92954 115308 93574 140000
rect 95514 115308 96134 140000
rect 99234 115308 99854 140000
rect 101794 115308 102414 140000
rect 102954 115308 103574 140000
rect 105514 115308 106134 140000
rect 109234 115308 109854 140000
rect 111794 115308 112414 140000
rect 112954 115308 113574 140000
rect 115514 115308 116134 140000
rect 119234 115308 119854 140000
rect 121794 115308 122414 140000
rect 122954 115308 123574 140000
rect 125514 115308 126134 140000
rect 129234 115308 129854 140000
rect 131794 115308 132414 140000
rect 132954 115308 133574 140000
rect 135514 115308 136134 140000
rect 139234 115308 139854 140000
rect 141794 115308 142414 140000
rect 142954 115308 143574 140000
rect 145514 115308 146134 140000
rect 149234 115308 149854 140000
rect 151794 115308 152414 140000
rect 152954 115308 153574 140000
rect 155514 115308 156134 140000
rect 159234 115308 159854 140000
rect 161794 115308 162414 140000
rect 162954 115308 163574 140000
rect 165514 115308 166134 140000
rect 29234 -5734 29854 28000
rect 31794 -1894 32414 28000
rect 32954 -7654 33574 28000
rect 35514 -3814 36134 28000
rect 39234 -5734 39854 28000
rect 41794 -1894 42414 28000
rect 42954 -7654 43574 28000
rect 45514 -3814 46134 28000
rect 49234 -5734 49854 28000
rect 51794 -1894 52414 28000
rect 52954 -7654 53574 28000
rect 55514 -3814 56134 28000
rect 59234 -5734 59854 28000
rect 61794 -1894 62414 28000
rect 62954 -7654 63574 28000
rect 65514 -3814 66134 28000
rect 69234 -5734 69854 28000
rect 71794 -1894 72414 28000
rect 72954 -7654 73574 28000
rect 75514 -3814 76134 28000
rect 79234 -5734 79854 28000
rect 81794 -1894 82414 28000
rect 82954 -7654 83574 28000
rect 85514 -3814 86134 28000
rect 89234 -5734 89854 28000
rect 91794 -1894 92414 28000
rect 92954 -7654 93574 28000
rect 95514 -3814 96134 28000
rect 99234 -5734 99854 28000
rect 101794 -1894 102414 28000
rect 102954 -7654 103574 28000
rect 105514 -3814 106134 28000
rect 109234 -5734 109854 28000
rect 111794 -1894 112414 28000
rect 112954 -7654 113574 28000
rect 115514 -3814 116134 28000
rect 119234 -5734 119854 28000
rect 121794 -1894 122414 28000
rect 122954 -7654 123574 28000
rect 125514 -3814 126134 28000
rect 129234 -5734 129854 28000
rect 131794 -1894 132414 28000
rect 132954 -7654 133574 28000
rect 135514 -3814 136134 28000
rect 139234 -5734 139854 28000
rect 141794 -1894 142414 28000
rect 142954 -7654 143574 28000
rect 145514 -3814 146134 28000
rect 149234 -5734 149854 28000
rect 151794 -1894 152414 28000
rect 152954 -7654 153574 28000
rect 155514 -3814 156134 28000
rect 159234 -5734 159854 28000
rect 161794 -1894 162414 28000
rect 162954 -7654 163574 28000
rect 165514 -3814 166134 28000
rect 169234 -5734 169854 709670
rect 171794 -1894 172414 705830
rect 172954 -7654 173574 711590
rect 175514 -3814 176134 707750
rect 179234 -5734 179854 709670
rect 181794 -1894 182414 705830
rect 182954 -7654 183574 711590
rect 185514 -3814 186134 707750
rect 189234 -5734 189854 709670
rect 191794 -1894 192414 705830
rect 192954 -7654 193574 711590
rect 195514 -3814 196134 707750
rect 199234 539308 199854 709670
rect 201794 539308 202414 705830
rect 202954 539308 203574 711590
rect 205514 539308 206134 707750
rect 209234 539308 209854 709670
rect 211794 539308 212414 705830
rect 212954 539308 213574 711590
rect 215514 539308 216134 707750
rect 219234 539308 219854 709670
rect 221794 539308 222414 705830
rect 222954 539308 223574 711590
rect 225514 539308 226134 707750
rect 229234 539308 229854 709670
rect 231794 539308 232414 705830
rect 232954 539308 233574 711590
rect 235514 539308 236134 707750
rect 239234 659500 239854 709670
rect 241794 659500 242414 705830
rect 242954 659500 243574 711590
rect 245514 659500 246134 707750
rect 249234 659500 249854 709670
rect 251794 659500 252414 705830
rect 252954 659500 253574 711590
rect 255514 659500 256134 707750
rect 259234 659500 259854 709670
rect 261794 659500 262414 705830
rect 262954 659500 263574 711590
rect 265514 659500 266134 707750
rect 269234 659500 269854 709670
rect 271794 659500 272414 705830
rect 272954 659500 273574 711590
rect 275514 659500 276134 707750
rect 279234 659500 279854 709670
rect 281794 659500 282414 705830
rect 282954 659500 283574 711590
rect 285514 659500 286134 707750
rect 289234 659500 289854 709670
rect 291794 659500 292414 705830
rect 292954 659500 293574 711590
rect 295514 659500 296134 707750
rect 299234 659500 299854 709670
rect 301794 659500 302414 705830
rect 302954 659500 303574 711590
rect 305514 659500 306134 707750
rect 309234 659500 309854 709670
rect 311794 659500 312414 705830
rect 312954 659500 313574 711590
rect 315514 659500 316134 707750
rect 319234 659500 319854 709670
rect 321794 659500 322414 705830
rect 322954 659500 323574 711590
rect 325514 659500 326134 707750
rect 329234 659500 329854 709670
rect 331794 659500 332414 705830
rect 332954 659500 333574 711590
rect 335514 659500 336134 707750
rect 239234 539308 239854 576000
rect 241794 539308 242414 576000
rect 242954 539308 243574 576000
rect 245514 539308 246134 576000
rect 249234 539308 249854 576000
rect 251794 539308 252414 576000
rect 252954 539308 253574 576000
rect 255514 539308 256134 576000
rect 259234 539308 259854 576000
rect 261794 539308 262414 576000
rect 262954 539308 263574 576000
rect 265514 539308 266134 576000
rect 269234 539308 269854 576000
rect 271794 539308 272414 576000
rect 272954 539308 273574 576000
rect 275514 539308 276134 576000
rect 279234 539308 279854 576000
rect 281794 539308 282414 576000
rect 282954 539308 283574 576000
rect 285514 539308 286134 576000
rect 289234 539308 289854 576000
rect 291794 539308 292414 576000
rect 292954 539308 293574 576000
rect 295514 539308 296134 576000
rect 299234 539308 299854 576000
rect 301794 539308 302414 576000
rect 302954 539308 303574 576000
rect 305514 539308 306134 576000
rect 309234 539308 309854 576000
rect 311794 539308 312414 576000
rect 312954 539308 313574 576000
rect 315514 539308 316134 576000
rect 319234 539308 319854 576000
rect 321794 539308 322414 576000
rect 322954 539308 323574 576000
rect 325514 539308 326134 576000
rect 329234 539308 329854 576000
rect 331794 539308 332414 576000
rect 332954 539308 333574 576000
rect 335514 539308 336134 576000
rect 199234 421162 199854 452000
rect 201794 421162 202414 452000
rect 202954 421162 203574 452000
rect 205514 421162 206134 452000
rect 209234 421162 209854 452000
rect 211794 421162 212414 452000
rect 212954 421162 213574 452000
rect 215514 421162 216134 452000
rect 219234 421162 219854 452000
rect 221794 421162 222414 452000
rect 222954 421162 223574 452000
rect 225514 421162 226134 452000
rect 229234 421162 229854 452000
rect 231794 421162 232414 452000
rect 232954 421162 233574 452000
rect 235514 421162 236134 452000
rect 239234 421162 239854 452000
rect 241794 421162 242414 452000
rect 242954 421162 243574 452000
rect 245514 421162 246134 452000
rect 249234 421162 249854 452000
rect 251794 421162 252414 452000
rect 252954 421162 253574 452000
rect 255514 421162 256134 452000
rect 259234 421162 259854 452000
rect 261794 421162 262414 452000
rect 262954 421162 263574 452000
rect 265514 421162 266134 452000
rect 269234 421162 269854 452000
rect 271794 421162 272414 452000
rect 272954 421162 273574 452000
rect 275514 421162 276134 452000
rect 279234 421162 279854 452000
rect 281794 421162 282414 452000
rect 282954 421162 283574 452000
rect 285514 421162 286134 452000
rect 289234 421162 289854 452000
rect 291794 421162 292414 452000
rect 292954 421162 293574 452000
rect 295514 421162 296134 452000
rect 299234 421162 299854 452000
rect 301794 421162 302414 452000
rect 302954 421162 303574 452000
rect 305514 421162 306134 452000
rect 309234 421162 309854 452000
rect 311794 421162 312414 452000
rect 312954 421162 313574 452000
rect 315514 421162 316134 452000
rect 319234 421162 319854 452000
rect 321794 421162 322414 452000
rect 322954 421162 323574 452000
rect 325514 421162 326134 452000
rect 329234 421162 329854 452000
rect 331794 421162 332414 452000
rect 332954 421162 333574 452000
rect 335514 421162 336134 452000
rect 339234 421162 339854 709670
rect 341794 421162 342414 705830
rect 342954 421162 343574 711590
rect 345514 421162 346134 707750
rect 349234 421162 349854 709670
rect 351794 421162 352414 705830
rect 352954 421162 353574 711590
rect 355514 421162 356134 707750
rect 359234 421162 359854 709670
rect 361794 421162 362414 705830
rect 362954 421162 363574 711590
rect 365514 421162 366134 707750
rect 369234 421162 369854 709670
rect 371794 421162 372414 705830
rect 372954 421162 373574 711590
rect 375514 421162 376134 707750
rect 379234 421162 379854 709670
rect 381794 421162 382414 705830
rect 382954 421162 383574 711590
rect 385514 421162 386134 707750
rect 389234 421162 389854 709670
rect 391794 421162 392414 705830
rect 392954 421162 393574 711590
rect 395514 421162 396134 707750
rect 399234 421162 399854 709670
rect 401794 421162 402414 705830
rect 402954 421162 403574 711590
rect 405514 421162 406134 707750
rect 409234 659500 409854 709670
rect 411794 659500 412414 705830
rect 412954 659500 413574 711590
rect 415514 659500 416134 707750
rect 419234 659500 419854 709670
rect 421794 659500 422414 705830
rect 422954 659500 423574 711590
rect 425514 659500 426134 707750
rect 429234 659500 429854 709670
rect 431794 659500 432414 705830
rect 432954 659500 433574 711590
rect 435514 659500 436134 707750
rect 439234 659500 439854 709670
rect 441794 659500 442414 705830
rect 442954 659500 443574 711590
rect 445514 659500 446134 707750
rect 449234 659500 449854 709670
rect 451794 659500 452414 705830
rect 452954 659500 453574 711590
rect 455514 659500 456134 707750
rect 459234 659500 459854 709670
rect 461794 659500 462414 705830
rect 462954 659500 463574 711590
rect 465514 659500 466134 707750
rect 469234 659500 469854 709670
rect 471794 659500 472414 705830
rect 472954 659500 473574 711590
rect 475514 659500 476134 707750
rect 479234 659500 479854 709670
rect 481794 659500 482414 705830
rect 482954 659500 483574 711590
rect 485514 659500 486134 707750
rect 489234 659500 489854 709670
rect 491794 659500 492414 705830
rect 492954 659500 493574 711590
rect 495514 659500 496134 707750
rect 499234 659500 499854 709670
rect 501794 659500 502414 705830
rect 502954 659500 503574 711590
rect 505514 659500 506134 707750
rect 409234 539308 409854 576000
rect 411794 539308 412414 576000
rect 412954 539308 413574 576000
rect 415514 539308 416134 576000
rect 419234 539308 419854 576000
rect 421794 539308 422414 576000
rect 422954 539308 423574 576000
rect 425514 539308 426134 576000
rect 429234 539308 429854 576000
rect 431794 539308 432414 576000
rect 432954 539308 433574 576000
rect 435514 539308 436134 576000
rect 439234 539308 439854 576000
rect 441794 539308 442414 576000
rect 442954 539308 443574 576000
rect 445514 539308 446134 576000
rect 449234 539308 449854 576000
rect 451794 539308 452414 576000
rect 452954 539308 453574 576000
rect 455514 539308 456134 576000
rect 459234 539308 459854 576000
rect 461794 539308 462414 576000
rect 462954 539308 463574 576000
rect 465514 539308 466134 576000
rect 469234 539308 469854 576000
rect 471794 539308 472414 576000
rect 472954 539308 473574 576000
rect 475514 539308 476134 576000
rect 479234 539308 479854 576000
rect 481794 539308 482414 576000
rect 482954 539308 483574 576000
rect 485514 539308 486134 576000
rect 489234 539308 489854 576000
rect 491794 539308 492414 576000
rect 492954 539308 493574 576000
rect 495514 539308 496134 576000
rect 499234 539308 499854 576000
rect 501794 539308 502414 576000
rect 502954 539308 503574 576000
rect 505514 539308 506134 576000
rect 509234 539308 509854 709670
rect 511794 539308 512414 705830
rect 512954 539308 513574 711590
rect 515514 539308 516134 707750
rect 519234 539308 519854 709670
rect 521794 539308 522414 705830
rect 522954 539308 523574 711590
rect 525514 539308 526134 707750
rect 529234 539308 529854 709670
rect 531794 539308 532414 705830
rect 532954 539308 533574 711590
rect 535514 539308 536134 707750
rect 539234 539308 539854 709670
rect 541794 539308 542414 705830
rect 542954 539308 543574 711590
rect 545514 539308 546134 707750
rect 409234 421162 409854 452000
rect 411794 421162 412414 452000
rect 412954 421162 413574 452000
rect 415514 421162 416134 452000
rect 419234 421162 419854 452000
rect 421794 421162 422414 452000
rect 422954 421162 423574 452000
rect 425514 421162 426134 452000
rect 429234 421162 429854 452000
rect 431794 421162 432414 452000
rect 432954 421162 433574 452000
rect 435514 421162 436134 452000
rect 439234 421162 439854 452000
rect 441794 421162 442414 452000
rect 442954 421162 443574 452000
rect 445514 421162 446134 452000
rect 449234 421162 449854 452000
rect 451794 421162 452414 452000
rect 452954 421162 453574 452000
rect 455514 421162 456134 452000
rect 459234 421162 459854 452000
rect 461794 421162 462414 452000
rect 462954 421162 463574 452000
rect 465514 421162 466134 452000
rect 469234 421162 469854 452000
rect 471794 421162 472414 452000
rect 472954 421162 473574 452000
rect 475514 421162 476134 452000
rect 479234 421162 479854 452000
rect 481794 421162 482414 452000
rect 482954 421162 483574 452000
rect 485514 421162 486134 452000
rect 489234 421162 489854 452000
rect 491794 421162 492414 452000
rect 492954 421162 493574 452000
rect 495514 421162 496134 452000
rect 499234 421162 499854 452000
rect 501794 421162 502414 452000
rect 502954 421162 503574 452000
rect 505514 421162 506134 452000
rect 509234 421162 509854 452000
rect 511794 421162 512414 452000
rect 512954 421162 513574 452000
rect 515514 421162 516134 452000
rect 519234 421162 519854 452000
rect 521794 421162 522414 452000
rect 522954 421162 523574 452000
rect 525514 421162 526134 452000
rect 529234 421162 529854 452000
rect 531794 421162 532414 452000
rect 532954 421162 533574 452000
rect 535514 421162 536134 452000
rect 539234 421162 539854 452000
rect 541794 421162 542414 452000
rect 542954 421162 543574 452000
rect 545514 421162 546134 452000
rect 549234 421162 549854 709670
rect 551794 421162 552414 705830
rect 552954 421162 553574 711590
rect 555514 421162 556134 707750
rect 199234 -5734 199854 58000
rect 201794 -1894 202414 58000
rect 202954 -7654 203574 58000
rect 205514 -3814 206134 58000
rect 209234 -5734 209854 58000
rect 211794 -1894 212414 58000
rect 212954 -7654 213574 58000
rect 215514 -3814 216134 58000
rect 219234 -5734 219854 58000
rect 221794 -1894 222414 58000
rect 222954 -7654 223574 58000
rect 225514 -3814 226134 58000
rect 229234 -5734 229854 58000
rect 231794 -1894 232414 58000
rect 232954 -7654 233574 58000
rect 235514 -3814 236134 58000
rect 239234 -5734 239854 58000
rect 241794 -1894 242414 58000
rect 242954 -7654 243574 58000
rect 245514 -3814 246134 58000
rect 249234 -5734 249854 58000
rect 251794 -1894 252414 58000
rect 252954 -7654 253574 58000
rect 255514 -3814 256134 58000
rect 259234 -5734 259854 58000
rect 261794 -1894 262414 58000
rect 262954 -7654 263574 58000
rect 265514 -3814 266134 58000
rect 269234 -5734 269854 58000
rect 271794 -1894 272414 58000
rect 272954 -7654 273574 58000
rect 275514 -3814 276134 58000
rect 279234 -5734 279854 58000
rect 281794 -1894 282414 58000
rect 282954 -7654 283574 58000
rect 285514 -3814 286134 58000
rect 289234 -5734 289854 58000
rect 291794 -1894 292414 58000
rect 292954 -7654 293574 58000
rect 295514 -3814 296134 58000
rect 299234 -5734 299854 58000
rect 301794 -1894 302414 58000
rect 302954 -7654 303574 58000
rect 305514 -3814 306134 58000
rect 309234 -5734 309854 58000
rect 311794 -1894 312414 58000
rect 312954 -7654 313574 58000
rect 315514 -3814 316134 58000
rect 319234 -5734 319854 58000
rect 321794 -1894 322414 58000
rect 322954 -7654 323574 58000
rect 325514 -3814 326134 58000
rect 329234 -5734 329854 58000
rect 331794 -1894 332414 58000
rect 332954 -7654 333574 58000
rect 335514 -3814 336134 58000
rect 339234 -5734 339854 58000
rect 341794 -1894 342414 58000
rect 342954 -7654 343574 58000
rect 345514 -3814 346134 58000
rect 349234 -5734 349854 58000
rect 351794 -1894 352414 58000
rect 352954 -7654 353574 58000
rect 355514 -3814 356134 58000
rect 359234 -5734 359854 58000
rect 361794 -1894 362414 58000
rect 362954 -7654 363574 58000
rect 365514 -3814 366134 58000
rect 369234 -5734 369854 58000
rect 371794 -1894 372414 58000
rect 372954 -7654 373574 58000
rect 375514 -3814 376134 58000
rect 379234 -5734 379854 58000
rect 381794 -1894 382414 58000
rect 382954 -7654 383574 58000
rect 385514 -3814 386134 58000
rect 389234 -5734 389854 58000
rect 391794 -1894 392414 58000
rect 392954 -7654 393574 58000
rect 395514 -3814 396134 58000
rect 399234 -5734 399854 58000
rect 401794 -1894 402414 58000
rect 402954 -7654 403574 58000
rect 405514 -3814 406134 58000
rect 409234 -5734 409854 58000
rect 411794 -1894 412414 58000
rect 412954 -7654 413574 58000
rect 415514 -3814 416134 58000
rect 419234 -5734 419854 58000
rect 421794 -1894 422414 58000
rect 422954 -7654 423574 58000
rect 425514 -3814 426134 58000
rect 429234 -5734 429854 58000
rect 431794 -1894 432414 58000
rect 432954 -7654 433574 58000
rect 435514 -3814 436134 58000
rect 439234 -5734 439854 58000
rect 441794 -1894 442414 58000
rect 442954 -7654 443574 58000
rect 445514 -3814 446134 58000
rect 449234 -5734 449854 58000
rect 451794 -1894 452414 58000
rect 452954 -7654 453574 58000
rect 455514 -3814 456134 58000
rect 459234 -5734 459854 58000
rect 461794 -1894 462414 58000
rect 462954 -7654 463574 58000
rect 465514 -3814 466134 58000
rect 469234 -5734 469854 58000
rect 471794 -1894 472414 58000
rect 472954 -7654 473574 58000
rect 475514 -3814 476134 58000
rect 479234 -5734 479854 58000
rect 481794 -1894 482414 58000
rect 482954 -7654 483574 58000
rect 485514 -3814 486134 58000
rect 489234 -5734 489854 58000
rect 491794 -1894 492414 58000
rect 492954 -7654 493574 58000
rect 495514 -3814 496134 58000
rect 499234 -5734 499854 58000
rect 501794 -1894 502414 58000
rect 502954 -7654 503574 58000
rect 505514 -3814 506134 58000
rect 509234 -5734 509854 58000
rect 511794 -1894 512414 58000
rect 512954 -7654 513574 58000
rect 515514 -3814 516134 58000
rect 519234 -5734 519854 58000
rect 521794 -1894 522414 58000
rect 522954 -7654 523574 58000
rect 525514 -3814 526134 58000
rect 529234 -5734 529854 58000
rect 531794 -1894 532414 58000
rect 532954 -7654 533574 58000
rect 535514 -3814 536134 58000
rect 539234 -5734 539854 58000
rect 541794 -1894 542414 58000
rect 542954 -7654 543574 58000
rect 545514 -3814 546134 58000
rect 549234 -5734 549854 58000
rect 551794 -1894 552414 58000
rect 552954 -7654 553574 58000
rect 555514 -3814 556134 58000
rect 559234 -5734 559854 709670
rect 561794 -1894 562414 705830
rect 562954 -7654 563574 711590
rect 565514 -3814 566134 707750
rect 569234 -5734 569854 709670
rect 571794 -1894 572414 705830
rect 572954 -7654 573574 711590
rect 575514 -3814 576134 707750
rect 579234 -5734 579854 709670
rect 581794 -1894 582414 705830
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 30124 675228 31714 700637
rect 32494 675228 32874 700637
rect 33654 675228 35434 700637
rect 36214 675228 39154 700637
rect 39934 675228 41714 700637
rect 42494 675228 42874 700637
rect 43654 675228 45434 700637
rect 46214 675228 49154 700637
rect 49934 675228 51714 700637
rect 52494 675228 52874 700637
rect 53654 675228 55434 700637
rect 56214 675228 59154 700637
rect 59934 675228 61714 700637
rect 62494 675228 62874 700637
rect 63654 675228 65434 700637
rect 66214 675228 69154 700637
rect 69934 675228 71714 700637
rect 72494 675228 72874 700637
rect 73654 675228 75434 700637
rect 76214 675228 79154 700637
rect 79934 675228 81714 700637
rect 82494 675228 82874 700637
rect 83654 675228 85434 700637
rect 86214 675228 89154 700637
rect 89934 675228 91714 700637
rect 92494 675228 92874 700637
rect 93654 675228 95434 700637
rect 96214 675228 99154 700637
rect 99934 675228 101714 700637
rect 102494 675228 102874 700637
rect 103654 675228 105434 700637
rect 106214 675228 109154 700637
rect 109934 675228 111714 700637
rect 112494 675228 112874 700637
rect 113654 675228 115434 700637
rect 116214 675228 119154 700637
rect 119934 675228 121714 700637
rect 122494 675228 122874 700637
rect 123654 675228 125434 700637
rect 126214 675228 129154 700637
rect 129934 675228 131714 700637
rect 132494 675228 132874 700637
rect 133654 675228 135434 700637
rect 136214 675228 139154 700637
rect 139934 675228 141714 700637
rect 142494 675228 142874 700637
rect 143654 675228 145434 700637
rect 146214 675228 149154 700637
rect 149934 675228 151714 700637
rect 152494 675228 152874 700637
rect 153654 675228 155434 700637
rect 156214 675228 159154 700637
rect 159934 675228 161714 700637
rect 162494 675228 162874 700637
rect 163654 675228 165434 700637
rect 166214 675228 169154 700637
rect 30124 588080 169154 675228
rect 30124 563228 31714 588080
rect 32494 563228 32874 588080
rect 33654 563228 35434 588080
rect 36214 563228 39154 588080
rect 39934 563228 41714 588080
rect 42494 563228 42874 588080
rect 43654 563228 45434 588080
rect 46214 563228 49154 588080
rect 49934 563228 51714 588080
rect 52494 563228 52874 588080
rect 53654 563228 55434 588080
rect 56214 563228 59154 588080
rect 59934 563228 61714 588080
rect 62494 563228 62874 588080
rect 63654 563228 65434 588080
rect 66214 563228 69154 588080
rect 69934 563228 71714 588080
rect 72494 563228 72874 588080
rect 73654 563228 75434 588080
rect 76214 563228 79154 588080
rect 79934 563228 81714 588080
rect 82494 563228 82874 588080
rect 83654 563228 85434 588080
rect 86214 563228 89154 588080
rect 89934 563228 91714 588080
rect 92494 563228 92874 588080
rect 93654 563228 95434 588080
rect 96214 563228 99154 588080
rect 99934 563228 101714 588080
rect 102494 563228 102874 588080
rect 103654 563228 105434 588080
rect 106214 563228 109154 588080
rect 109934 563228 111714 588080
rect 112494 563228 112874 588080
rect 113654 563228 115434 588080
rect 116214 563228 119154 588080
rect 119934 563228 121714 588080
rect 122494 563228 122874 588080
rect 123654 563228 125434 588080
rect 126214 563228 129154 588080
rect 129934 563228 131714 588080
rect 132494 563228 132874 588080
rect 133654 563228 135434 588080
rect 136214 563228 139154 588080
rect 139934 563228 141714 588080
rect 142494 563228 142874 588080
rect 143654 563228 145434 588080
rect 146214 563228 149154 588080
rect 149934 563228 151714 588080
rect 152494 563228 152874 588080
rect 153654 563228 155434 588080
rect 156214 563228 159154 588080
rect 159934 563228 161714 588080
rect 162494 563228 162874 588080
rect 163654 563228 165434 588080
rect 166214 563228 169154 588080
rect 30124 476080 169154 563228
rect 30124 451228 31714 476080
rect 32494 451228 32874 476080
rect 33654 451228 35434 476080
rect 36214 451228 39154 476080
rect 39934 451228 41714 476080
rect 42494 451228 42874 476080
rect 43654 451228 45434 476080
rect 46214 451228 49154 476080
rect 49934 451228 51714 476080
rect 52494 451228 52874 476080
rect 53654 451228 55434 476080
rect 56214 451228 59154 476080
rect 59934 451228 61714 476080
rect 62494 451228 62874 476080
rect 63654 451228 65434 476080
rect 66214 451228 69154 476080
rect 69934 451228 71714 476080
rect 72494 451228 72874 476080
rect 73654 451228 75434 476080
rect 76214 451228 79154 476080
rect 79934 451228 81714 476080
rect 82494 451228 82874 476080
rect 83654 451228 85434 476080
rect 86214 451228 89154 476080
rect 89934 451228 91714 476080
rect 92494 451228 92874 476080
rect 93654 451228 95434 476080
rect 96214 451228 99154 476080
rect 99934 451228 101714 476080
rect 102494 451228 102874 476080
rect 103654 451228 105434 476080
rect 106214 451228 109154 476080
rect 109934 451228 111714 476080
rect 112494 451228 112874 476080
rect 113654 451228 115434 476080
rect 116214 451228 119154 476080
rect 119934 451228 121714 476080
rect 122494 451228 122874 476080
rect 123654 451228 125434 476080
rect 126214 451228 129154 476080
rect 129934 451228 131714 476080
rect 132494 451228 132874 476080
rect 133654 451228 135434 476080
rect 136214 451228 139154 476080
rect 139934 451228 141714 476080
rect 142494 451228 142874 476080
rect 143654 451228 145434 476080
rect 146214 451228 149154 476080
rect 149934 451228 151714 476080
rect 152494 451228 152874 476080
rect 153654 451228 155434 476080
rect 156214 451228 159154 476080
rect 159934 451228 161714 476080
rect 162494 451228 162874 476080
rect 163654 451228 165434 476080
rect 166214 451228 169154 476080
rect 30124 364080 169154 451228
rect 30124 339228 31714 364080
rect 32494 339228 32874 364080
rect 33654 339228 35434 364080
rect 36214 339228 39154 364080
rect 39934 339228 41714 364080
rect 42494 339228 42874 364080
rect 43654 339228 45434 364080
rect 46214 339228 49154 364080
rect 49934 339228 51714 364080
rect 52494 339228 52874 364080
rect 53654 339228 55434 364080
rect 56214 339228 59154 364080
rect 59934 339228 61714 364080
rect 62494 339228 62874 364080
rect 63654 339228 65434 364080
rect 66214 339228 69154 364080
rect 69934 339228 71714 364080
rect 72494 339228 72874 364080
rect 73654 339228 75434 364080
rect 76214 339228 79154 364080
rect 79934 339228 81714 364080
rect 82494 339228 82874 364080
rect 83654 339228 85434 364080
rect 86214 339228 89154 364080
rect 89934 339228 91714 364080
rect 92494 339228 92874 364080
rect 93654 339228 95434 364080
rect 96214 339228 99154 364080
rect 99934 339228 101714 364080
rect 102494 339228 102874 364080
rect 103654 339228 105434 364080
rect 106214 339228 109154 364080
rect 109934 339228 111714 364080
rect 112494 339228 112874 364080
rect 113654 339228 115434 364080
rect 116214 339228 119154 364080
rect 119934 339228 121714 364080
rect 122494 339228 122874 364080
rect 123654 339228 125434 364080
rect 126214 339228 129154 364080
rect 129934 339228 131714 364080
rect 132494 339228 132874 364080
rect 133654 339228 135434 364080
rect 136214 339228 139154 364080
rect 139934 339228 141714 364080
rect 142494 339228 142874 364080
rect 143654 339228 145434 364080
rect 146214 339228 149154 364080
rect 149934 339228 151714 364080
rect 152494 339228 152874 364080
rect 153654 339228 155434 364080
rect 156214 339228 159154 364080
rect 159934 339228 161714 364080
rect 162494 339228 162874 364080
rect 163654 339228 165434 364080
rect 166214 339228 169154 364080
rect 30124 252080 169154 339228
rect 30124 227228 31714 252080
rect 32494 227228 32874 252080
rect 33654 227228 35434 252080
rect 36214 227228 39154 252080
rect 39934 227228 41714 252080
rect 42494 227228 42874 252080
rect 43654 227228 45434 252080
rect 46214 227228 49154 252080
rect 49934 227228 51714 252080
rect 52494 227228 52874 252080
rect 53654 227228 55434 252080
rect 56214 227228 59154 252080
rect 59934 227228 61714 252080
rect 62494 227228 62874 252080
rect 63654 227228 65434 252080
rect 66214 227228 69154 252080
rect 69934 227228 71714 252080
rect 72494 227228 72874 252080
rect 73654 227228 75434 252080
rect 76214 227228 79154 252080
rect 79934 227228 81714 252080
rect 82494 227228 82874 252080
rect 83654 227228 85434 252080
rect 86214 227228 89154 252080
rect 89934 227228 91714 252080
rect 92494 227228 92874 252080
rect 93654 227228 95434 252080
rect 96214 227228 99154 252080
rect 99934 227228 101714 252080
rect 102494 227228 102874 252080
rect 103654 227228 105434 252080
rect 106214 227228 109154 252080
rect 109934 227228 111714 252080
rect 112494 227228 112874 252080
rect 113654 227228 115434 252080
rect 116214 227228 119154 252080
rect 119934 227228 121714 252080
rect 122494 227228 122874 252080
rect 123654 227228 125434 252080
rect 126214 227228 129154 252080
rect 129934 227228 131714 252080
rect 132494 227228 132874 252080
rect 133654 227228 135434 252080
rect 136214 227228 139154 252080
rect 139934 227228 141714 252080
rect 142494 227228 142874 252080
rect 143654 227228 145434 252080
rect 146214 227228 149154 252080
rect 149934 227228 151714 252080
rect 152494 227228 152874 252080
rect 153654 227228 155434 252080
rect 156214 227228 159154 252080
rect 159934 227228 161714 252080
rect 162494 227228 162874 252080
rect 163654 227228 165434 252080
rect 166214 227228 169154 252080
rect 30124 140080 169154 227228
rect 30124 115228 31714 140080
rect 32494 115228 32874 140080
rect 33654 115228 35434 140080
rect 36214 115228 39154 140080
rect 39934 115228 41714 140080
rect 42494 115228 42874 140080
rect 43654 115228 45434 140080
rect 46214 115228 49154 140080
rect 49934 115228 51714 140080
rect 52494 115228 52874 140080
rect 53654 115228 55434 140080
rect 56214 115228 59154 140080
rect 59934 115228 61714 140080
rect 62494 115228 62874 140080
rect 63654 115228 65434 140080
rect 66214 115228 69154 140080
rect 69934 115228 71714 140080
rect 72494 115228 72874 140080
rect 73654 115228 75434 140080
rect 76214 115228 79154 140080
rect 79934 115228 81714 140080
rect 82494 115228 82874 140080
rect 83654 115228 85434 140080
rect 86214 115228 89154 140080
rect 89934 115228 91714 140080
rect 92494 115228 92874 140080
rect 93654 115228 95434 140080
rect 96214 115228 99154 140080
rect 99934 115228 101714 140080
rect 102494 115228 102874 140080
rect 103654 115228 105434 140080
rect 106214 115228 109154 140080
rect 109934 115228 111714 140080
rect 112494 115228 112874 140080
rect 113654 115228 115434 140080
rect 116214 115228 119154 140080
rect 119934 115228 121714 140080
rect 122494 115228 122874 140080
rect 123654 115228 125434 140080
rect 126214 115228 129154 140080
rect 129934 115228 131714 140080
rect 132494 115228 132874 140080
rect 133654 115228 135434 140080
rect 136214 115228 139154 140080
rect 139934 115228 141714 140080
rect 142494 115228 142874 140080
rect 143654 115228 145434 140080
rect 146214 115228 149154 140080
rect 149934 115228 151714 140080
rect 152494 115228 152874 140080
rect 153654 115228 155434 140080
rect 156214 115228 159154 140080
rect 159934 115228 161714 140080
rect 162494 115228 162874 140080
rect 163654 115228 165434 140080
rect 166214 115228 169154 140080
rect 30124 28080 169154 115228
rect 30124 5611 31714 28080
rect 32494 5611 32874 28080
rect 33654 5611 35434 28080
rect 36214 5611 39154 28080
rect 39934 5611 41714 28080
rect 42494 5611 42874 28080
rect 43654 5611 45434 28080
rect 46214 5611 49154 28080
rect 49934 5611 51714 28080
rect 52494 5611 52874 28080
rect 53654 5611 55434 28080
rect 56214 5611 59154 28080
rect 59934 5611 61714 28080
rect 62494 5611 62874 28080
rect 63654 5611 65434 28080
rect 66214 5611 69154 28080
rect 69934 5611 71714 28080
rect 72494 5611 72874 28080
rect 73654 5611 75434 28080
rect 76214 5611 79154 28080
rect 79934 5611 81714 28080
rect 82494 5611 82874 28080
rect 83654 5611 85434 28080
rect 86214 5611 89154 28080
rect 89934 5611 91714 28080
rect 92494 5611 92874 28080
rect 93654 5611 95434 28080
rect 96214 5611 99154 28080
rect 99934 5611 101714 28080
rect 102494 5611 102874 28080
rect 103654 5611 105434 28080
rect 106214 5611 109154 28080
rect 109934 5611 111714 28080
rect 112494 5611 112874 28080
rect 113654 5611 115434 28080
rect 116214 5611 119154 28080
rect 119934 5611 121714 28080
rect 122494 5611 122874 28080
rect 123654 5611 125434 28080
rect 126214 5611 129154 28080
rect 129934 5611 131714 28080
rect 132494 5611 132874 28080
rect 133654 5611 135434 28080
rect 136214 5611 139154 28080
rect 139934 5611 141714 28080
rect 142494 5611 142874 28080
rect 143654 5611 145434 28080
rect 146214 5611 149154 28080
rect 149934 5611 151714 28080
rect 152494 5611 152874 28080
rect 153654 5611 155434 28080
rect 156214 5611 159154 28080
rect 159934 5611 161714 28080
rect 162494 5611 162874 28080
rect 163654 5611 165434 28080
rect 166214 5611 169154 28080
rect 169934 5611 171714 700637
rect 172494 5611 172874 700637
rect 173654 5611 175434 700637
rect 176214 5611 179154 700637
rect 179934 5611 181714 700637
rect 182494 5611 182874 700637
rect 183654 5611 185434 700637
rect 186214 5611 189154 700637
rect 189934 5611 191714 700637
rect 192494 5611 192874 700637
rect 193654 5611 195434 700637
rect 196214 539228 199154 700637
rect 199934 539228 201714 700637
rect 202494 539228 202874 700637
rect 203654 539228 205434 700637
rect 206214 539228 209154 700637
rect 209934 539228 211714 700637
rect 212494 539228 212874 700637
rect 213654 539228 215434 700637
rect 216214 539228 219154 700637
rect 219934 539228 221714 700637
rect 222494 539228 222874 700637
rect 223654 539228 225434 700637
rect 226214 539228 229154 700637
rect 229934 539228 231714 700637
rect 232494 539228 232874 700637
rect 233654 539228 235434 700637
rect 236214 659420 239154 700637
rect 239934 659420 241714 700637
rect 242494 659420 242874 700637
rect 243654 659420 245434 700637
rect 246214 659420 249154 700637
rect 249934 659420 251714 700637
rect 252494 659420 252874 700637
rect 253654 659420 255434 700637
rect 256214 659420 259154 700637
rect 259934 659420 261714 700637
rect 262494 659420 262874 700637
rect 263654 659420 265434 700637
rect 266214 659420 269154 700637
rect 269934 659420 271714 700637
rect 272494 659420 272874 700637
rect 273654 659420 275434 700637
rect 276214 659420 279154 700637
rect 279934 659420 281714 700637
rect 282494 659420 282874 700637
rect 283654 659420 285434 700637
rect 286214 659420 289154 700637
rect 289934 659420 291714 700637
rect 292494 659420 292874 700637
rect 293654 659420 295434 700637
rect 296214 659420 299154 700637
rect 299934 659420 301714 700637
rect 302494 659420 302874 700637
rect 303654 659420 305434 700637
rect 306214 659420 309154 700637
rect 309934 659420 311714 700637
rect 312494 659420 312874 700637
rect 313654 659420 315434 700637
rect 316214 659420 319154 700637
rect 319934 659420 321714 700637
rect 322494 659420 322874 700637
rect 323654 659420 325434 700637
rect 326214 659420 329154 700637
rect 329934 659420 331714 700637
rect 332494 659420 332874 700637
rect 333654 659420 335434 700637
rect 336214 659420 339154 700637
rect 236214 576080 339154 659420
rect 236214 539228 239154 576080
rect 239934 539228 241714 576080
rect 242494 539228 242874 576080
rect 243654 539228 245434 576080
rect 246214 539228 249154 576080
rect 249934 539228 251714 576080
rect 252494 539228 252874 576080
rect 253654 539228 255434 576080
rect 256214 539228 259154 576080
rect 259934 539228 261714 576080
rect 262494 539228 262874 576080
rect 263654 539228 265434 576080
rect 266214 539228 269154 576080
rect 269934 539228 271714 576080
rect 272494 539228 272874 576080
rect 273654 539228 275434 576080
rect 276214 539228 279154 576080
rect 279934 539228 281714 576080
rect 282494 539228 282874 576080
rect 283654 539228 285434 576080
rect 286214 539228 289154 576080
rect 289934 539228 291714 576080
rect 292494 539228 292874 576080
rect 293654 539228 295434 576080
rect 296214 539228 299154 576080
rect 299934 539228 301714 576080
rect 302494 539228 302874 576080
rect 303654 539228 305434 576080
rect 306214 539228 309154 576080
rect 309934 539228 311714 576080
rect 312494 539228 312874 576080
rect 313654 539228 315434 576080
rect 316214 539228 319154 576080
rect 319934 539228 321714 576080
rect 322494 539228 322874 576080
rect 323654 539228 325434 576080
rect 326214 539228 329154 576080
rect 329934 539228 331714 576080
rect 332494 539228 332874 576080
rect 333654 539228 335434 576080
rect 336214 539228 339154 576080
rect 196214 452080 339154 539228
rect 196214 421082 199154 452080
rect 199934 421082 201714 452080
rect 202494 421082 202874 452080
rect 203654 421082 205434 452080
rect 206214 421082 209154 452080
rect 209934 421082 211714 452080
rect 212494 421082 212874 452080
rect 213654 421082 215434 452080
rect 216214 421082 219154 452080
rect 219934 421082 221714 452080
rect 222494 421082 222874 452080
rect 223654 421082 225434 452080
rect 226214 421082 229154 452080
rect 229934 421082 231714 452080
rect 232494 421082 232874 452080
rect 233654 421082 235434 452080
rect 236214 421082 239154 452080
rect 239934 421082 241714 452080
rect 242494 421082 242874 452080
rect 243654 421082 245434 452080
rect 246214 421082 249154 452080
rect 249934 421082 251714 452080
rect 252494 421082 252874 452080
rect 253654 421082 255434 452080
rect 256214 421082 259154 452080
rect 259934 421082 261714 452080
rect 262494 421082 262874 452080
rect 263654 421082 265434 452080
rect 266214 421082 269154 452080
rect 269934 421082 271714 452080
rect 272494 421082 272874 452080
rect 273654 421082 275434 452080
rect 276214 421082 279154 452080
rect 279934 421082 281714 452080
rect 282494 421082 282874 452080
rect 283654 421082 285434 452080
rect 286214 421082 289154 452080
rect 289934 421082 291714 452080
rect 292494 421082 292874 452080
rect 293654 421082 295434 452080
rect 296214 421082 299154 452080
rect 299934 421082 301714 452080
rect 302494 421082 302874 452080
rect 303654 421082 305434 452080
rect 306214 421082 309154 452080
rect 309934 421082 311714 452080
rect 312494 421082 312874 452080
rect 313654 421082 315434 452080
rect 316214 421082 319154 452080
rect 319934 421082 321714 452080
rect 322494 421082 322874 452080
rect 323654 421082 325434 452080
rect 326214 421082 329154 452080
rect 329934 421082 331714 452080
rect 332494 421082 332874 452080
rect 333654 421082 335434 452080
rect 336214 421082 339154 452080
rect 339934 421082 341714 700637
rect 342494 421082 342874 700637
rect 343654 421082 345434 700637
rect 346214 421082 349154 700637
rect 349934 421082 351714 700637
rect 352494 421082 352874 700637
rect 353654 421082 355434 700637
rect 356214 421082 359154 700637
rect 359934 421082 361714 700637
rect 362494 421082 362874 700637
rect 363654 421082 365434 700637
rect 366214 421082 369154 700637
rect 369934 421082 371714 700637
rect 372494 421082 372874 700637
rect 373654 421082 375434 700637
rect 376214 421082 379154 700637
rect 379934 421082 381714 700637
rect 382494 421082 382874 700637
rect 383654 421082 385434 700637
rect 386214 421082 389154 700637
rect 389934 421082 391714 700637
rect 392494 421082 392874 700637
rect 393654 421082 395434 700637
rect 396214 421082 399154 700637
rect 399934 421082 401714 700637
rect 402494 421082 402874 700637
rect 403654 421082 405434 700637
rect 406214 659420 409154 700637
rect 409934 659420 411714 700637
rect 412494 659420 412874 700637
rect 413654 659420 415434 700637
rect 416214 659420 419154 700637
rect 419934 659420 421714 700637
rect 422494 659420 422874 700637
rect 423654 659420 425434 700637
rect 426214 659420 429154 700637
rect 429934 659420 431714 700637
rect 432494 659420 432874 700637
rect 433654 659420 435434 700637
rect 436214 659420 439154 700637
rect 439934 659420 441714 700637
rect 442494 659420 442874 700637
rect 443654 659420 445434 700637
rect 446214 659420 449154 700637
rect 449934 659420 451714 700637
rect 452494 659420 452874 700637
rect 453654 659420 455434 700637
rect 456214 659420 459154 700637
rect 459934 659420 461714 700637
rect 462494 659420 462874 700637
rect 463654 659420 465434 700637
rect 466214 659420 469154 700637
rect 469934 659420 471714 700637
rect 472494 659420 472874 700637
rect 473654 659420 475434 700637
rect 476214 659420 479154 700637
rect 479934 659420 481714 700637
rect 482494 659420 482874 700637
rect 483654 659420 485434 700637
rect 486214 659420 489154 700637
rect 489934 659420 491714 700637
rect 492494 659420 492874 700637
rect 493654 659420 495434 700637
rect 496214 659420 499154 700637
rect 499934 659420 501714 700637
rect 502494 659420 502874 700637
rect 503654 659420 505434 700637
rect 506214 659420 509154 700637
rect 406214 576080 509154 659420
rect 406214 539228 409154 576080
rect 409934 539228 411714 576080
rect 412494 539228 412874 576080
rect 413654 539228 415434 576080
rect 416214 539228 419154 576080
rect 419934 539228 421714 576080
rect 422494 539228 422874 576080
rect 423654 539228 425434 576080
rect 426214 539228 429154 576080
rect 429934 539228 431714 576080
rect 432494 539228 432874 576080
rect 433654 539228 435434 576080
rect 436214 539228 439154 576080
rect 439934 539228 441714 576080
rect 442494 539228 442874 576080
rect 443654 539228 445434 576080
rect 446214 539228 449154 576080
rect 449934 539228 451714 576080
rect 452494 539228 452874 576080
rect 453654 539228 455434 576080
rect 456214 539228 459154 576080
rect 459934 539228 461714 576080
rect 462494 539228 462874 576080
rect 463654 539228 465434 576080
rect 466214 539228 469154 576080
rect 469934 539228 471714 576080
rect 472494 539228 472874 576080
rect 473654 539228 475434 576080
rect 476214 539228 479154 576080
rect 479934 539228 481714 576080
rect 482494 539228 482874 576080
rect 483654 539228 485434 576080
rect 486214 539228 489154 576080
rect 489934 539228 491714 576080
rect 492494 539228 492874 576080
rect 493654 539228 495434 576080
rect 496214 539228 499154 576080
rect 499934 539228 501714 576080
rect 502494 539228 502874 576080
rect 503654 539228 505434 576080
rect 506214 539228 509154 576080
rect 509934 539228 511714 700637
rect 512494 539228 512874 700637
rect 513654 539228 515434 700637
rect 516214 539228 519154 700637
rect 519934 539228 521714 700637
rect 522494 539228 522874 700637
rect 523654 539228 525434 700637
rect 526214 539228 529154 700637
rect 529934 539228 531714 700637
rect 532494 539228 532874 700637
rect 533654 539228 535434 700637
rect 536214 539228 539154 700637
rect 539934 539228 541714 700637
rect 542494 539228 542874 700637
rect 543654 539228 545434 700637
rect 546214 539228 546496 700637
rect 406214 452080 546496 539228
rect 406214 421082 409154 452080
rect 409934 421082 411714 452080
rect 412494 421082 412874 452080
rect 413654 421082 415434 452080
rect 416214 421082 419154 452080
rect 419934 421082 421714 452080
rect 422494 421082 422874 452080
rect 423654 421082 425434 452080
rect 426214 421082 429154 452080
rect 429934 421082 431714 452080
rect 432494 421082 432874 452080
rect 433654 421082 435434 452080
rect 436214 421082 439154 452080
rect 439934 421082 441714 452080
rect 442494 421082 442874 452080
rect 443654 421082 445434 452080
rect 446214 421082 449154 452080
rect 449934 421082 451714 452080
rect 452494 421082 452874 452080
rect 453654 421082 455434 452080
rect 456214 421082 459154 452080
rect 459934 421082 461714 452080
rect 462494 421082 462874 452080
rect 463654 421082 465434 452080
rect 466214 421082 469154 452080
rect 469934 421082 471714 452080
rect 472494 421082 472874 452080
rect 473654 421082 475434 452080
rect 476214 421082 479154 452080
rect 479934 421082 481714 452080
rect 482494 421082 482874 452080
rect 483654 421082 485434 452080
rect 486214 421082 489154 452080
rect 489934 421082 491714 452080
rect 492494 421082 492874 452080
rect 493654 421082 495434 452080
rect 496214 421082 499154 452080
rect 499934 421082 501714 452080
rect 502494 421082 502874 452080
rect 503654 421082 505434 452080
rect 506214 421082 509154 452080
rect 509934 421082 511714 452080
rect 512494 421082 512874 452080
rect 513654 421082 515434 452080
rect 516214 421082 519154 452080
rect 519934 421082 521714 452080
rect 522494 421082 522874 452080
rect 523654 421082 525434 452080
rect 526214 421082 529154 452080
rect 529934 421082 531714 452080
rect 532494 421082 532874 452080
rect 533654 421082 535434 452080
rect 536214 421082 539154 452080
rect 539934 421082 541714 452080
rect 542494 421082 542874 452080
rect 543654 421082 545434 452080
rect 546214 421082 546496 452080
rect 196214 58080 546496 421082
rect 196214 5611 199154 58080
rect 199934 5611 201714 58080
rect 202494 5611 202874 58080
rect 203654 5611 205434 58080
rect 206214 5611 209154 58080
rect 209934 5611 211714 58080
rect 212494 5611 212874 58080
rect 213654 5611 215434 58080
rect 216214 5611 219154 58080
rect 219934 5611 221714 58080
rect 222494 5611 222874 58080
rect 223654 5611 225434 58080
rect 226214 5611 229154 58080
rect 229934 5611 231714 58080
rect 232494 5611 232874 58080
rect 233654 5611 235434 58080
rect 236214 5611 239154 58080
rect 239934 5611 241714 58080
rect 242494 5611 242874 58080
rect 243654 5611 245434 58080
rect 246214 5611 249154 58080
rect 249934 5611 251714 58080
rect 252494 5611 252874 58080
rect 253654 5611 255434 58080
rect 256214 5611 259154 58080
rect 259934 5611 261714 58080
rect 262494 5611 262874 58080
rect 263654 5611 265434 58080
rect 266214 5611 269154 58080
rect 269934 5611 271714 58080
rect 272494 5611 272874 58080
rect 273654 5611 275434 58080
rect 276214 5611 279154 58080
rect 279934 5611 281714 58080
rect 282494 5611 282874 58080
rect 283654 5611 285434 58080
rect 286214 5611 289154 58080
rect 289934 5611 291714 58080
rect 292494 5611 292874 58080
rect 293654 5611 295434 58080
rect 296214 5611 299154 58080
rect 299934 5611 301714 58080
rect 302494 5611 302874 58080
rect 303654 5611 305434 58080
rect 306214 5611 309154 58080
rect 309934 5611 311714 58080
rect 312494 5611 312874 58080
rect 313654 5611 315434 58080
rect 316214 5611 319154 58080
rect 319934 5611 321714 58080
rect 322494 5611 322874 58080
rect 323654 5611 325434 58080
rect 326214 5611 329154 58080
rect 329934 5611 331714 58080
rect 332494 5611 332874 58080
rect 333654 5611 335434 58080
rect 336214 5611 339154 58080
rect 339934 5611 341714 58080
rect 342494 5611 342874 58080
rect 343654 5611 345434 58080
rect 346214 5611 349154 58080
rect 349934 5611 351714 58080
rect 352494 5611 352874 58080
rect 353654 5611 355434 58080
rect 356214 5611 359154 58080
rect 359934 5611 361714 58080
rect 362494 5611 362874 58080
rect 363654 5611 365434 58080
rect 366214 5611 369154 58080
rect 369934 5611 371714 58080
rect 372494 5611 372874 58080
rect 373654 5611 375434 58080
rect 376214 5611 379154 58080
rect 379934 5611 381714 58080
rect 382494 5611 382874 58080
rect 383654 5611 385434 58080
rect 386214 5611 389154 58080
rect 389934 5611 391714 58080
rect 392494 5611 392874 58080
rect 393654 5611 395434 58080
rect 396214 5611 399154 58080
rect 399934 5611 401714 58080
rect 402494 5611 402874 58080
rect 403654 5611 405434 58080
rect 406214 5611 409154 58080
rect 409934 5611 411714 58080
rect 412494 5611 412874 58080
rect 413654 5611 415434 58080
rect 416214 5611 419154 58080
rect 419934 5611 421714 58080
rect 422494 5611 422874 58080
rect 423654 5611 425434 58080
rect 426214 5611 429154 58080
rect 429934 5611 431714 58080
rect 432494 5611 432874 58080
rect 433654 5611 435434 58080
rect 436214 5611 439154 58080
rect 439934 5611 441714 58080
rect 442494 5611 442874 58080
rect 443654 5611 445434 58080
rect 446214 5611 449154 58080
rect 449934 5611 451714 58080
rect 452494 5611 452874 58080
rect 453654 5611 455434 58080
rect 456214 5611 459154 58080
rect 459934 5611 461714 58080
rect 462494 5611 462874 58080
rect 463654 5611 465434 58080
rect 466214 5611 469154 58080
rect 469934 5611 471714 58080
rect 472494 5611 472874 58080
rect 473654 5611 475434 58080
rect 476214 5611 479154 58080
rect 479934 5611 481714 58080
rect 482494 5611 482874 58080
rect 483654 5611 485434 58080
rect 486214 5611 489154 58080
rect 489934 5611 491714 58080
rect 492494 5611 492874 58080
rect 493654 5611 495434 58080
rect 496214 5611 499154 58080
rect 499934 5611 501714 58080
rect 502494 5611 502874 58080
rect 503654 5611 505434 58080
rect 506214 5611 509154 58080
rect 509934 5611 511714 58080
rect 512494 5611 512874 58080
rect 513654 5611 515434 58080
rect 516214 5611 519154 58080
rect 519934 5611 521714 58080
rect 522494 5611 522874 58080
rect 523654 5611 525434 58080
rect 526214 5611 529154 58080
rect 529934 5611 531714 58080
rect 532494 5611 532874 58080
rect 533654 5611 535434 58080
rect 536214 5611 539154 58080
rect 539934 5611 541714 58080
rect 542494 5611 542874 58080
rect 543654 5611 545434 58080
rect 546214 5611 546496 58080
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -6806 700306 590730 700926
rect -4886 696586 588810 697206
rect -8726 694026 592650 694646
rect -2966 692866 586890 693486
rect -6806 690306 590730 690926
rect -4886 686586 588810 687206
rect -8726 684026 592650 684646
rect -2966 682866 586890 683486
rect -6806 680306 590730 680926
rect -4886 676586 588810 677206
rect -8726 674026 592650 674646
rect -2966 672866 586890 673486
rect -6806 670306 590730 670926
rect -4886 666586 588810 667206
rect -8726 664026 592650 664646
rect -2966 662866 586890 663486
rect -6806 660306 590730 660926
rect -4886 656586 588810 657206
rect -8726 654026 592650 654646
rect -2966 652866 586890 653486
rect -6806 650306 590730 650926
rect -4886 646586 588810 647206
rect -8726 644026 592650 644646
rect -2966 642866 586890 643486
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -8726 634026 592650 634646
rect -2966 632866 586890 633486
rect -6806 630306 590730 630926
rect -4886 626586 588810 627206
rect -8726 624026 592650 624646
rect -2966 622866 586890 623486
rect -6806 620306 590730 620926
rect -4886 616586 588810 617206
rect -8726 614026 592650 614646
rect -2966 612866 586890 613486
rect -6806 610306 590730 610926
rect -4886 606586 588810 607206
rect -8726 604026 592650 604646
rect -2966 602866 586890 603486
rect -6806 600306 590730 600926
rect -4886 596586 588810 597206
rect -8726 594026 592650 594646
rect -2966 592866 586890 593486
rect -6806 590306 590730 590926
rect -4886 586586 588810 587206
rect -8726 584026 592650 584646
rect -2966 582866 586890 583486
rect -6806 580306 590730 580926
rect -4886 576586 588810 577206
rect -8726 574026 592650 574646
rect -2966 572866 586890 573486
rect -6806 570306 590730 570926
rect -4886 566586 588810 567206
rect -8726 564026 592650 564646
rect -2966 562866 586890 563486
rect -6806 560306 590730 560926
rect -4886 556586 588810 557206
rect -8726 554026 592650 554646
rect -2966 552866 586890 553486
rect -6806 550306 590730 550926
rect -4886 546586 588810 547206
rect -8726 544026 592650 544646
rect -2966 542866 586890 543486
rect -6806 540306 590730 540926
rect -4886 536586 588810 537206
rect -8726 534026 592650 534646
rect -2966 532866 586890 533486
rect -6806 530306 590730 530926
rect -4886 526586 588810 527206
rect -8726 524026 592650 524646
rect -2966 522866 586890 523486
rect -6806 520306 590730 520926
rect -4886 516586 588810 517206
rect -8726 514026 592650 514646
rect -2966 512866 586890 513486
rect -6806 510306 590730 510926
rect -4886 506586 588810 507206
rect -8726 504026 592650 504646
rect -2966 502866 586890 503486
rect -6806 500306 590730 500926
rect -4886 496586 588810 497206
rect -8726 494026 592650 494646
rect -2966 492866 586890 493486
rect -6806 490306 590730 490926
rect -4886 486586 588810 487206
rect -8726 484026 592650 484646
rect -2966 482866 586890 483486
rect -6806 480306 590730 480926
rect -4886 476586 588810 477206
rect -8726 474026 592650 474646
rect -2966 472866 586890 473486
rect -6806 470306 590730 470926
rect -4886 466586 588810 467206
rect -8726 464026 592650 464646
rect -2966 462866 586890 463486
rect -6806 460306 590730 460926
rect -4886 456586 588810 457206
rect -8726 454026 592650 454646
rect -2966 452866 586890 453486
rect -6806 450306 590730 450926
rect -4886 446586 588810 447206
rect -8726 444026 592650 444646
rect -2966 442866 586890 443486
rect -6806 440306 590730 440926
rect -4886 436586 588810 437206
rect -8726 434026 592650 434646
rect -2966 432866 586890 433486
rect -6806 430306 590730 430926
rect -4886 426586 588810 427206
rect -8726 424026 592650 424646
rect -2966 422866 586890 423486
rect -6806 420306 590730 420926
rect -4886 416586 588810 417206
rect -8726 414026 592650 414646
rect -2966 412866 586890 413486
rect -6806 410306 590730 410926
rect -4886 406586 588810 407206
rect -8726 404026 592650 404646
rect -2966 402866 586890 403486
rect -6806 400306 590730 400926
rect -4886 396586 588810 397206
rect -8726 394026 592650 394646
rect -2966 392866 586890 393486
rect -6806 390306 590730 390926
rect -4886 386586 588810 387206
rect -8726 384026 592650 384646
rect -2966 382866 586890 383486
rect -6806 380306 590730 380926
rect -4886 376586 588810 377206
rect -8726 374026 592650 374646
rect -2966 372866 586890 373486
rect -6806 370306 590730 370926
rect -4886 366586 588810 367206
rect -8726 364026 592650 364646
rect -2966 362866 586890 363486
rect -6806 360306 590730 360926
rect -4886 356586 588810 357206
rect -8726 354026 592650 354646
rect -2966 352866 586890 353486
rect -6806 350306 590730 350926
rect -4886 346586 588810 347206
rect -8726 344026 592650 344646
rect -2966 342866 586890 343486
rect -6806 340306 590730 340926
rect -4886 336586 588810 337206
rect -8726 334026 592650 334646
rect -2966 332866 586890 333486
rect -6806 330306 590730 330926
rect -4886 326586 588810 327206
rect -8726 324026 592650 324646
rect -2966 322866 586890 323486
rect -6806 320306 590730 320926
rect -4886 316586 588810 317206
rect -8726 314026 592650 314646
rect -2966 312866 586890 313486
rect -6806 310306 590730 310926
rect -4886 306586 588810 307206
rect -8726 304026 592650 304646
rect -2966 302866 586890 303486
rect -6806 300306 590730 300926
rect -4886 296586 588810 297206
rect -8726 294026 592650 294646
rect -2966 292866 586890 293486
rect -6806 290306 590730 290926
rect -4886 286586 588810 287206
rect -8726 284026 592650 284646
rect -2966 282866 586890 283486
rect -6806 280306 590730 280926
rect -4886 276586 588810 277206
rect -8726 274026 592650 274646
rect -2966 272866 586890 273486
rect -6806 270306 590730 270926
rect -4886 266586 588810 267206
rect -8726 264026 592650 264646
rect -2966 262866 586890 263486
rect -6806 260306 590730 260926
rect -4886 256586 588810 257206
rect -8726 254026 592650 254646
rect -2966 252866 586890 253486
rect -6806 250306 590730 250926
rect -4886 246586 588810 247206
rect -8726 244026 592650 244646
rect -2966 242866 586890 243486
rect -6806 240306 590730 240926
rect -4886 236586 588810 237206
rect -8726 234026 592650 234646
rect -2966 232866 586890 233486
rect -6806 230306 590730 230926
rect -4886 226586 588810 227206
rect -8726 224026 592650 224646
rect -2966 222866 586890 223486
rect -6806 220306 590730 220926
rect -4886 216586 588810 217206
rect -8726 214026 592650 214646
rect -2966 212866 586890 213486
rect -6806 210306 590730 210926
rect -4886 206586 588810 207206
rect -8726 204026 592650 204646
rect -2966 202866 586890 203486
rect -6806 200306 590730 200926
rect -4886 196586 588810 197206
rect -8726 194026 592650 194646
rect -2966 192866 586890 193486
rect -6806 190306 590730 190926
rect -4886 186586 588810 187206
rect -8726 184026 592650 184646
rect -2966 182866 586890 183486
rect -6806 180306 590730 180926
rect -4886 176586 588810 177206
rect -8726 174026 592650 174646
rect -2966 172866 586890 173486
rect -6806 170306 590730 170926
rect -4886 166586 588810 167206
rect -8726 164026 592650 164646
rect -2966 162866 586890 163486
rect -6806 160306 590730 160926
rect -4886 156586 588810 157206
rect -8726 154026 592650 154646
rect -2966 152866 586890 153486
rect -6806 150306 590730 150926
rect -4886 146586 588810 147206
rect -8726 144026 592650 144646
rect -2966 142866 586890 143486
rect -6806 140306 590730 140926
rect -4886 136586 588810 137206
rect -8726 134026 592650 134646
rect -2966 132866 586890 133486
rect -6806 130306 590730 130926
rect -4886 126586 588810 127206
rect -8726 124026 592650 124646
rect -2966 122866 586890 123486
rect -6806 120306 590730 120926
rect -4886 116586 588810 117206
rect -8726 114026 592650 114646
rect -2966 112866 586890 113486
rect -6806 110306 590730 110926
rect -4886 106586 588810 107206
rect -8726 104026 592650 104646
rect -2966 102866 586890 103486
rect -6806 100306 590730 100926
rect -4886 96586 588810 97206
rect -8726 94026 592650 94646
rect -2966 92866 586890 93486
rect -6806 90306 590730 90926
rect -4886 86586 588810 87206
rect -8726 84026 592650 84646
rect -2966 82866 586890 83486
rect -6806 80306 590730 80926
rect -4886 76586 588810 77206
rect -8726 74026 592650 74646
rect -2966 72866 586890 73486
rect -6806 70306 590730 70926
rect -4886 66586 588810 67206
rect -8726 64026 592650 64646
rect -2966 62866 586890 63486
rect -6806 60306 590730 60926
rect -4886 56586 588810 57206
rect -8726 54026 592650 54646
rect -2966 52866 586890 53486
rect -6806 50306 590730 50926
rect -4886 46586 588810 47206
rect -8726 44026 592650 44646
rect -2966 42866 586890 43486
rect -6806 40306 590730 40926
rect -4886 36586 588810 37206
rect -8726 34026 592650 34646
rect -2966 32866 586890 33486
rect -6806 30306 590730 30926
rect -4886 26586 588810 27206
rect -8726 24026 592650 24646
rect -2966 22866 586890 23486
rect -6806 20306 590730 20926
rect -4886 16586 588810 17206
rect -8726 14026 592650 14646
rect -2966 12866 586890 13486
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 22866 586890 23486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 42866 586890 43486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 62866 586890 63486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 82866 586890 83486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 102866 586890 103486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 122866 586890 123486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 142866 586890 143486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 162866 586890 163486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 202866 586890 203486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 222866 586890 223486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 242866 586890 243486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 262866 586890 263486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 282866 586890 283486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 302866 586890 303486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 322866 586890 323486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 342866 586890 343486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 382866 586890 383486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 402866 586890 403486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 422866 586890 423486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 442866 586890 443486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 462866 586890 463486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 482866 586890 483486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 502866 586890 503486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 522866 586890 523486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 562866 586890 563486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 582866 586890 583486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 602866 586890 603486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 622866 586890 623486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 642866 586890 643486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 662866 586890 663486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 682866 586890 683486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 41794 -1894 42414 28000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 -1894 62414 28000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 -1894 82414 28000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 -1894 102414 28000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 -1894 122414 28000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 -1894 142414 28000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 -1894 162414 28000 6 vccd1
port 532 nsew power input
rlabel metal4 s 201794 -1894 202414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 221794 -1894 222414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 -1894 242414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 -1894 262414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 -1894 282414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 -1894 302414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 -1894 322414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 341794 -1894 342414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 -1894 362414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 381794 -1894 382414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 401794 -1894 402414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 -1894 422414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 441794 -1894 442414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 -1894 462414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 -1894 482414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 -1894 502414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 521794 -1894 522414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 -1894 542414 58000 6 vccd1
port 532 nsew power input
rlabel metal4 s 41794 115308 42414 140000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 115308 62414 140000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 115308 82414 140000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 115308 102414 140000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 115308 122414 140000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 115308 142414 140000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 115308 162414 140000 6 vccd1
port 532 nsew power input
rlabel metal4 s 41794 227308 42414 252000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 227308 62414 252000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 227308 82414 252000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 227308 102414 252000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 227308 122414 252000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 227308 142414 252000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 227308 162414 252000 6 vccd1
port 532 nsew power input
rlabel metal4 s 41794 339308 42414 364000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 339308 62414 364000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 339308 82414 364000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 339308 102414 364000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 339308 122414 364000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 339308 142414 364000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 339308 162414 364000 6 vccd1
port 532 nsew power input
rlabel metal4 s 201794 421162 202414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 221794 421162 222414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 421162 242414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 421162 262414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 421162 282414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 421162 302414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 421162 322414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 421162 422414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 441794 421162 442414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 421162 462414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 421162 482414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 421162 502414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 521794 421162 522414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 421162 542414 452000 6 vccd1
port 532 nsew power input
rlabel metal4 s 41794 451308 42414 476000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 451308 62414 476000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 451308 82414 476000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 451308 102414 476000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 451308 122414 476000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 451308 142414 476000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 451308 162414 476000 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 539308 242414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 539308 262414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 539308 282414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 539308 302414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 539308 322414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 539308 422414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 441794 539308 442414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 539308 462414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 539308 482414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 539308 502414 576000 6 vccd1
port 532 nsew power input
rlabel metal4 s 41794 563308 42414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 563308 62414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 563308 82414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 563308 102414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 563308 122414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 563308 142414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 563308 162414 588000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 21794 -1894 22414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 41794 675308 42414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 61794 675308 62414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 81794 675308 82414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 101794 675308 102414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 121794 675308 122414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 141794 675308 142414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 161794 675308 162414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 201794 539308 202414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 221794 539308 222414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 241794 659500 242414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 261794 659500 262414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 281794 659500 282414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 301794 659500 302414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 321794 659500 322414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 341794 421162 342414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 421162 362414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 381794 421162 382414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 401794 421162 402414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 421794 659500 422414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 441794 659500 442414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 461794 659500 462414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 481794 659500 482414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 501794 659500 502414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 521794 539308 522414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 539308 542414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 561794 -1894 562414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 581794 -1894 582414 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 26586 588810 27206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 46586 588810 47206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 66586 588810 67206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 86586 588810 87206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 106586 588810 107206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 126586 588810 127206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 146586 588810 147206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 166586 588810 167206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 206586 588810 207206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 226586 588810 227206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 246586 588810 247206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 266586 588810 267206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 286586 588810 287206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 306586 588810 307206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 326586 588810 327206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 346586 588810 347206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 386586 588810 387206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 406586 588810 407206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 426586 588810 427206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 446586 588810 447206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 466586 588810 467206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 486586 588810 487206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 506586 588810 507206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 526586 588810 527206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 566586 588810 567206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 586586 588810 587206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 606586 588810 607206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 626586 588810 627206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 646586 588810 647206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 666586 588810 667206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 686586 588810 687206 6 vccd2
port 533 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 45514 -3814 46134 28000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 -3814 66134 28000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 -3814 86134 28000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 -3814 106134 28000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 -3814 126134 28000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 -3814 146134 28000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 -3814 166134 28000 6 vccd2
port 533 nsew power input
rlabel metal4 s 205514 -3814 206134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 225514 -3814 226134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 -3814 246134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 -3814 266134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 -3814 286134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 -3814 306134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 325514 -3814 326134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 345514 -3814 346134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 -3814 366134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 385514 -3814 386134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 405514 -3814 406134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 -3814 426134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 445514 -3814 446134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 -3814 466134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 -3814 486134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 -3814 506134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 525514 -3814 526134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 545514 -3814 546134 58000 6 vccd2
port 533 nsew power input
rlabel metal4 s 45514 115308 46134 140000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 115308 66134 140000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 115308 86134 140000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 115308 106134 140000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 115308 126134 140000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 115308 146134 140000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 115308 166134 140000 6 vccd2
port 533 nsew power input
rlabel metal4 s 45514 227308 46134 252000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 227308 66134 252000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 227308 86134 252000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 227308 106134 252000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 227308 126134 252000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 227308 146134 252000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 227308 166134 252000 6 vccd2
port 533 nsew power input
rlabel metal4 s 45514 339308 46134 364000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 339308 66134 364000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 339308 86134 364000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 339308 106134 364000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 339308 126134 364000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 339308 146134 364000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 339308 166134 364000 6 vccd2
port 533 nsew power input
rlabel metal4 s 205514 421162 206134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 225514 421162 226134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 421162 246134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 421162 266134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 421162 286134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 421162 306134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 325514 421162 326134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 421162 426134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 445514 421162 446134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 421162 466134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 421162 486134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 421162 506134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 525514 421162 526134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 545514 421162 546134 452000 6 vccd2
port 533 nsew power input
rlabel metal4 s 45514 451308 46134 476000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 451308 66134 476000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 451308 86134 476000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 451308 106134 476000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 451308 126134 476000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 451308 146134 476000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 451308 166134 476000 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 539308 246134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 539308 266134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 539308 286134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 539308 306134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 325514 539308 326134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 539308 426134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 445514 539308 446134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 539308 466134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 539308 486134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 539308 506134 576000 6 vccd2
port 533 nsew power input
rlabel metal4 s 45514 563308 46134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 563308 66134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 563308 86134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 563308 106134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 563308 126134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 563308 146134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 563308 166134 588000 6 vccd2
port 533 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 25514 -3814 26134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 45514 675308 46134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 65514 675308 66134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 85514 675308 86134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 105514 675308 106134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 125514 675308 126134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 145514 675308 146134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 165514 675308 166134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 205514 539308 206134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 225514 539308 226134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 245514 659500 246134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 265514 659500 266134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 285514 659500 286134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 305514 659500 306134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 325514 659500 326134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 345514 421162 346134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 421162 366134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 385514 421162 386134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 405514 421162 406134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 425514 659500 426134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 445514 659500 446134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 465514 659500 466134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 485514 659500 486134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 505514 659500 506134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 525514 539308 526134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 545514 539308 546134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 565514 -3814 566134 707750 6 vccd2
port 533 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 30306 590730 30926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 50306 590730 50926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 70306 590730 70926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 90306 590730 90926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 110306 590730 110926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 130306 590730 130926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 150306 590730 150926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 170306 590730 170926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 210306 590730 210926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 230306 590730 230926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 250306 590730 250926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 270306 590730 270926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 290306 590730 290926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 310306 590730 310926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 330306 590730 330926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 350306 590730 350926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 390306 590730 390926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 410306 590730 410926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 430306 590730 430926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 450306 590730 450926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 470306 590730 470926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 490306 590730 490926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 510306 590730 510926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 530306 590730 530926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 570306 590730 570926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 590306 590730 590926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 610306 590730 610926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 630306 590730 630926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 650306 590730 650926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 670306 590730 670926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 690306 590730 690926 6 vdda1
port 534 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 29234 -5734 29854 28000 6 vdda1
port 534 nsew power input
rlabel metal4 s 49234 -5734 49854 28000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 -5734 69854 28000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 -5734 89854 28000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 -5734 109854 28000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 -5734 129854 28000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 -5734 149854 28000 6 vdda1
port 534 nsew power input
rlabel metal4 s 209234 -5734 209854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 229234 -5734 229854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 -5734 249854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 -5734 269854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 -5734 289854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 -5734 309854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 329234 -5734 329854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 349234 -5734 349854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 -5734 369854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 389234 -5734 389854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 -5734 409854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 -5734 429854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 -5734 449854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 -5734 469854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 -5734 489854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 509234 -5734 509854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 529234 -5734 529854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 549234 -5734 549854 58000 6 vdda1
port 534 nsew power input
rlabel metal4 s 29234 115308 29854 140000 6 vdda1
port 534 nsew power input
rlabel metal4 s 49234 115308 49854 140000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 115308 69854 140000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 115308 89854 140000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 115308 109854 140000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 115308 129854 140000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 115308 149854 140000 6 vdda1
port 534 nsew power input
rlabel metal4 s 29234 227308 29854 252000 6 vdda1
port 534 nsew power input
rlabel metal4 s 49234 227308 49854 252000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 227308 69854 252000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 227308 89854 252000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 227308 109854 252000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 227308 129854 252000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 227308 149854 252000 6 vdda1
port 534 nsew power input
rlabel metal4 s 29234 339308 29854 364000 6 vdda1
port 534 nsew power input
rlabel metal4 s 49234 339308 49854 364000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 339308 69854 364000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 339308 89854 364000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 339308 109854 364000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 339308 129854 364000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 339308 149854 364000 6 vdda1
port 534 nsew power input
rlabel metal4 s 209234 421162 209854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 229234 421162 229854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 421162 249854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 421162 269854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 421162 289854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 421162 309854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 329234 421162 329854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 421162 409854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 421162 429854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 421162 449854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 421162 469854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 421162 489854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 509234 421162 509854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 529234 421162 529854 452000 6 vdda1
port 534 nsew power input
rlabel metal4 s 29234 451308 29854 476000 6 vdda1
port 534 nsew power input
rlabel metal4 s 49234 451308 49854 476000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 451308 69854 476000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 451308 89854 476000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 451308 109854 476000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 451308 129854 476000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 451308 149854 476000 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 539308 249854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 539308 269854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 539308 289854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 539308 309854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 329234 539308 329854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 539308 409854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 539308 429854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 539308 449854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 539308 469854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 539308 489854 576000 6 vdda1
port 534 nsew power input
rlabel metal4 s 29234 563308 29854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 49234 563308 49854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 563308 69854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 563308 89854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 563308 109854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 563308 129854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 563308 149854 588000 6 vdda1
port 534 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 29234 675308 29854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 49234 675308 49854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 69234 675308 69854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 89234 675308 89854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 109234 675308 109854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 129234 675308 129854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 149234 675308 149854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 169234 -5734 169854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 209234 539308 209854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 229234 539308 229854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 249234 659500 249854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 269234 659500 269854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 289234 659500 289854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 309234 659500 309854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 329234 659500 329854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 349234 421162 349854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 421162 369854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 389234 421162 389854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 409234 659500 409854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 429234 659500 429854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 449234 659500 449854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 469234 659500 469854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 489234 659500 489854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 509234 539308 509854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 529234 539308 529854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 549234 421162 549854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 569234 -5734 569854 709670 6 vdda1
port 534 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 34026 592650 34646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 54026 592650 54646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 74026 592650 74646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 94026 592650 94646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 114026 592650 114646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 134026 592650 134646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 154026 592650 154646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 174026 592650 174646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 214026 592650 214646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 234026 592650 234646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 254026 592650 254646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 274026 592650 274646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 294026 592650 294646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 314026 592650 314646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 334026 592650 334646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 354026 592650 354646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 394026 592650 394646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 414026 592650 414646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 434026 592650 434646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 454026 592650 454646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 474026 592650 474646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 494026 592650 494646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 514026 592650 514646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 534026 592650 534646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 574026 592650 574646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 594026 592650 594646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 614026 592650 614646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 634026 592650 634646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 654026 592650 654646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 674026 592650 674646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 694026 592650 694646 6 vdda2
port 535 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 32954 -7654 33574 28000 6 vdda2
port 535 nsew power input
rlabel metal4 s 52954 -7654 53574 28000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 -7654 73574 28000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 -7654 93574 28000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 -7654 113574 28000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 -7654 133574 28000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 -7654 153574 28000 6 vdda2
port 535 nsew power input
rlabel metal4 s 212954 -7654 213574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 232954 -7654 233574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 -7654 253574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 -7654 273574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 -7654 293574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 -7654 313574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 332954 -7654 333574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 352954 -7654 353574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 -7654 373574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 392954 -7654 393574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 -7654 413574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 -7654 433574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 -7654 453574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 -7654 473574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 -7654 493574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 512954 -7654 513574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 532954 -7654 533574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 552954 -7654 553574 58000 6 vdda2
port 535 nsew power input
rlabel metal4 s 32954 115308 33574 140000 6 vdda2
port 535 nsew power input
rlabel metal4 s 52954 115308 53574 140000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 115308 73574 140000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 115308 93574 140000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 115308 113574 140000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 115308 133574 140000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 115308 153574 140000 6 vdda2
port 535 nsew power input
rlabel metal4 s 32954 227308 33574 252000 6 vdda2
port 535 nsew power input
rlabel metal4 s 52954 227308 53574 252000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 227308 73574 252000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 227308 93574 252000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 227308 113574 252000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 227308 133574 252000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 227308 153574 252000 6 vdda2
port 535 nsew power input
rlabel metal4 s 32954 339308 33574 364000 6 vdda2
port 535 nsew power input
rlabel metal4 s 52954 339308 53574 364000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 339308 73574 364000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 339308 93574 364000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 339308 113574 364000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 339308 133574 364000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 339308 153574 364000 6 vdda2
port 535 nsew power input
rlabel metal4 s 212954 421162 213574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 232954 421162 233574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 421162 253574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 421162 273574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 421162 293574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 421162 313574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 332954 421162 333574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 421162 413574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 421162 433574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 421162 453574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 421162 473574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 421162 493574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 512954 421162 513574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 532954 421162 533574 452000 6 vdda2
port 535 nsew power input
rlabel metal4 s 32954 451308 33574 476000 6 vdda2
port 535 nsew power input
rlabel metal4 s 52954 451308 53574 476000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 451308 73574 476000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 451308 93574 476000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 451308 113574 476000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 451308 133574 476000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 451308 153574 476000 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 539308 253574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 539308 273574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 539308 293574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 539308 313574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 332954 539308 333574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 539308 413574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 539308 433574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 539308 453574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 539308 473574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 539308 493574 576000 6 vdda2
port 535 nsew power input
rlabel metal4 s 32954 563308 33574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 52954 563308 53574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 563308 73574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 563308 93574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 563308 113574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 563308 133574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 563308 153574 588000 6 vdda2
port 535 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 32954 675308 33574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 52954 675308 53574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 72954 675308 73574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 92954 675308 93574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 112954 675308 113574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 132954 675308 133574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 152954 675308 153574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 172954 -7654 173574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 212954 539308 213574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 232954 539308 233574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 252954 659500 253574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 272954 659500 273574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 292954 659500 293574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 312954 659500 313574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 332954 659500 333574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 352954 421162 353574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 421162 373574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 392954 421162 393574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 412954 659500 413574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 432954 659500 433574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 452954 659500 453574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 472954 659500 473574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 492954 659500 493574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 512954 539308 513574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 532954 539308 533574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 552954 421162 553574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 572954 -7654 573574 711590 6 vdda2
port 535 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 20306 590730 20926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 40306 590730 40926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 60306 590730 60926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 80306 590730 80926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 120306 590730 120926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 140306 590730 140926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 160306 590730 160926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 180306 590730 180926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 200306 590730 200926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 220306 590730 220926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 240306 590730 240926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 260306 590730 260926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 300306 590730 300926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 320306 590730 320926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 340306 590730 340926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 360306 590730 360926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 380306 590730 380926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 400306 590730 400926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 420306 590730 420926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 440306 590730 440926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 480306 590730 480926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 500306 590730 500926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 520306 590730 520926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 540306 590730 540926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 560306 590730 560926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 580306 590730 580926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 600306 590730 600926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 620306 590730 620926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 660306 590730 660926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 680306 590730 680926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 700306 590730 700926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 39234 -5734 39854 28000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 -5734 59854 28000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 -5734 79854 28000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 -5734 99854 28000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 -5734 119854 28000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 -5734 139854 28000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 -5734 159854 28000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 199234 -5734 199854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 -5734 219854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 -5734 239854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 -5734 259854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 -5734 299854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 -5734 319854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 339234 -5734 339854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 359234 -5734 359854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 379234 -5734 379854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 399234 -5734 399854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 419234 -5734 419854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439234 -5734 439854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 -5734 479854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 -5734 499854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 519234 -5734 519854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 539234 -5734 539854 58000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 39234 115308 39854 140000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 115308 59854 140000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 115308 79854 140000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 115308 99854 140000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 115308 119854 140000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 115308 139854 140000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 115308 159854 140000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 39234 227308 39854 252000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 227308 59854 252000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 227308 79854 252000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 227308 99854 252000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 227308 119854 252000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 227308 139854 252000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 227308 159854 252000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 39234 339308 39854 364000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 339308 59854 364000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 339308 79854 364000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 339308 99854 364000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 339308 119854 364000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 339308 139854 364000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 339308 159854 364000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 199234 421162 199854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 421162 219854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 421162 239854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 421162 259854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 421162 279854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 421162 299854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 421162 319854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 419234 421162 419854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439234 421162 439854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 421162 459854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 421162 479854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 421162 499854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 519234 421162 519854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 539234 421162 539854 452000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 39234 451308 39854 476000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 451308 59854 476000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 451308 79854 476000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 451308 99854 476000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 451308 119854 476000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 451308 139854 476000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 451308 159854 476000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 539308 239854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 539308 259854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 539308 279854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 539308 299854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 539308 319854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 419234 539308 419854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439234 539308 439854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 539308 459854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 539308 479854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 539308 499854 576000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 39234 563308 39854 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 563308 59854 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 563308 79854 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 563308 99854 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 563308 119854 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 563308 139854 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 563308 159854 588000 6 vssa1
port 536 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground input
rlabel metal4 s 19234 -5734 19854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 39234 675308 39854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 59234 675308 59854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 79234 675308 79854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 675308 99854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 119234 675308 119854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139234 675308 139854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 159234 675308 159854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 179234 -5734 179854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 199234 539308 199854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219234 539308 219854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239234 659500 239854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 259234 659500 259854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 659500 279854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 299234 659500 299854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 319234 659500 319854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 339234 421162 339854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 359234 421162 359854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 379234 421162 379854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 399234 421162 399854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 419234 659500 419854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 439234 659500 439854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 659500 459854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 479234 659500 479854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 499234 659500 499854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 519234 539308 519854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 539234 539308 539854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 559234 -5734 559854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 579234 -5734 579854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 24026 592650 24646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 44026 592650 44646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 64026 592650 64646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 84026 592650 84646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 124026 592650 124646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 144026 592650 144646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 164026 592650 164646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 184026 592650 184646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 204026 592650 204646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 224026 592650 224646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 244026 592650 244646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 264026 592650 264646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 304026 592650 304646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 324026 592650 324646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 344026 592650 344646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 364026 592650 364646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 384026 592650 384646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 404026 592650 404646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 424026 592650 424646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 444026 592650 444646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 484026 592650 484646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 504026 592650 504646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 524026 592650 524646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 544026 592650 544646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 564026 592650 564646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 584026 592650 584646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 604026 592650 604646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 624026 592650 624646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 664026 592650 664646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 684026 592650 684646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 42954 -7654 43574 28000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 -7654 63574 28000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 -7654 83574 28000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 -7654 103574 28000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 -7654 123574 28000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 -7654 143574 28000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 -7654 163574 28000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 202954 -7654 203574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 -7654 223574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 -7654 243574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 -7654 263574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 -7654 303574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 322954 -7654 323574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 342954 -7654 343574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 362954 -7654 363574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 382954 -7654 383574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 402954 -7654 403574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422954 -7654 423574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 442954 -7654 443574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 -7654 483574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 -7654 503574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 522954 -7654 523574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 542954 -7654 543574 58000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 42954 115308 43574 140000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 115308 63574 140000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 115308 83574 140000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 115308 103574 140000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 115308 123574 140000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 115308 143574 140000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 115308 163574 140000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 42954 227308 43574 252000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 227308 63574 252000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 227308 83574 252000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 227308 103574 252000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 227308 123574 252000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 227308 143574 252000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 227308 163574 252000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 42954 339308 43574 364000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 339308 63574 364000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 339308 83574 364000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 339308 103574 364000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 339308 123574 364000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 339308 143574 364000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 339308 163574 364000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 202954 421162 203574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 421162 223574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 421162 243574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 421162 263574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 421162 283574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 421162 303574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 322954 421162 323574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422954 421162 423574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 442954 421162 443574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 421162 463574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 421162 483574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 421162 503574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 522954 421162 523574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 542954 421162 543574 452000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 42954 451308 43574 476000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 451308 63574 476000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 451308 83574 476000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 451308 103574 476000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 451308 123574 476000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 451308 143574 476000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 451308 163574 476000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 539308 243574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 539308 263574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 539308 283574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 539308 303574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 322954 539308 323574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422954 539308 423574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 442954 539308 443574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 539308 463574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 539308 483574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 539308 503574 576000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 42954 563308 43574 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 563308 63574 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 563308 83574 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 563308 103574 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 563308 123574 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 563308 143574 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 563308 163574 588000 6 vssa2
port 537 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground input
rlabel metal4 s 22954 -7654 23574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 42954 675308 43574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 62954 675308 63574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 82954 675308 83574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 675308 103574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 122954 675308 123574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 142954 675308 143574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 162954 675308 163574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 182954 -7654 183574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 202954 539308 203574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222954 539308 223574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 242954 659500 243574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 262954 659500 263574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 659500 283574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 302954 659500 303574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 322954 659500 323574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 342954 421162 343574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 362954 421162 363574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 382954 421162 383574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 402954 421162 403574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 422954 659500 423574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 442954 659500 443574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 659500 463574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 482954 659500 483574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 502954 659500 503574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 522954 539308 523574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 542954 539308 543574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 562954 -7654 563574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 12866 586890 13486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 32866 586890 33486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 52866 586890 53486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 72866 586890 73486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 112866 586890 113486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 132866 586890 133486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 152866 586890 153486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 172866 586890 173486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 192866 586890 193486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 212866 586890 213486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 232866 586890 233486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 252866 586890 253486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 292866 586890 293486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 312866 586890 313486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 332866 586890 333486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 352866 586890 353486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 372866 586890 373486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 392866 586890 393486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 412866 586890 413486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 432866 586890 433486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 472866 586890 473486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 492866 586890 493486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 512866 586890 513486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 532866 586890 533486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 552866 586890 553486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 572866 586890 573486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 592866 586890 593486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 612866 586890 613486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 652866 586890 653486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 672866 586890 673486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 692866 586890 693486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 31794 -1894 32414 28000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 51794 -1894 52414 28000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 -1894 72414 28000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 -1894 92414 28000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 -1894 112414 28000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 -1894 132414 28000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 -1894 152414 28000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 211794 -1894 212414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 231794 -1894 232414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 -1894 252414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 -1894 292414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 -1894 312414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 331794 -1894 332414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 -1894 352414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 371794 -1894 372414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 391794 -1894 392414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 -1894 412414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 431794 -1894 432414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 -1894 472414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 -1894 492414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 511794 -1894 512414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 531794 -1894 532414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 551794 -1894 552414 58000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 31794 115308 32414 140000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 51794 115308 52414 140000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 115308 72414 140000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 115308 92414 140000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 115308 112414 140000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 115308 132414 140000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 115308 152414 140000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 31794 227308 32414 252000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 51794 227308 52414 252000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 227308 72414 252000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 227308 92414 252000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 227308 112414 252000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 227308 132414 252000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 227308 152414 252000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 31794 339308 32414 364000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 51794 339308 52414 364000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 339308 72414 364000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 339308 92414 364000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 339308 112414 364000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 339308 132414 364000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 339308 152414 364000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 211794 421162 212414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 231794 421162 232414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 421162 252414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 421162 272414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 421162 292414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 421162 312414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 331794 421162 332414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 421162 412414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 431794 421162 432414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 421162 452414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 421162 472414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 421162 492414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 511794 421162 512414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 531794 421162 532414 452000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 31794 451308 32414 476000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 51794 451308 52414 476000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 451308 72414 476000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 451308 92414 476000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 451308 112414 476000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 451308 132414 476000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 451308 152414 476000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 539308 252414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 539308 272414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 539308 292414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 539308 312414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 331794 539308 332414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 539308 412414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 431794 539308 432414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 539308 452414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 539308 472414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 539308 492414 576000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 31794 563308 32414 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 51794 563308 52414 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 563308 72414 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 563308 92414 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 563308 112414 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 563308 132414 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 563308 152414 588000 6 vssd1
port 538 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground input
rlabel metal4 s 11794 -1894 12414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 31794 675308 32414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 51794 675308 52414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 71794 675308 72414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 675308 92414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 111794 675308 112414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 131794 675308 132414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 151794 675308 152414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 171794 -1894 172414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 191794 -1894 192414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 211794 539308 212414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 231794 539308 232414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 251794 659500 252414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 659500 272414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 291794 659500 292414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 311794 659500 312414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 331794 659500 332414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 351794 421162 352414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 371794 421162 372414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 391794 421162 392414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 411794 659500 412414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 431794 659500 432414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 659500 452414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 471794 659500 472414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 491794 659500 492414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 511794 539308 512414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 531794 539308 532414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 551794 421162 552414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 571794 -1894 572414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 16586 588810 17206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 36586 588810 37206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 56586 588810 57206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 76586 588810 77206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 116586 588810 117206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 136586 588810 137206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 156586 588810 157206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 176586 588810 177206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 196586 588810 197206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 216586 588810 217206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 236586 588810 237206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 256586 588810 257206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 296586 588810 297206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 316586 588810 317206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 336586 588810 337206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 356586 588810 357206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 376586 588810 377206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 396586 588810 397206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 416586 588810 417206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 436586 588810 437206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 476586 588810 477206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 496586 588810 497206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 516586 588810 517206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 536586 588810 537206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 556586 588810 557206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 576586 588810 577206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 596586 588810 597206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 616586 588810 617206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 656586 588810 657206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 676586 588810 677206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 696586 588810 697206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 35514 -3814 36134 28000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 55514 -3814 56134 28000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 -3814 76134 28000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 -3814 96134 28000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 -3814 116134 28000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 -3814 136134 28000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 -3814 156134 28000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 215514 -3814 216134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235514 -3814 236134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 -3814 256134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 -3814 296134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 -3814 316134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 335514 -3814 336134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 -3814 356134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 375514 -3814 376134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 395514 -3814 396134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 -3814 416134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 435514 -3814 436134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 -3814 476134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 -3814 496134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 515514 -3814 516134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 535514 -3814 536134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 555514 -3814 556134 58000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 35514 115308 36134 140000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 55514 115308 56134 140000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 115308 76134 140000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 115308 96134 140000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 115308 116134 140000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 115308 136134 140000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 115308 156134 140000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 35514 227308 36134 252000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 55514 227308 56134 252000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 227308 76134 252000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 227308 96134 252000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 227308 116134 252000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 227308 136134 252000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 227308 156134 252000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 35514 339308 36134 364000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 55514 339308 56134 364000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 339308 76134 364000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 339308 96134 364000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 339308 116134 364000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 339308 136134 364000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 339308 156134 364000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 215514 421162 216134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235514 421162 236134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 421162 256134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 421162 276134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 421162 296134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 421162 316134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 335514 421162 336134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 421162 416134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 435514 421162 436134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 421162 456134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 421162 476134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 421162 496134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 515514 421162 516134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 535514 421162 536134 452000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 35514 451308 36134 476000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 55514 451308 56134 476000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 451308 76134 476000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 451308 96134 476000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 451308 116134 476000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 451308 136134 476000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 451308 156134 476000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 539308 256134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 539308 276134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 539308 296134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 539308 316134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 335514 539308 336134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 539308 416134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 435514 539308 436134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 539308 456134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 539308 476134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 539308 496134 576000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 35514 563308 36134 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 55514 563308 56134 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 563308 76134 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 563308 96134 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 563308 116134 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 563308 136134 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 563308 156134 588000 6 vssd2
port 539 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground input
rlabel metal4 s 15514 -3814 16134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 35514 675308 36134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 55514 675308 56134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 75514 675308 76134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 675308 96134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 115514 675308 116134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 135514 675308 136134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155514 675308 156134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 175514 -3814 176134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 195514 -3814 196134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 215514 539308 216134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235514 539308 236134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 255514 659500 256134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 659500 276134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 295514 659500 296134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 315514 659500 316134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 335514 659500 336134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 355514 421162 356134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 375514 421162 376134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 395514 421162 396134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 415514 659500 416134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 435514 659500 436134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 659500 456134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 475514 659500 476134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 495514 659500 496134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 515514 539308 516134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 535514 539308 536134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 555514 421162 556134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 575514 -3814 576134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29081168
string GDS_FILE /home/shc/Development/efabless/marmot_asic/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 25150374
<< end >>

