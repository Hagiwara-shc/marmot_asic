VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.330 2934.450 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 114.330 2934.450 117.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 214.330 2934.450 217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 314.330 2934.450 317.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 414.330 2934.450 417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 514.330 2934.450 517.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 614.330 2934.450 617.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 714.330 2934.450 717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 814.330 2934.450 817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 914.330 2934.450 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1014.330 2934.450 1017.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1114.330 2934.450 1117.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1214.330 2934.450 1217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1314.330 2934.450 1317.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1414.330 2934.450 1417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1514.330 2934.450 1517.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1614.330 2934.450 1617.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1714.330 2934.450 1717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1814.330 2934.450 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1914.330 2934.450 1917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2014.330 2934.450 2017.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2114.330 2934.450 2117.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2214.330 2934.450 2217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2314.330 2934.450 2317.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2414.330 2934.450 2417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2514.330 2934.450 2517.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2614.330 2934.450 2617.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2714.330 2934.450 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2814.330 2934.450 2817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2914.330 2934.450 2917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3014.330 2934.450 3017.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3114.330 2934.450 3117.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3214.330 2934.450 3217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3314.330 2934.450 3317.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3414.330 2934.450 3417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 -9.470 212.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 -9.470 312.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 -9.470 412.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.970 -9.470 512.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 -9.470 612.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 -9.470 712.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 -9.470 812.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.970 -9.470 1012.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1108.970 -9.470 1112.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.970 -9.470 1212.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1308.970 -9.470 1312.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 -9.470 1412.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1508.970 -9.470 1512.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.970 -9.470 1612.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1708.970 -9.470 1712.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -9.470 1812.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1908.970 -9.470 1912.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.970 -9.470 2012.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 -9.470 2112.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.970 -9.470 2212.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2308.970 -9.470 2312.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.970 -9.470 2412.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.970 -9.470 2512.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.970 -9.470 2612.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -9.470 2712.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 576.540 212.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 576.540 312.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 576.540 412.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.970 576.540 512.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 576.540 612.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 576.540 712.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 576.540 812.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 1136.540 212.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 1136.540 312.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 1136.540 412.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.970 1136.540 512.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 1136.540 612.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 1136.540 712.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 1136.540 812.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 1696.540 212.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 1696.540 312.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 1696.540 412.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.970 1696.540 512.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 1696.540 612.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 1696.540 712.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 1696.540 812.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.970 2077.100 1012.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1108.970 2077.100 1112.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.970 2077.100 1212.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1308.970 2077.100 1312.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 2077.100 1412.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1508.970 2077.100 1512.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.970 2077.100 1612.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 2077.100 2112.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.970 2077.100 2212.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2308.970 2077.100 2312.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.970 2077.100 2412.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.970 2077.100 2512.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.970 2077.100 2612.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 2077.100 2712.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 2256.540 212.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 2256.540 312.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 2256.540 412.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.970 2256.540 512.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 2256.540 612.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 2256.540 712.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 2256.540 812.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.970 2696.540 1212.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1308.970 2696.540 1312.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 2696.540 1412.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1508.970 2696.540 1512.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.970 2696.540 1612.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 2696.540 2112.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.970 2696.540 2212.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2308.970 2696.540 2312.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.970 2696.540 2412.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.970 2696.540 2512.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 2816.540 212.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 2816.540 312.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 2816.540 412.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.970 2816.540 512.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 2816.540 612.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 2816.540 712.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 2816.540 812.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.970 -9.470 112.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 3376.540 212.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 3376.540 312.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 3376.540 412.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.970 3376.540 512.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 3376.540 612.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 3376.540 712.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 3376.540 812.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -9.470 912.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.970 2696.540 1012.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1108.970 2696.540 1112.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.970 3297.500 1212.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1308.970 3297.500 1312.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 3297.500 1412.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1508.970 3297.500 1512.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.970 3297.500 1612.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1708.970 2077.100 1712.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 2077.100 1812.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1908.970 2077.100 1912.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.970 2077.100 2012.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.970 3297.500 2112.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.970 3297.500 2212.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2308.970 3297.500 2312.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.970 3297.500 2412.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.970 3297.500 2512.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.970 2696.540 2612.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 2696.540 2712.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.970 -9.470 2812.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2908.970 -9.470 2912.070 3529.150 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 32.930 2944.050 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 132.930 2944.050 136.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 232.930 2944.050 236.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 332.930 2944.050 336.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 432.930 2944.050 436.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 532.930 2944.050 536.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 632.930 2944.050 636.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 732.930 2944.050 736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 832.930 2944.050 836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 932.930 2944.050 936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1032.930 2944.050 1036.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1132.930 2944.050 1136.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1232.930 2944.050 1236.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1332.930 2944.050 1336.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1432.930 2944.050 1436.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1532.930 2944.050 1536.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1632.930 2944.050 1636.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1732.930 2944.050 1736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1832.930 2944.050 1836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1932.930 2944.050 1936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2032.930 2944.050 2036.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2132.930 2944.050 2136.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2232.930 2944.050 2236.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2332.930 2944.050 2336.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2432.930 2944.050 2436.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2532.930 2944.050 2536.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2632.930 2944.050 2636.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2732.930 2944.050 2736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2832.930 2944.050 2836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2932.930 2944.050 2936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3032.930 2944.050 3036.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3132.930 2944.050 3136.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3232.930 2944.050 3236.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3332.930 2944.050 3336.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3432.930 2944.050 3436.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 -19.070 230.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 -19.070 330.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 -19.070 430.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.570 -19.070 530.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.570 -19.070 630.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 -19.070 730.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 827.570 -19.070 830.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1027.570 -19.070 1030.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1127.570 -19.070 1130.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1227.570 -19.070 1230.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1327.570 -19.070 1330.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 -19.070 1430.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1527.570 -19.070 1530.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1627.570 -19.070 1630.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1727.570 -19.070 1730.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 -19.070 1830.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1927.570 -19.070 1930.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2027.570 -19.070 2030.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2127.570 -19.070 2130.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2227.570 -19.070 2230.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2327.570 -19.070 2330.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2427.570 -19.070 2430.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2527.570 -19.070 2530.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2627.570 -19.070 2630.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 -19.070 2730.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 576.540 230.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 576.540 330.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 576.540 430.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.570 576.540 530.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.570 576.540 630.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 576.540 730.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 827.570 576.540 830.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 1136.540 230.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 1136.540 330.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 1136.540 430.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.570 1136.540 530.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.570 1136.540 630.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 1136.540 730.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 827.570 1136.540 830.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 1696.540 230.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 1696.540 330.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 1696.540 430.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.570 1696.540 530.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.570 1696.540 630.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 1696.540 730.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 827.570 1696.540 830.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1027.570 2077.100 1030.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1127.570 2077.100 1130.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1227.570 2077.100 1230.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1327.570 2077.100 1330.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 2077.100 1430.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1527.570 2077.100 1530.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1627.570 2077.100 1630.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2127.570 2077.100 2130.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2227.570 2077.100 2230.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2327.570 2077.100 2330.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2427.570 2077.100 2430.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2527.570 2077.100 2530.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2627.570 2077.100 2630.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 2077.100 2730.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 2256.540 230.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 2256.540 330.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 2256.540 430.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.570 2256.540 530.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.570 2256.540 630.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 2256.540 730.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 827.570 2256.540 830.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1227.570 2696.540 1230.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1327.570 2696.540 1330.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 2696.540 1430.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1527.570 2696.540 1530.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1627.570 2696.540 1630.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2127.570 2696.540 2130.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2227.570 2696.540 2230.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2327.570 2696.540 2330.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2427.570 2696.540 2430.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2527.570 2696.540 2530.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 2816.540 230.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 2816.540 330.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 2816.540 430.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.570 2816.540 530.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.570 2816.540 630.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 2816.540 730.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 827.570 2816.540 830.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -19.070 30.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 127.570 -19.070 130.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 3376.540 230.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 3376.540 330.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 3376.540 430.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.570 3376.540 530.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.570 3376.540 630.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 3376.540 730.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 827.570 3376.540 830.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 -19.070 930.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1027.570 2696.540 1030.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1127.570 2696.540 1130.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1227.570 3297.500 1230.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1327.570 3297.500 1330.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1427.570 3297.500 1430.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1527.570 3297.500 1530.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1627.570 3297.500 1630.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1727.570 2077.100 1730.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 2077.100 1830.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1927.570 2077.100 1930.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2027.570 2077.100 2030.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2127.570 3297.500 2130.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2227.570 3297.500 2230.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2327.570 3297.500 2330.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2427.570 3297.500 2430.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2527.570 3297.500 2530.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2627.570 2696.540 2630.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 2696.540 2730.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2827.570 -19.070 2830.670 3538.750 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 51.530 2953.650 54.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 151.530 2953.650 154.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 251.530 2953.650 254.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 351.530 2953.650 354.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 451.530 2953.650 454.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 551.530 2953.650 554.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 651.530 2953.650 654.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 751.530 2953.650 754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 851.530 2953.650 854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 951.530 2953.650 954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1051.530 2953.650 1054.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1151.530 2953.650 1154.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1251.530 2953.650 1254.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1351.530 2953.650 1354.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1451.530 2953.650 1454.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1551.530 2953.650 1554.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1651.530 2953.650 1654.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1751.530 2953.650 1754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1851.530 2953.650 1854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1951.530 2953.650 1954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2051.530 2953.650 2054.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2151.530 2953.650 2154.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2251.530 2953.650 2254.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2351.530 2953.650 2354.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2451.530 2953.650 2454.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2551.530 2953.650 2554.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2651.530 2953.650 2654.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2751.530 2953.650 2754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2851.530 2953.650 2854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2951.530 2953.650 2954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3051.530 2953.650 3054.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3151.530 2953.650 3154.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3251.530 2953.650 3254.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3351.530 2953.650 3354.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3451.530 2953.650 3454.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.170 -28.670 149.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.170 -28.670 249.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.170 -28.670 349.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.170 -28.670 449.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.170 -28.670 549.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.170 -28.670 649.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 -28.670 749.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1046.170 -28.670 1049.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.170 -28.670 1149.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.170 -28.670 1249.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1346.170 -28.670 1349.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 -28.670 1449.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1546.170 -28.670 1549.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1646.170 -28.670 1649.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.170 -28.670 1749.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 -28.670 1849.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1946.170 -28.670 1949.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2046.170 -28.670 2049.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.170 -28.670 2149.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2246.170 -28.670 2249.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.170 -28.670 2349.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2446.170 -28.670 2449.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2546.170 -28.670 2549.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2646.170 -28.670 2649.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 -28.670 2749.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.170 576.540 149.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.170 576.540 249.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.170 576.540 349.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.170 576.540 449.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.170 576.540 549.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.170 576.540 649.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 576.540 749.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.170 1136.540 149.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.170 1136.540 249.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.170 1136.540 349.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.170 1136.540 449.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.170 1136.540 549.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.170 1136.540 649.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 1136.540 749.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.170 1696.540 149.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.170 1696.540 249.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.170 1696.540 349.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.170 1696.540 449.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.170 1696.540 549.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.170 1696.540 649.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 1696.540 749.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1046.170 2077.100 1049.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.170 2077.100 1149.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.170 2077.100 1249.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1346.170 2077.100 1349.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 2077.100 1449.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1546.170 2077.100 1549.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1646.170 2077.100 1649.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2046.170 2077.100 2049.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.170 2077.100 2149.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2246.170 2077.100 2249.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.170 2077.100 2349.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2446.170 2077.100 2449.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2546.170 2077.100 2549.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2646.170 2077.100 2649.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.170 2256.540 149.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.170 2256.540 249.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.170 2256.540 349.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.170 2256.540 449.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.170 2256.540 549.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.170 2256.540 649.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 2256.540 749.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.170 2696.540 1249.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1346.170 2696.540 1349.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 2696.540 1449.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1546.170 2696.540 1549.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1646.170 2696.540 1649.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2046.170 2696.540 2049.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.170 2696.540 2149.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2246.170 2696.540 2249.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.170 2696.540 2349.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2446.170 2696.540 2449.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.170 2816.540 149.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.170 2816.540 249.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.170 2816.540 349.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.170 2816.540 449.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.170 2816.540 549.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.170 2816.540 649.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 2816.540 749.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 -28.670 49.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.170 3376.540 149.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.170 3376.540 249.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.170 3376.540 349.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.170 3376.540 449.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.170 3376.540 549.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.170 3376.540 649.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.170 3376.540 749.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.170 -28.670 849.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 -28.670 949.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1046.170 2696.540 1049.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.170 2696.540 1149.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.170 3297.500 1249.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1346.170 3297.500 1349.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.170 3297.500 1449.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1546.170 3297.500 1549.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1646.170 3297.500 1649.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.170 2077.100 1749.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 2077.100 1849.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1946.170 2077.100 1949.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2046.170 3297.500 2049.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.170 3297.500 2149.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2246.170 3297.500 2249.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.170 3297.500 2349.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2446.170 3297.500 2449.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2546.170 2696.540 2549.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2646.170 2696.540 2649.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 2077.100 2749.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2846.170 -28.670 2849.270 3548.350 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 170.130 2963.250 173.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 270.130 2963.250 273.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 370.130 2963.250 373.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 470.130 2963.250 473.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 570.130 2963.250 573.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 670.130 2963.250 673.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 770.130 2963.250 773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 870.130 2963.250 873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 970.130 2963.250 973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1070.130 2963.250 1073.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1170.130 2963.250 1173.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1270.130 2963.250 1273.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1370.130 2963.250 1373.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1470.130 2963.250 1473.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1570.130 2963.250 1573.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1670.130 2963.250 1673.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1770.130 2963.250 1773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1970.130 2963.250 1973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2070.130 2963.250 2073.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2170.130 2963.250 2173.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2270.130 2963.250 2273.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2370.130 2963.250 2373.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2470.130 2963.250 2473.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2570.130 2963.250 2573.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2670.130 2963.250 2673.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2870.130 2963.250 2873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2970.130 2963.250 2973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3070.130 2963.250 3073.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3170.130 2963.250 3173.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3270.130 2963.250 3273.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3370.130 2963.250 3373.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3470.130 2963.250 3473.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.770 -38.270 167.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.770 -38.270 267.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.770 -38.270 367.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.770 -38.270 467.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.770 -38.270 567.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.770 -38.270 667.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 -38.270 767.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1064.770 -38.270 1067.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.770 -38.270 1167.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1264.770 -38.270 1267.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1364.770 -38.270 1367.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 -38.270 1467.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1564.770 -38.270 1567.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1664.770 -38.270 1667.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1764.770 -38.270 1767.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 -38.270 1867.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1964.770 -38.270 1967.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2064.770 -38.270 2067.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.770 -38.270 2167.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2264.770 -38.270 2267.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2364.770 -38.270 2367.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2464.770 -38.270 2467.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2564.770 -38.270 2567.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2664.770 -38.270 2667.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 -38.270 2767.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.770 576.540 167.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.770 576.540 267.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.770 576.540 367.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.770 576.540 467.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.770 576.540 567.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.770 576.540 667.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 576.540 767.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.770 1136.540 167.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.770 1136.540 267.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.770 1136.540 367.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.770 1136.540 467.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.770 1136.540 567.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.770 1136.540 667.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 1136.540 767.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.770 1696.540 167.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.770 1696.540 267.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.770 1696.540 367.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.770 1696.540 467.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.770 1696.540 567.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.770 1696.540 667.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 1696.540 767.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1064.770 2077.100 1067.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.770 2077.100 1167.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1264.770 2077.100 1267.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1364.770 2077.100 1367.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 2077.100 1467.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1564.770 2077.100 1567.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1664.770 2077.100 1667.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2064.770 2077.100 2067.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.770 2077.100 2167.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2264.770 2077.100 2267.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2364.770 2077.100 2367.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2464.770 2077.100 2467.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2564.770 2077.100 2567.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2664.770 2077.100 2667.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.770 2256.540 167.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.770 2256.540 267.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.770 2256.540 367.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.770 2256.540 467.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.770 2256.540 567.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.770 2256.540 667.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 2256.540 767.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1264.770 2696.540 1267.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1364.770 2696.540 1367.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 2696.540 1467.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1564.770 2696.540 1567.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1664.770 2696.540 1667.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2064.770 2696.540 2067.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.770 2696.540 2167.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2264.770 2696.540 2267.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2364.770 2696.540 2367.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2464.770 2696.540 2467.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.770 2816.540 167.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.770 2816.540 267.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.770 2816.540 367.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.770 2816.540 467.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.770 2816.540 567.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.770 2816.540 667.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 2816.540 767.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.770 3376.540 167.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.770 3376.540 267.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.770 3376.540 367.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.770 3376.540 467.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.770 3376.540 567.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.770 3376.540 667.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 764.770 3376.540 767.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.770 -38.270 867.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 -38.270 967.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1064.770 2696.540 1067.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.770 2696.540 1167.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1264.770 3297.500 1267.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1364.770 3297.500 1367.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.770 3297.500 1467.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1564.770 3297.500 1567.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1664.770 3297.500 1667.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1764.770 2077.100 1767.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 2077.100 1867.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1964.770 2077.100 1967.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2064.770 3297.500 2067.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2164.770 3297.500 2167.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2264.770 3297.500 2267.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2364.770 3297.500 2367.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2464.770 3297.500 2467.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2564.770 2696.540 2567.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2664.770 2696.540 2667.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 2077.100 2767.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2864.770 -38.270 2867.870 3557.950 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 101.530 2953.650 104.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 201.530 2953.650 204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 301.530 2953.650 304.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 401.530 2953.650 404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 501.530 2953.650 504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 601.530 2953.650 604.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 701.530 2953.650 704.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 801.530 2953.650 804.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 901.530 2953.650 904.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1001.530 2953.650 1004.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1101.530 2953.650 1104.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1201.530 2953.650 1204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1301.530 2953.650 1304.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1401.530 2953.650 1404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1501.530 2953.650 1504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1601.530 2953.650 1604.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1701.530 2953.650 1704.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1801.530 2953.650 1804.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1901.530 2953.650 1904.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2001.530 2953.650 2004.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2101.530 2953.650 2104.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2201.530 2953.650 2204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2301.530 2953.650 2304.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2401.530 2953.650 2404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2501.530 2953.650 2504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2601.530 2953.650 2604.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2701.530 2953.650 2704.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2801.530 2953.650 2804.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2901.530 2953.650 2904.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3001.530 2953.650 3004.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3101.530 2953.650 3104.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3301.530 2953.650 3304.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3401.530 2953.650 3404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3501.530 2953.650 3504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.170 -28.670 199.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.170 -28.670 299.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 -28.670 399.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 -28.670 499.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.170 -28.670 599.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.170 -28.670 699.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.170 -28.670 799.270 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.170 -28.670 999.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.170 -28.670 1099.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1196.170 -28.670 1199.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1296.170 -28.670 1299.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 -28.670 1399.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.170 -28.670 1499.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1596.170 -28.670 1599.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1696.170 -28.670 1699.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1796.170 -28.670 1799.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1896.170 -28.670 1899.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1996.170 -28.670 1999.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2096.170 -28.670 2099.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2196.170 -28.670 2199.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 -28.670 2299.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2396.170 -28.670 2399.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 -28.670 2499.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2596.170 -28.670 2599.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2696.170 -28.670 2699.270 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.170 576.540 199.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.170 576.540 299.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 576.540 399.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 576.540 499.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.170 576.540 599.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.170 576.540 699.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.170 576.540 799.270 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.170 1136.540 199.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.170 1136.540 299.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 1136.540 399.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 1136.540 499.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.170 1136.540 599.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.170 1136.540 699.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.170 1136.540 799.270 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.170 1696.540 199.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.170 1696.540 299.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 1696.540 399.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 1696.540 499.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.170 1696.540 599.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.170 1696.540 699.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.170 1696.540 799.270 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.170 2077.100 999.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.170 2077.100 1099.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1196.170 2077.100 1199.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1296.170 2077.100 1299.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 2077.100 1399.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.170 2077.100 1499.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1596.170 2077.100 1599.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2096.170 2077.100 2099.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2196.170 2077.100 2199.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 2077.100 2299.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2396.170 2077.100 2399.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 2077.100 2499.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2596.170 2077.100 2599.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2696.170 2077.100 2699.270 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.170 2256.540 199.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.170 2256.540 299.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 2256.540 399.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 2256.540 499.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.170 2256.540 599.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.170 2256.540 699.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.170 2256.540 799.270 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1196.170 2696.540 1199.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1296.170 2696.540 1299.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 2696.540 1399.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.170 2696.540 1499.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1596.170 2696.540 1599.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2096.170 2696.540 2099.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2196.170 2696.540 2199.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 2696.540 2299.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2396.170 2696.540 2399.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 2696.540 2499.270 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.170 2816.540 199.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.170 2816.540 299.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 2816.540 399.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 2816.540 499.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.170 2816.540 599.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.170 2816.540 699.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.170 2816.540 799.270 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.170 -28.670 99.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.170 3376.540 199.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.170 3376.540 299.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.170 3376.540 399.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 3376.540 499.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.170 3376.540 599.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.170 3376.540 699.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.170 3376.540 799.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 896.170 -28.670 899.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.170 2696.540 999.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.170 2696.540 1099.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1196.170 3297.500 1199.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1296.170 3297.500 1299.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 3297.500 1399.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.170 3297.500 1499.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1596.170 3297.500 1599.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1696.170 2077.100 1699.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1796.170 2077.100 1799.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1896.170 2077.100 1899.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1996.170 2077.100 1999.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2096.170 3297.500 2099.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2196.170 3297.500 2199.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 3297.500 2299.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2396.170 3297.500 2399.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.170 3297.500 2499.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2596.170 2696.540 2599.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2696.170 2696.540 2699.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2796.170 -28.670 2799.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2896.170 -28.670 2899.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 120.130 2963.250 123.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 220.130 2963.250 223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 320.130 2963.250 323.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 420.130 2963.250 423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 520.130 2963.250 523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 620.130 2963.250 623.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 720.130 2963.250 723.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 820.130 2963.250 823.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 920.130 2963.250 923.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1020.130 2963.250 1023.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1120.130 2963.250 1123.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1220.130 2963.250 1223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1320.130 2963.250 1323.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1420.130 2963.250 1423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1520.130 2963.250 1523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1620.130 2963.250 1623.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1720.130 2963.250 1723.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1820.130 2963.250 1823.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1920.130 2963.250 1923.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2020.130 2963.250 2023.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2120.130 2963.250 2123.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2220.130 2963.250 2223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2320.130 2963.250 2323.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2420.130 2963.250 2423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2520.130 2963.250 2523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2620.130 2963.250 2623.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2720.130 2963.250 2723.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2820.130 2963.250 2823.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2920.130 2963.250 2923.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3020.130 2963.250 3023.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3120.130 2963.250 3123.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3320.130 2963.250 3323.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3420.130 2963.250 3423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.770 -38.270 217.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.770 -38.270 317.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 -38.270 417.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 -38.270 517.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.770 -38.270 617.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 714.770 -38.270 717.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.770 -38.270 817.870 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1014.770 -38.270 1017.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.770 -38.270 1117.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1214.770 -38.270 1217.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1314.770 -38.270 1317.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 -38.270 1417.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1514.770 -38.270 1517.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.770 -38.270 1617.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1714.770 -38.270 1717.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1814.770 -38.270 1817.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1914.770 -38.270 1917.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2014.770 -38.270 2017.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.770 -38.270 2117.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.770 -38.270 2217.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 -38.270 2317.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2414.770 -38.270 2417.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 -38.270 2517.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2614.770 -38.270 2617.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2714.770 -38.270 2717.870 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.770 576.540 217.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.770 576.540 317.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 576.540 417.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 576.540 517.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.770 576.540 617.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 714.770 576.540 717.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.770 576.540 817.870 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.770 1136.540 217.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.770 1136.540 317.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 1136.540 417.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 1136.540 517.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.770 1136.540 617.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 714.770 1136.540 717.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.770 1136.540 817.870 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.770 1696.540 217.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.770 1696.540 317.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 1696.540 417.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 1696.540 517.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.770 1696.540 617.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 714.770 1696.540 717.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.770 1696.540 817.870 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1014.770 2077.100 1017.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.770 2077.100 1117.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1214.770 2077.100 1217.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1314.770 2077.100 1317.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 2077.100 1417.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1514.770 2077.100 1517.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.770 2077.100 1617.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.770 2077.100 2117.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.770 2077.100 2217.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 2077.100 2317.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2414.770 2077.100 2417.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 2077.100 2517.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2614.770 2077.100 2617.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2714.770 2077.100 2717.870 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.770 2256.540 217.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.770 2256.540 317.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 2256.540 417.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 2256.540 517.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.770 2256.540 617.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 714.770 2256.540 717.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.770 2256.540 817.870 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1214.770 2696.540 1217.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1314.770 2696.540 1317.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 2696.540 1417.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1514.770 2696.540 1517.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.770 2696.540 1617.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.770 2696.540 2117.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.770 2696.540 2217.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 2696.540 2317.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2414.770 2696.540 2417.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 2696.540 2517.870 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.770 2816.540 217.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.770 2816.540 317.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 2816.540 417.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 2816.540 517.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.770 2816.540 617.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 714.770 2816.540 717.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.770 2816.540 817.870 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.770 -38.270 117.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.770 3376.540 217.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.770 3376.540 317.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.770 3376.540 417.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 3376.540 517.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.770 3376.540 617.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 714.770 3376.540 717.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.770 3376.540 817.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 914.770 -38.270 917.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1014.770 2696.540 1017.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.770 2696.540 1117.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1214.770 3297.500 1217.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1314.770 3297.500 1317.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 3297.500 1417.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1514.770 3297.500 1517.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.770 3297.500 1617.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1714.770 2077.100 1717.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1814.770 2077.100 1817.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1914.770 2077.100 1917.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2014.770 2077.100 2017.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.770 3297.500 2117.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.770 3297.500 2217.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 3297.500 2317.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2414.770 3297.500 2417.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2514.770 3297.500 2517.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2614.770 2696.540 2617.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2714.770 2696.540 2717.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2814.770 -38.270 2817.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 64.330 2934.450 67.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 164.330 2934.450 167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 264.330 2934.450 267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 364.330 2934.450 367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 464.330 2934.450 467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 564.330 2934.450 567.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 664.330 2934.450 667.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 764.330 2934.450 767.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 864.330 2934.450 867.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 964.330 2934.450 967.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1064.330 2934.450 1067.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1164.330 2934.450 1167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1264.330 2934.450 1267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1364.330 2934.450 1367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1464.330 2934.450 1467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1564.330 2934.450 1567.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1664.330 2934.450 1667.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1764.330 2934.450 1767.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1864.330 2934.450 1867.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1964.330 2934.450 1967.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2064.330 2934.450 2067.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2164.330 2934.450 2167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2264.330 2934.450 2267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2364.330 2934.450 2367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2464.330 2934.450 2467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2564.330 2934.450 2567.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2664.330 2934.450 2667.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2764.330 2934.450 2767.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2864.330 2934.450 2867.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2964.330 2934.450 2967.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3064.330 2934.450 3067.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3164.330 2934.450 3167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3264.330 2934.450 3267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3364.330 2934.450 3367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3464.330 2934.450 3467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.970 -9.470 162.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.970 -9.470 262.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 -9.470 362.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 -9.470 462.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.970 -9.470 562.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.970 -9.470 662.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.970 -9.470 762.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.970 -9.470 1062.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1158.970 -9.470 1162.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.970 -9.470 1262.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 -9.470 1362.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1458.970 -9.470 1462.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1558.970 -9.470 1562.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.970 -9.470 1662.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.970 -9.470 1762.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1858.970 -9.470 1862.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 -9.470 1962.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2058.970 -9.470 2062.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2158.970 -9.470 2162.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 -9.470 2262.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2358.970 -9.470 2362.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 -9.470 2462.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.970 -9.470 2562.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.970 -9.470 2662.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.970 -9.470 2762.070 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.970 576.540 162.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.970 576.540 262.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 576.540 362.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 576.540 462.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.970 576.540 562.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.970 576.540 662.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.970 576.540 762.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.970 1136.540 162.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.970 1136.540 262.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 1136.540 362.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1136.540 462.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.970 1136.540 562.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.970 1136.540 662.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.970 1136.540 762.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.970 1696.540 162.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.970 1696.540 262.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 1696.540 362.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1696.540 462.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.970 1696.540 562.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.970 1696.540 662.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.970 1696.540 762.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.970 2077.100 1062.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1158.970 2077.100 1162.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.970 2077.100 1262.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 2077.100 1362.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1458.970 2077.100 1462.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1558.970 2077.100 1562.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.970 2077.100 1662.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2058.970 2077.100 2062.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2158.970 2077.100 2162.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2077.100 2262.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2358.970 2077.100 2362.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 2077.100 2462.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.970 2077.100 2562.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.970 2077.100 2662.070 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.970 2256.540 162.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.970 2256.540 262.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 2256.540 362.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2256.540 462.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.970 2256.540 562.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.970 2256.540 662.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.970 2256.540 762.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.970 2696.540 1262.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 2696.540 1362.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1458.970 2696.540 1462.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1558.970 2696.540 1562.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.970 2696.540 1662.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2058.970 2696.540 2062.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2158.970 2696.540 2162.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2696.540 2262.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2358.970 2696.540 2362.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 2696.540 2462.070 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.970 2816.540 162.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.970 2816.540 262.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 2816.540 362.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2816.540 462.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.970 2816.540 562.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.970 2816.540 662.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.970 2816.540 762.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.970 -9.470 62.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.970 3376.540 162.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.970 3376.540 262.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.970 3376.540 362.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 3376.540 462.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.970 3376.540 562.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.970 3376.540 662.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.970 3376.540 762.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.970 -9.470 862.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 958.970 -9.470 962.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.970 2696.540 1062.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1158.970 2696.540 1162.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.970 3297.500 1262.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 3297.500 1362.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1458.970 3297.500 1462.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1558.970 3297.500 1562.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.970 3297.500 1662.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.970 2077.100 1762.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1858.970 2077.100 1862.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 2077.100 1962.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2058.970 3297.500 2062.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2158.970 3297.500 2162.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 3297.500 2262.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2358.970 3297.500 2362.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.970 3297.500 2462.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.970 2696.540 2562.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.970 2696.540 2662.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.970 2077.100 2762.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2858.970 -9.470 2862.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 82.930 2944.050 86.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 182.930 2944.050 186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 282.930 2944.050 286.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 382.930 2944.050 386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 482.930 2944.050 486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 582.930 2944.050 586.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 682.930 2944.050 686.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 782.930 2944.050 786.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 882.930 2944.050 886.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 982.930 2944.050 986.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1082.930 2944.050 1086.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1182.930 2944.050 1186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1282.930 2944.050 1286.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1382.930 2944.050 1386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1482.930 2944.050 1486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1582.930 2944.050 1586.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1682.930 2944.050 1686.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1782.930 2944.050 1786.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1882.930 2944.050 1886.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1982.930 2944.050 1986.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2082.930 2944.050 2086.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2182.930 2944.050 2186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2282.930 2944.050 2286.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2382.930 2944.050 2386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2482.930 2944.050 2486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2582.930 2944.050 2586.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2682.930 2944.050 2686.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2782.930 2944.050 2786.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2882.930 2944.050 2886.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2982.930 2944.050 2986.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3082.930 2944.050 3086.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3282.930 2944.050 3286.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3382.930 2944.050 3386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3482.930 2944.050 3486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.570 -19.070 180.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 277.570 -19.070 280.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 -19.070 380.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 -19.070 480.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 577.570 -19.070 580.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 677.570 -19.070 680.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.570 -19.070 780.670 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1077.570 -19.070 1080.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1177.570 -19.070 1180.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1277.570 -19.070 1280.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 -19.070 1380.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1477.570 -19.070 1480.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1577.570 -19.070 1580.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1677.570 -19.070 1680.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1777.570 -19.070 1780.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1877.570 -19.070 1880.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1977.570 -19.070 1980.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2077.570 -19.070 2080.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.570 -19.070 2180.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 -19.070 2280.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2377.570 -19.070 2380.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 -19.070 2480.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2577.570 -19.070 2580.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2677.570 -19.070 2680.670 290.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.570 576.540 180.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 277.570 576.540 280.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 576.540 380.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 576.540 480.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 577.570 576.540 580.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 677.570 576.540 680.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.570 576.540 780.670 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.570 1136.540 180.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 277.570 1136.540 280.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 1136.540 380.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 1136.540 480.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 577.570 1136.540 580.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 677.570 1136.540 680.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.570 1136.540 780.670 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.570 1696.540 180.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 277.570 1696.540 280.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 1696.540 380.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 1696.540 480.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 577.570 1696.540 580.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 677.570 1696.540 680.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.570 1696.540 780.670 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1077.570 2077.100 1080.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1177.570 2077.100 1180.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1277.570 2077.100 1280.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 2077.100 1380.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1477.570 2077.100 1480.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1577.570 2077.100 1580.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1677.570 2077.100 1680.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2077.570 2077.100 2080.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.570 2077.100 2180.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 2077.100 2280.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2377.570 2077.100 2380.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 2077.100 2480.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2577.570 2077.100 2580.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2677.570 2077.100 2680.670 2260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.570 2256.540 180.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 277.570 2256.540 280.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 2256.540 380.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 2256.540 480.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 577.570 2256.540 580.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 677.570 2256.540 680.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.570 2256.540 780.670 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1277.570 2696.540 1280.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 2696.540 1380.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1477.570 2696.540 1480.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1577.570 2696.540 1580.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1677.570 2696.540 1680.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2077.570 2696.540 2080.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.570 2696.540 2180.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 2696.540 2280.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2377.570 2696.540 2380.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 2696.540 2480.670 2880.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.570 2816.540 180.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 277.570 2816.540 280.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 2816.540 380.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 2816.540 480.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 577.570 2816.540 580.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 677.570 2816.540 680.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.570 2816.540 780.670 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 77.570 -19.070 80.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.570 3376.540 180.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 277.570 3376.540 280.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 377.570 3376.540 380.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 3376.540 480.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 577.570 3376.540 580.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 677.570 3376.540 680.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.570 3376.540 780.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 877.570 -19.070 880.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 977.570 -19.070 980.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1077.570 2696.540 1080.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1177.570 2696.540 1180.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1277.570 3297.500 1280.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 3297.500 1380.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1477.570 3297.500 1480.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1577.570 3297.500 1580.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1677.570 3297.500 1680.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1777.570 2077.100 1780.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1877.570 2077.100 1880.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1977.570 2077.100 1980.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2077.570 3297.500 2080.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.570 3297.500 2180.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 3297.500 2280.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2377.570 3297.500 2380.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2477.570 3297.500 2480.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2577.570 2696.540 2580.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2677.570 2696.540 2680.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2777.570 -19.070 2780.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2877.570 -19.070 2880.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 1005.520 310.795 2750.760 2054.485 ;
      LAYER met1 ;
        RECT 2.830 13.980 2912.190 3503.660 ;
      LAYER met2 ;
        RECT 2.860 3517.320 40.150 3518.050 ;
        RECT 41.270 3517.320 121.110 3518.050 ;
        RECT 122.230 3517.320 202.070 3518.050 ;
        RECT 203.190 3517.320 283.490 3518.050 ;
        RECT 284.610 3517.320 364.450 3518.050 ;
        RECT 365.570 3517.320 445.410 3518.050 ;
        RECT 446.530 3517.320 526.830 3518.050 ;
        RECT 527.950 3517.320 607.790 3518.050 ;
        RECT 608.910 3517.320 688.750 3518.050 ;
        RECT 689.870 3517.320 770.170 3518.050 ;
        RECT 771.290 3517.320 851.130 3518.050 ;
        RECT 852.250 3517.320 932.090 3518.050 ;
        RECT 933.210 3517.320 1013.510 3518.050 ;
        RECT 1014.630 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1175.430 3518.050 ;
        RECT 1176.550 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1500.190 3518.050 ;
        RECT 1501.310 3517.320 1581.150 3518.050 ;
        RECT 1582.270 3517.320 1662.110 3518.050 ;
        RECT 1663.230 3517.320 1743.530 3518.050 ;
        RECT 1744.650 3517.320 1824.490 3518.050 ;
        RECT 1825.610 3517.320 1905.450 3518.050 ;
        RECT 1906.570 3517.320 1986.870 3518.050 ;
        RECT 1987.990 3517.320 2067.830 3518.050 ;
        RECT 2068.950 3517.320 2148.790 3518.050 ;
        RECT 2149.910 3517.320 2230.210 3518.050 ;
        RECT 2231.330 3517.320 2311.170 3518.050 ;
        RECT 2312.290 3517.320 2392.130 3518.050 ;
        RECT 2393.250 3517.320 2473.550 3518.050 ;
        RECT 2474.670 3517.320 2554.510 3518.050 ;
        RECT 2555.630 3517.320 2635.470 3518.050 ;
        RECT 2636.590 3517.320 2716.890 3518.050 ;
        RECT 2718.010 3517.320 2797.850 3518.050 ;
        RECT 2798.970 3517.320 2878.810 3518.050 ;
        RECT 2879.930 3517.320 2917.160 3518.050 ;
        RECT 2.860 2.680 2917.160 3517.320 ;
        RECT 3.550 1.630 7.950 2.680 ;
        RECT 9.070 1.630 13.930 2.680 ;
        RECT 15.050 1.630 19.910 2.680 ;
        RECT 21.030 1.630 25.890 2.680 ;
        RECT 27.010 1.630 31.870 2.680 ;
        RECT 32.990 1.630 37.850 2.680 ;
        RECT 38.970 1.630 43.370 2.680 ;
        RECT 44.490 1.630 49.350 2.680 ;
        RECT 50.470 1.630 55.330 2.680 ;
        RECT 56.450 1.630 61.310 2.680 ;
        RECT 62.430 1.630 67.290 2.680 ;
        RECT 68.410 1.630 73.270 2.680 ;
        RECT 74.390 1.630 79.250 2.680 ;
        RECT 80.370 1.630 84.770 2.680 ;
        RECT 85.890 1.630 90.750 2.680 ;
        RECT 91.870 1.630 96.730 2.680 ;
        RECT 97.850 1.630 102.710 2.680 ;
        RECT 103.830 1.630 108.690 2.680 ;
        RECT 109.810 1.630 114.670 2.680 ;
        RECT 115.790 1.630 120.650 2.680 ;
        RECT 121.770 1.630 126.170 2.680 ;
        RECT 127.290 1.630 132.150 2.680 ;
        RECT 133.270 1.630 138.130 2.680 ;
        RECT 139.250 1.630 144.110 2.680 ;
        RECT 145.230 1.630 150.090 2.680 ;
        RECT 151.210 1.630 156.070 2.680 ;
        RECT 157.190 1.630 161.590 2.680 ;
        RECT 162.710 1.630 167.570 2.680 ;
        RECT 168.690 1.630 173.550 2.680 ;
        RECT 174.670 1.630 179.530 2.680 ;
        RECT 180.650 1.630 185.510 2.680 ;
        RECT 186.630 1.630 191.490 2.680 ;
        RECT 192.610 1.630 197.470 2.680 ;
        RECT 198.590 1.630 202.990 2.680 ;
        RECT 204.110 1.630 208.970 2.680 ;
        RECT 210.090 1.630 214.950 2.680 ;
        RECT 216.070 1.630 220.930 2.680 ;
        RECT 222.050 1.630 226.910 2.680 ;
        RECT 228.030 1.630 232.890 2.680 ;
        RECT 234.010 1.630 238.870 2.680 ;
        RECT 239.990 1.630 244.390 2.680 ;
        RECT 245.510 1.630 250.370 2.680 ;
        RECT 251.490 1.630 256.350 2.680 ;
        RECT 257.470 1.630 262.330 2.680 ;
        RECT 263.450 1.630 268.310 2.680 ;
        RECT 269.430 1.630 274.290 2.680 ;
        RECT 275.410 1.630 279.810 2.680 ;
        RECT 280.930 1.630 285.790 2.680 ;
        RECT 286.910 1.630 291.770 2.680 ;
        RECT 292.890 1.630 297.750 2.680 ;
        RECT 298.870 1.630 303.730 2.680 ;
        RECT 304.850 1.630 309.710 2.680 ;
        RECT 310.830 1.630 315.690 2.680 ;
        RECT 316.810 1.630 321.210 2.680 ;
        RECT 322.330 1.630 327.190 2.680 ;
        RECT 328.310 1.630 333.170 2.680 ;
        RECT 334.290 1.630 339.150 2.680 ;
        RECT 340.270 1.630 345.130 2.680 ;
        RECT 346.250 1.630 351.110 2.680 ;
        RECT 352.230 1.630 357.090 2.680 ;
        RECT 358.210 1.630 362.610 2.680 ;
        RECT 363.730 1.630 368.590 2.680 ;
        RECT 369.710 1.630 374.570 2.680 ;
        RECT 375.690 1.630 380.550 2.680 ;
        RECT 381.670 1.630 386.530 2.680 ;
        RECT 387.650 1.630 392.510 2.680 ;
        RECT 393.630 1.630 398.030 2.680 ;
        RECT 399.150 1.630 404.010 2.680 ;
        RECT 405.130 1.630 409.990 2.680 ;
        RECT 411.110 1.630 415.970 2.680 ;
        RECT 417.090 1.630 421.950 2.680 ;
        RECT 423.070 1.630 427.930 2.680 ;
        RECT 429.050 1.630 433.910 2.680 ;
        RECT 435.030 1.630 439.430 2.680 ;
        RECT 440.550 1.630 445.410 2.680 ;
        RECT 446.530 1.630 451.390 2.680 ;
        RECT 452.510 1.630 457.370 2.680 ;
        RECT 458.490 1.630 463.350 2.680 ;
        RECT 464.470 1.630 469.330 2.680 ;
        RECT 470.450 1.630 475.310 2.680 ;
        RECT 476.430 1.630 480.830 2.680 ;
        RECT 481.950 1.630 486.810 2.680 ;
        RECT 487.930 1.630 492.790 2.680 ;
        RECT 493.910 1.630 498.770 2.680 ;
        RECT 499.890 1.630 504.750 2.680 ;
        RECT 505.870 1.630 510.730 2.680 ;
        RECT 511.850 1.630 516.250 2.680 ;
        RECT 517.370 1.630 522.230 2.680 ;
        RECT 523.350 1.630 528.210 2.680 ;
        RECT 529.330 1.630 534.190 2.680 ;
        RECT 535.310 1.630 540.170 2.680 ;
        RECT 541.290 1.630 546.150 2.680 ;
        RECT 547.270 1.630 552.130 2.680 ;
        RECT 553.250 1.630 557.650 2.680 ;
        RECT 558.770 1.630 563.630 2.680 ;
        RECT 564.750 1.630 569.610 2.680 ;
        RECT 570.730 1.630 575.590 2.680 ;
        RECT 576.710 1.630 581.570 2.680 ;
        RECT 582.690 1.630 587.550 2.680 ;
        RECT 588.670 1.630 593.530 2.680 ;
        RECT 594.650 1.630 599.050 2.680 ;
        RECT 600.170 1.630 605.030 2.680 ;
        RECT 606.150 1.630 611.010 2.680 ;
        RECT 612.130 1.630 616.990 2.680 ;
        RECT 618.110 1.630 622.970 2.680 ;
        RECT 624.090 1.630 628.950 2.680 ;
        RECT 630.070 1.630 634.470 2.680 ;
        RECT 635.590 1.630 640.450 2.680 ;
        RECT 641.570 1.630 646.430 2.680 ;
        RECT 647.550 1.630 652.410 2.680 ;
        RECT 653.530 1.630 658.390 2.680 ;
        RECT 659.510 1.630 664.370 2.680 ;
        RECT 665.490 1.630 670.350 2.680 ;
        RECT 671.470 1.630 675.870 2.680 ;
        RECT 676.990 1.630 681.850 2.680 ;
        RECT 682.970 1.630 687.830 2.680 ;
        RECT 688.950 1.630 693.810 2.680 ;
        RECT 694.930 1.630 699.790 2.680 ;
        RECT 700.910 1.630 705.770 2.680 ;
        RECT 706.890 1.630 711.750 2.680 ;
        RECT 712.870 1.630 717.270 2.680 ;
        RECT 718.390 1.630 723.250 2.680 ;
        RECT 724.370 1.630 729.230 2.680 ;
        RECT 730.350 1.630 735.210 2.680 ;
        RECT 736.330 1.630 741.190 2.680 ;
        RECT 742.310 1.630 747.170 2.680 ;
        RECT 748.290 1.630 752.690 2.680 ;
        RECT 753.810 1.630 758.670 2.680 ;
        RECT 759.790 1.630 764.650 2.680 ;
        RECT 765.770 1.630 770.630 2.680 ;
        RECT 771.750 1.630 776.610 2.680 ;
        RECT 777.730 1.630 782.590 2.680 ;
        RECT 783.710 1.630 788.570 2.680 ;
        RECT 789.690 1.630 794.090 2.680 ;
        RECT 795.210 1.630 800.070 2.680 ;
        RECT 801.190 1.630 806.050 2.680 ;
        RECT 807.170 1.630 812.030 2.680 ;
        RECT 813.150 1.630 818.010 2.680 ;
        RECT 819.130 1.630 823.990 2.680 ;
        RECT 825.110 1.630 829.970 2.680 ;
        RECT 831.090 1.630 835.490 2.680 ;
        RECT 836.610 1.630 841.470 2.680 ;
        RECT 842.590 1.630 847.450 2.680 ;
        RECT 848.570 1.630 853.430 2.680 ;
        RECT 854.550 1.630 859.410 2.680 ;
        RECT 860.530 1.630 865.390 2.680 ;
        RECT 866.510 1.630 870.910 2.680 ;
        RECT 872.030 1.630 876.890 2.680 ;
        RECT 878.010 1.630 882.870 2.680 ;
        RECT 883.990 1.630 888.850 2.680 ;
        RECT 889.970 1.630 894.830 2.680 ;
        RECT 895.950 1.630 900.810 2.680 ;
        RECT 901.930 1.630 906.790 2.680 ;
        RECT 907.910 1.630 912.310 2.680 ;
        RECT 913.430 1.630 918.290 2.680 ;
        RECT 919.410 1.630 924.270 2.680 ;
        RECT 925.390 1.630 930.250 2.680 ;
        RECT 931.370 1.630 936.230 2.680 ;
        RECT 937.350 1.630 942.210 2.680 ;
        RECT 943.330 1.630 948.190 2.680 ;
        RECT 949.310 1.630 953.710 2.680 ;
        RECT 954.830 1.630 959.690 2.680 ;
        RECT 960.810 1.630 965.670 2.680 ;
        RECT 966.790 1.630 971.650 2.680 ;
        RECT 972.770 1.630 977.630 2.680 ;
        RECT 978.750 1.630 983.610 2.680 ;
        RECT 984.730 1.630 989.130 2.680 ;
        RECT 990.250 1.630 995.110 2.680 ;
        RECT 996.230 1.630 1001.090 2.680 ;
        RECT 1002.210 1.630 1007.070 2.680 ;
        RECT 1008.190 1.630 1013.050 2.680 ;
        RECT 1014.170 1.630 1019.030 2.680 ;
        RECT 1020.150 1.630 1025.010 2.680 ;
        RECT 1026.130 1.630 1030.530 2.680 ;
        RECT 1031.650 1.630 1036.510 2.680 ;
        RECT 1037.630 1.630 1042.490 2.680 ;
        RECT 1043.610 1.630 1048.470 2.680 ;
        RECT 1049.590 1.630 1054.450 2.680 ;
        RECT 1055.570 1.630 1060.430 2.680 ;
        RECT 1061.550 1.630 1066.410 2.680 ;
        RECT 1067.530 1.630 1071.930 2.680 ;
        RECT 1073.050 1.630 1077.910 2.680 ;
        RECT 1079.030 1.630 1083.890 2.680 ;
        RECT 1085.010 1.630 1089.870 2.680 ;
        RECT 1090.990 1.630 1095.850 2.680 ;
        RECT 1096.970 1.630 1101.830 2.680 ;
        RECT 1102.950 1.630 1107.350 2.680 ;
        RECT 1108.470 1.630 1113.330 2.680 ;
        RECT 1114.450 1.630 1119.310 2.680 ;
        RECT 1120.430 1.630 1125.290 2.680 ;
        RECT 1126.410 1.630 1131.270 2.680 ;
        RECT 1132.390 1.630 1137.250 2.680 ;
        RECT 1138.370 1.630 1143.230 2.680 ;
        RECT 1144.350 1.630 1148.750 2.680 ;
        RECT 1149.870 1.630 1154.730 2.680 ;
        RECT 1155.850 1.630 1160.710 2.680 ;
        RECT 1161.830 1.630 1166.690 2.680 ;
        RECT 1167.810 1.630 1172.670 2.680 ;
        RECT 1173.790 1.630 1178.650 2.680 ;
        RECT 1179.770 1.630 1184.630 2.680 ;
        RECT 1185.750 1.630 1190.150 2.680 ;
        RECT 1191.270 1.630 1196.130 2.680 ;
        RECT 1197.250 1.630 1202.110 2.680 ;
        RECT 1203.230 1.630 1208.090 2.680 ;
        RECT 1209.210 1.630 1214.070 2.680 ;
        RECT 1215.190 1.630 1220.050 2.680 ;
        RECT 1221.170 1.630 1225.570 2.680 ;
        RECT 1226.690 1.630 1231.550 2.680 ;
        RECT 1232.670 1.630 1237.530 2.680 ;
        RECT 1238.650 1.630 1243.510 2.680 ;
        RECT 1244.630 1.630 1249.490 2.680 ;
        RECT 1250.610 1.630 1255.470 2.680 ;
        RECT 1256.590 1.630 1261.450 2.680 ;
        RECT 1262.570 1.630 1266.970 2.680 ;
        RECT 1268.090 1.630 1272.950 2.680 ;
        RECT 1274.070 1.630 1278.930 2.680 ;
        RECT 1280.050 1.630 1284.910 2.680 ;
        RECT 1286.030 1.630 1290.890 2.680 ;
        RECT 1292.010 1.630 1296.870 2.680 ;
        RECT 1297.990 1.630 1302.850 2.680 ;
        RECT 1303.970 1.630 1308.370 2.680 ;
        RECT 1309.490 1.630 1314.350 2.680 ;
        RECT 1315.470 1.630 1320.330 2.680 ;
        RECT 1321.450 1.630 1326.310 2.680 ;
        RECT 1327.430 1.630 1332.290 2.680 ;
        RECT 1333.410 1.630 1338.270 2.680 ;
        RECT 1339.390 1.630 1343.790 2.680 ;
        RECT 1344.910 1.630 1349.770 2.680 ;
        RECT 1350.890 1.630 1355.750 2.680 ;
        RECT 1356.870 1.630 1361.730 2.680 ;
        RECT 1362.850 1.630 1367.710 2.680 ;
        RECT 1368.830 1.630 1373.690 2.680 ;
        RECT 1374.810 1.630 1379.670 2.680 ;
        RECT 1380.790 1.630 1385.190 2.680 ;
        RECT 1386.310 1.630 1391.170 2.680 ;
        RECT 1392.290 1.630 1397.150 2.680 ;
        RECT 1398.270 1.630 1403.130 2.680 ;
        RECT 1404.250 1.630 1409.110 2.680 ;
        RECT 1410.230 1.630 1415.090 2.680 ;
        RECT 1416.210 1.630 1421.070 2.680 ;
        RECT 1422.190 1.630 1426.590 2.680 ;
        RECT 1427.710 1.630 1432.570 2.680 ;
        RECT 1433.690 1.630 1438.550 2.680 ;
        RECT 1439.670 1.630 1444.530 2.680 ;
        RECT 1445.650 1.630 1450.510 2.680 ;
        RECT 1451.630 1.630 1456.490 2.680 ;
        RECT 1457.610 1.630 1462.470 2.680 ;
        RECT 1463.590 1.630 1467.990 2.680 ;
        RECT 1469.110 1.630 1473.970 2.680 ;
        RECT 1475.090 1.630 1479.950 2.680 ;
        RECT 1481.070 1.630 1485.930 2.680 ;
        RECT 1487.050 1.630 1491.910 2.680 ;
        RECT 1493.030 1.630 1497.890 2.680 ;
        RECT 1499.010 1.630 1503.410 2.680 ;
        RECT 1504.530 1.630 1509.390 2.680 ;
        RECT 1510.510 1.630 1515.370 2.680 ;
        RECT 1516.490 1.630 1521.350 2.680 ;
        RECT 1522.470 1.630 1527.330 2.680 ;
        RECT 1528.450 1.630 1533.310 2.680 ;
        RECT 1534.430 1.630 1539.290 2.680 ;
        RECT 1540.410 1.630 1544.810 2.680 ;
        RECT 1545.930 1.630 1550.790 2.680 ;
        RECT 1551.910 1.630 1556.770 2.680 ;
        RECT 1557.890 1.630 1562.750 2.680 ;
        RECT 1563.870 1.630 1568.730 2.680 ;
        RECT 1569.850 1.630 1574.710 2.680 ;
        RECT 1575.830 1.630 1580.690 2.680 ;
        RECT 1581.810 1.630 1586.210 2.680 ;
        RECT 1587.330 1.630 1592.190 2.680 ;
        RECT 1593.310 1.630 1598.170 2.680 ;
        RECT 1599.290 1.630 1604.150 2.680 ;
        RECT 1605.270 1.630 1610.130 2.680 ;
        RECT 1611.250 1.630 1616.110 2.680 ;
        RECT 1617.230 1.630 1621.630 2.680 ;
        RECT 1622.750 1.630 1627.610 2.680 ;
        RECT 1628.730 1.630 1633.590 2.680 ;
        RECT 1634.710 1.630 1639.570 2.680 ;
        RECT 1640.690 1.630 1645.550 2.680 ;
        RECT 1646.670 1.630 1651.530 2.680 ;
        RECT 1652.650 1.630 1657.510 2.680 ;
        RECT 1658.630 1.630 1663.030 2.680 ;
        RECT 1664.150 1.630 1669.010 2.680 ;
        RECT 1670.130 1.630 1674.990 2.680 ;
        RECT 1676.110 1.630 1680.970 2.680 ;
        RECT 1682.090 1.630 1686.950 2.680 ;
        RECT 1688.070 1.630 1692.930 2.680 ;
        RECT 1694.050 1.630 1698.910 2.680 ;
        RECT 1700.030 1.630 1704.430 2.680 ;
        RECT 1705.550 1.630 1710.410 2.680 ;
        RECT 1711.530 1.630 1716.390 2.680 ;
        RECT 1717.510 1.630 1722.370 2.680 ;
        RECT 1723.490 1.630 1728.350 2.680 ;
        RECT 1729.470 1.630 1734.330 2.680 ;
        RECT 1735.450 1.630 1739.850 2.680 ;
        RECT 1740.970 1.630 1745.830 2.680 ;
        RECT 1746.950 1.630 1751.810 2.680 ;
        RECT 1752.930 1.630 1757.790 2.680 ;
        RECT 1758.910 1.630 1763.770 2.680 ;
        RECT 1764.890 1.630 1769.750 2.680 ;
        RECT 1770.870 1.630 1775.730 2.680 ;
        RECT 1776.850 1.630 1781.250 2.680 ;
        RECT 1782.370 1.630 1787.230 2.680 ;
        RECT 1788.350 1.630 1793.210 2.680 ;
        RECT 1794.330 1.630 1799.190 2.680 ;
        RECT 1800.310 1.630 1805.170 2.680 ;
        RECT 1806.290 1.630 1811.150 2.680 ;
        RECT 1812.270 1.630 1817.130 2.680 ;
        RECT 1818.250 1.630 1822.650 2.680 ;
        RECT 1823.770 1.630 1828.630 2.680 ;
        RECT 1829.750 1.630 1834.610 2.680 ;
        RECT 1835.730 1.630 1840.590 2.680 ;
        RECT 1841.710 1.630 1846.570 2.680 ;
        RECT 1847.690 1.630 1852.550 2.680 ;
        RECT 1853.670 1.630 1858.070 2.680 ;
        RECT 1859.190 1.630 1864.050 2.680 ;
        RECT 1865.170 1.630 1870.030 2.680 ;
        RECT 1871.150 1.630 1876.010 2.680 ;
        RECT 1877.130 1.630 1881.990 2.680 ;
        RECT 1883.110 1.630 1887.970 2.680 ;
        RECT 1889.090 1.630 1893.950 2.680 ;
        RECT 1895.070 1.630 1899.470 2.680 ;
        RECT 1900.590 1.630 1905.450 2.680 ;
        RECT 1906.570 1.630 1911.430 2.680 ;
        RECT 1912.550 1.630 1917.410 2.680 ;
        RECT 1918.530 1.630 1923.390 2.680 ;
        RECT 1924.510 1.630 1929.370 2.680 ;
        RECT 1930.490 1.630 1935.350 2.680 ;
        RECT 1936.470 1.630 1940.870 2.680 ;
        RECT 1941.990 1.630 1946.850 2.680 ;
        RECT 1947.970 1.630 1952.830 2.680 ;
        RECT 1953.950 1.630 1958.810 2.680 ;
        RECT 1959.930 1.630 1964.790 2.680 ;
        RECT 1965.910 1.630 1970.770 2.680 ;
        RECT 1971.890 1.630 1976.290 2.680 ;
        RECT 1977.410 1.630 1982.270 2.680 ;
        RECT 1983.390 1.630 1988.250 2.680 ;
        RECT 1989.370 1.630 1994.230 2.680 ;
        RECT 1995.350 1.630 2000.210 2.680 ;
        RECT 2001.330 1.630 2006.190 2.680 ;
        RECT 2007.310 1.630 2012.170 2.680 ;
        RECT 2013.290 1.630 2017.690 2.680 ;
        RECT 2018.810 1.630 2023.670 2.680 ;
        RECT 2024.790 1.630 2029.650 2.680 ;
        RECT 2030.770 1.630 2035.630 2.680 ;
        RECT 2036.750 1.630 2041.610 2.680 ;
        RECT 2042.730 1.630 2047.590 2.680 ;
        RECT 2048.710 1.630 2053.570 2.680 ;
        RECT 2054.690 1.630 2059.090 2.680 ;
        RECT 2060.210 1.630 2065.070 2.680 ;
        RECT 2066.190 1.630 2071.050 2.680 ;
        RECT 2072.170 1.630 2077.030 2.680 ;
        RECT 2078.150 1.630 2083.010 2.680 ;
        RECT 2084.130 1.630 2088.990 2.680 ;
        RECT 2090.110 1.630 2094.510 2.680 ;
        RECT 2095.630 1.630 2100.490 2.680 ;
        RECT 2101.610 1.630 2106.470 2.680 ;
        RECT 2107.590 1.630 2112.450 2.680 ;
        RECT 2113.570 1.630 2118.430 2.680 ;
        RECT 2119.550 1.630 2124.410 2.680 ;
        RECT 2125.530 1.630 2130.390 2.680 ;
        RECT 2131.510 1.630 2135.910 2.680 ;
        RECT 2137.030 1.630 2141.890 2.680 ;
        RECT 2143.010 1.630 2147.870 2.680 ;
        RECT 2148.990 1.630 2153.850 2.680 ;
        RECT 2154.970 1.630 2159.830 2.680 ;
        RECT 2160.950 1.630 2165.810 2.680 ;
        RECT 2166.930 1.630 2171.790 2.680 ;
        RECT 2172.910 1.630 2177.310 2.680 ;
        RECT 2178.430 1.630 2183.290 2.680 ;
        RECT 2184.410 1.630 2189.270 2.680 ;
        RECT 2190.390 1.630 2195.250 2.680 ;
        RECT 2196.370 1.630 2201.230 2.680 ;
        RECT 2202.350 1.630 2207.210 2.680 ;
        RECT 2208.330 1.630 2212.730 2.680 ;
        RECT 2213.850 1.630 2218.710 2.680 ;
        RECT 2219.830 1.630 2224.690 2.680 ;
        RECT 2225.810 1.630 2230.670 2.680 ;
        RECT 2231.790 1.630 2236.650 2.680 ;
        RECT 2237.770 1.630 2242.630 2.680 ;
        RECT 2243.750 1.630 2248.610 2.680 ;
        RECT 2249.730 1.630 2254.130 2.680 ;
        RECT 2255.250 1.630 2260.110 2.680 ;
        RECT 2261.230 1.630 2266.090 2.680 ;
        RECT 2267.210 1.630 2272.070 2.680 ;
        RECT 2273.190 1.630 2278.050 2.680 ;
        RECT 2279.170 1.630 2284.030 2.680 ;
        RECT 2285.150 1.630 2290.010 2.680 ;
        RECT 2291.130 1.630 2295.530 2.680 ;
        RECT 2296.650 1.630 2301.510 2.680 ;
        RECT 2302.630 1.630 2307.490 2.680 ;
        RECT 2308.610 1.630 2313.470 2.680 ;
        RECT 2314.590 1.630 2319.450 2.680 ;
        RECT 2320.570 1.630 2325.430 2.680 ;
        RECT 2326.550 1.630 2330.950 2.680 ;
        RECT 2332.070 1.630 2336.930 2.680 ;
        RECT 2338.050 1.630 2342.910 2.680 ;
        RECT 2344.030 1.630 2348.890 2.680 ;
        RECT 2350.010 1.630 2354.870 2.680 ;
        RECT 2355.990 1.630 2360.850 2.680 ;
        RECT 2361.970 1.630 2366.830 2.680 ;
        RECT 2367.950 1.630 2372.350 2.680 ;
        RECT 2373.470 1.630 2378.330 2.680 ;
        RECT 2379.450 1.630 2384.310 2.680 ;
        RECT 2385.430 1.630 2390.290 2.680 ;
        RECT 2391.410 1.630 2396.270 2.680 ;
        RECT 2397.390 1.630 2402.250 2.680 ;
        RECT 2403.370 1.630 2408.230 2.680 ;
        RECT 2409.350 1.630 2413.750 2.680 ;
        RECT 2414.870 1.630 2419.730 2.680 ;
        RECT 2420.850 1.630 2425.710 2.680 ;
        RECT 2426.830 1.630 2431.690 2.680 ;
        RECT 2432.810 1.630 2437.670 2.680 ;
        RECT 2438.790 1.630 2443.650 2.680 ;
        RECT 2444.770 1.630 2449.170 2.680 ;
        RECT 2450.290 1.630 2455.150 2.680 ;
        RECT 2456.270 1.630 2461.130 2.680 ;
        RECT 2462.250 1.630 2467.110 2.680 ;
        RECT 2468.230 1.630 2473.090 2.680 ;
        RECT 2474.210 1.630 2479.070 2.680 ;
        RECT 2480.190 1.630 2485.050 2.680 ;
        RECT 2486.170 1.630 2490.570 2.680 ;
        RECT 2491.690 1.630 2496.550 2.680 ;
        RECT 2497.670 1.630 2502.530 2.680 ;
        RECT 2503.650 1.630 2508.510 2.680 ;
        RECT 2509.630 1.630 2514.490 2.680 ;
        RECT 2515.610 1.630 2520.470 2.680 ;
        RECT 2521.590 1.630 2526.450 2.680 ;
        RECT 2527.570 1.630 2531.970 2.680 ;
        RECT 2533.090 1.630 2537.950 2.680 ;
        RECT 2539.070 1.630 2543.930 2.680 ;
        RECT 2545.050 1.630 2549.910 2.680 ;
        RECT 2551.030 1.630 2555.890 2.680 ;
        RECT 2557.010 1.630 2561.870 2.680 ;
        RECT 2562.990 1.630 2567.390 2.680 ;
        RECT 2568.510 1.630 2573.370 2.680 ;
        RECT 2574.490 1.630 2579.350 2.680 ;
        RECT 2580.470 1.630 2585.330 2.680 ;
        RECT 2586.450 1.630 2591.310 2.680 ;
        RECT 2592.430 1.630 2597.290 2.680 ;
        RECT 2598.410 1.630 2603.270 2.680 ;
        RECT 2604.390 1.630 2608.790 2.680 ;
        RECT 2609.910 1.630 2614.770 2.680 ;
        RECT 2615.890 1.630 2620.750 2.680 ;
        RECT 2621.870 1.630 2626.730 2.680 ;
        RECT 2627.850 1.630 2632.710 2.680 ;
        RECT 2633.830 1.630 2638.690 2.680 ;
        RECT 2639.810 1.630 2644.670 2.680 ;
        RECT 2645.790 1.630 2650.190 2.680 ;
        RECT 2651.310 1.630 2656.170 2.680 ;
        RECT 2657.290 1.630 2662.150 2.680 ;
        RECT 2663.270 1.630 2668.130 2.680 ;
        RECT 2669.250 1.630 2674.110 2.680 ;
        RECT 2675.230 1.630 2680.090 2.680 ;
        RECT 2681.210 1.630 2685.610 2.680 ;
        RECT 2686.730 1.630 2691.590 2.680 ;
        RECT 2692.710 1.630 2697.570 2.680 ;
        RECT 2698.690 1.630 2703.550 2.680 ;
        RECT 2704.670 1.630 2709.530 2.680 ;
        RECT 2710.650 1.630 2715.510 2.680 ;
        RECT 2716.630 1.630 2721.490 2.680 ;
        RECT 2722.610 1.630 2727.010 2.680 ;
        RECT 2728.130 1.630 2732.990 2.680 ;
        RECT 2734.110 1.630 2738.970 2.680 ;
        RECT 2740.090 1.630 2744.950 2.680 ;
        RECT 2746.070 1.630 2750.930 2.680 ;
        RECT 2752.050 1.630 2756.910 2.680 ;
        RECT 2758.030 1.630 2762.890 2.680 ;
        RECT 2764.010 1.630 2768.410 2.680 ;
        RECT 2769.530 1.630 2774.390 2.680 ;
        RECT 2775.510 1.630 2780.370 2.680 ;
        RECT 2781.490 1.630 2786.350 2.680 ;
        RECT 2787.470 1.630 2792.330 2.680 ;
        RECT 2793.450 1.630 2798.310 2.680 ;
        RECT 2799.430 1.630 2803.830 2.680 ;
        RECT 2804.950 1.630 2809.810 2.680 ;
        RECT 2810.930 1.630 2815.790 2.680 ;
        RECT 2816.910 1.630 2821.770 2.680 ;
        RECT 2822.890 1.630 2827.750 2.680 ;
        RECT 2828.870 1.630 2833.730 2.680 ;
        RECT 2834.850 1.630 2839.710 2.680 ;
        RECT 2840.830 1.630 2845.230 2.680 ;
        RECT 2846.350 1.630 2851.210 2.680 ;
        RECT 2852.330 1.630 2857.190 2.680 ;
        RECT 2858.310 1.630 2863.170 2.680 ;
        RECT 2864.290 1.630 2869.150 2.680 ;
        RECT 2870.270 1.630 2875.130 2.680 ;
        RECT 2876.250 1.630 2881.110 2.680 ;
        RECT 2882.230 1.630 2886.630 2.680 ;
        RECT 2887.750 1.630 2892.610 2.680 ;
        RECT 2893.730 1.630 2898.590 2.680 ;
        RECT 2899.710 1.630 2904.570 2.680 ;
        RECT 2905.690 1.630 2910.550 2.680 ;
        RECT 2911.670 1.630 2916.530 2.680 ;
      LAYER met3 ;
        RECT 1.230 3487.700 2917.600 3501.825 ;
        RECT 2.800 3487.020 2917.600 3487.700 ;
        RECT 2.800 3485.700 2917.200 3487.020 ;
        RECT 1.230 3485.020 2917.200 3485.700 ;
        RECT 1.230 3422.420 2917.600 3485.020 ;
        RECT 2.800 3420.420 2917.600 3422.420 ;
        RECT 1.230 3420.380 2917.600 3420.420 ;
        RECT 1.230 3418.380 2917.200 3420.380 ;
        RECT 1.230 3357.140 2917.600 3418.380 ;
        RECT 2.800 3355.140 2917.600 3357.140 ;
        RECT 1.230 3354.420 2917.600 3355.140 ;
        RECT 1.230 3352.420 2917.200 3354.420 ;
        RECT 1.230 3291.860 2917.600 3352.420 ;
        RECT 2.800 3289.860 2917.600 3291.860 ;
        RECT 1.230 3287.780 2917.600 3289.860 ;
        RECT 1.230 3285.780 2917.200 3287.780 ;
        RECT 1.230 3226.580 2917.600 3285.780 ;
        RECT 2.800 3224.580 2917.600 3226.580 ;
        RECT 1.230 3221.140 2917.600 3224.580 ;
        RECT 1.230 3219.140 2917.200 3221.140 ;
        RECT 1.230 3161.300 2917.600 3219.140 ;
        RECT 2.800 3159.300 2917.600 3161.300 ;
        RECT 1.230 3155.180 2917.600 3159.300 ;
        RECT 1.230 3153.180 2917.200 3155.180 ;
        RECT 1.230 3096.700 2917.600 3153.180 ;
        RECT 2.800 3094.700 2917.600 3096.700 ;
        RECT 1.230 3088.540 2917.600 3094.700 ;
        RECT 1.230 3086.540 2917.200 3088.540 ;
        RECT 1.230 3031.420 2917.600 3086.540 ;
        RECT 2.800 3029.420 2917.600 3031.420 ;
        RECT 1.230 3021.900 2917.600 3029.420 ;
        RECT 1.230 3019.900 2917.200 3021.900 ;
        RECT 1.230 2966.140 2917.600 3019.900 ;
        RECT 2.800 2964.140 2917.600 2966.140 ;
        RECT 1.230 2955.940 2917.600 2964.140 ;
        RECT 1.230 2953.940 2917.200 2955.940 ;
        RECT 1.230 2900.860 2917.600 2953.940 ;
        RECT 2.800 2898.860 2917.600 2900.860 ;
        RECT 1.230 2889.300 2917.600 2898.860 ;
        RECT 1.230 2887.300 2917.200 2889.300 ;
        RECT 1.230 2835.580 2917.600 2887.300 ;
        RECT 2.800 2833.580 2917.600 2835.580 ;
        RECT 1.230 2822.660 2917.600 2833.580 ;
        RECT 1.230 2820.660 2917.200 2822.660 ;
        RECT 1.230 2770.300 2917.600 2820.660 ;
        RECT 2.800 2768.300 2917.600 2770.300 ;
        RECT 1.230 2756.700 2917.600 2768.300 ;
        RECT 1.230 2754.700 2917.200 2756.700 ;
        RECT 1.230 2705.020 2917.600 2754.700 ;
        RECT 2.800 2703.020 2917.600 2705.020 ;
        RECT 1.230 2690.060 2917.600 2703.020 ;
        RECT 1.230 2688.060 2917.200 2690.060 ;
        RECT 1.230 2640.420 2917.600 2688.060 ;
        RECT 2.800 2638.420 2917.600 2640.420 ;
        RECT 1.230 2623.420 2917.600 2638.420 ;
        RECT 1.230 2621.420 2917.200 2623.420 ;
        RECT 1.230 2575.140 2917.600 2621.420 ;
        RECT 2.800 2573.140 2917.600 2575.140 ;
        RECT 1.230 2557.460 2917.600 2573.140 ;
        RECT 1.230 2555.460 2917.200 2557.460 ;
        RECT 1.230 2509.860 2917.600 2555.460 ;
        RECT 2.800 2507.860 2917.600 2509.860 ;
        RECT 1.230 2490.820 2917.600 2507.860 ;
        RECT 1.230 2488.820 2917.200 2490.820 ;
        RECT 1.230 2444.580 2917.600 2488.820 ;
        RECT 2.800 2442.580 2917.600 2444.580 ;
        RECT 1.230 2424.180 2917.600 2442.580 ;
        RECT 1.230 2422.180 2917.200 2424.180 ;
        RECT 1.230 2379.300 2917.600 2422.180 ;
        RECT 2.800 2377.300 2917.600 2379.300 ;
        RECT 1.230 2358.220 2917.600 2377.300 ;
        RECT 1.230 2356.220 2917.200 2358.220 ;
        RECT 1.230 2314.020 2917.600 2356.220 ;
        RECT 2.800 2312.020 2917.600 2314.020 ;
        RECT 1.230 2291.580 2917.600 2312.020 ;
        RECT 1.230 2289.580 2917.200 2291.580 ;
        RECT 1.230 2248.740 2917.600 2289.580 ;
        RECT 2.800 2246.740 2917.600 2248.740 ;
        RECT 1.230 2224.940 2917.600 2246.740 ;
        RECT 1.230 2222.940 2917.200 2224.940 ;
        RECT 1.230 2184.140 2917.600 2222.940 ;
        RECT 2.800 2182.140 2917.600 2184.140 ;
        RECT 1.230 2158.980 2917.600 2182.140 ;
        RECT 1.230 2156.980 2917.200 2158.980 ;
        RECT 1.230 2118.860 2917.600 2156.980 ;
        RECT 2.800 2116.860 2917.600 2118.860 ;
        RECT 1.230 2092.340 2917.600 2116.860 ;
        RECT 1.230 2090.340 2917.200 2092.340 ;
        RECT 1.230 2053.580 2917.600 2090.340 ;
        RECT 2.800 2051.580 2917.600 2053.580 ;
        RECT 1.230 2025.700 2917.600 2051.580 ;
        RECT 1.230 2023.700 2917.200 2025.700 ;
        RECT 1.230 1988.300 2917.600 2023.700 ;
        RECT 2.800 1986.300 2917.600 1988.300 ;
        RECT 1.230 1959.740 2917.600 1986.300 ;
        RECT 1.230 1957.740 2917.200 1959.740 ;
        RECT 1.230 1923.020 2917.600 1957.740 ;
        RECT 2.800 1921.020 2917.600 1923.020 ;
        RECT 1.230 1893.100 2917.600 1921.020 ;
        RECT 1.230 1891.100 2917.200 1893.100 ;
        RECT 1.230 1857.740 2917.600 1891.100 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 1.230 1826.460 2917.600 1855.740 ;
        RECT 1.230 1824.460 2917.200 1826.460 ;
        RECT 1.230 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 1.230 1760.500 2917.600 1791.140 ;
        RECT 1.230 1758.500 2917.200 1760.500 ;
        RECT 1.230 1727.860 2917.600 1758.500 ;
        RECT 2.800 1725.860 2917.600 1727.860 ;
        RECT 1.230 1693.860 2917.600 1725.860 ;
        RECT 1.230 1691.860 2917.200 1693.860 ;
        RECT 1.230 1662.580 2917.600 1691.860 ;
        RECT 2.800 1660.580 2917.600 1662.580 ;
        RECT 1.230 1627.220 2917.600 1660.580 ;
        RECT 1.230 1625.220 2917.200 1627.220 ;
        RECT 1.230 1597.300 2917.600 1625.220 ;
        RECT 2.800 1595.300 2917.600 1597.300 ;
        RECT 1.230 1561.260 2917.600 1595.300 ;
        RECT 1.230 1559.260 2917.200 1561.260 ;
        RECT 1.230 1532.020 2917.600 1559.260 ;
        RECT 2.800 1530.020 2917.600 1532.020 ;
        RECT 1.230 1494.620 2917.600 1530.020 ;
        RECT 1.230 1492.620 2917.200 1494.620 ;
        RECT 1.230 1466.740 2917.600 1492.620 ;
        RECT 2.800 1464.740 2917.600 1466.740 ;
        RECT 1.230 1427.980 2917.600 1464.740 ;
        RECT 1.230 1425.980 2917.200 1427.980 ;
        RECT 1.230 1401.460 2917.600 1425.980 ;
        RECT 2.800 1399.460 2917.600 1401.460 ;
        RECT 1.230 1362.020 2917.600 1399.460 ;
        RECT 1.230 1360.020 2917.200 1362.020 ;
        RECT 1.230 1336.860 2917.600 1360.020 ;
        RECT 2.800 1334.860 2917.600 1336.860 ;
        RECT 1.230 1295.380 2917.600 1334.860 ;
        RECT 1.230 1293.380 2917.200 1295.380 ;
        RECT 1.230 1271.580 2917.600 1293.380 ;
        RECT 2.800 1269.580 2917.600 1271.580 ;
        RECT 1.230 1228.740 2917.600 1269.580 ;
        RECT 1.230 1226.740 2917.200 1228.740 ;
        RECT 1.230 1206.300 2917.600 1226.740 ;
        RECT 2.800 1204.300 2917.600 1206.300 ;
        RECT 1.230 1162.780 2917.600 1204.300 ;
        RECT 1.230 1160.780 2917.200 1162.780 ;
        RECT 1.230 1141.020 2917.600 1160.780 ;
        RECT 2.800 1139.020 2917.600 1141.020 ;
        RECT 1.230 1096.140 2917.600 1139.020 ;
        RECT 1.230 1094.140 2917.200 1096.140 ;
        RECT 1.230 1075.740 2917.600 1094.140 ;
        RECT 2.800 1073.740 2917.600 1075.740 ;
        RECT 1.230 1029.500 2917.600 1073.740 ;
        RECT 1.230 1027.500 2917.200 1029.500 ;
        RECT 1.230 1010.460 2917.600 1027.500 ;
        RECT 2.800 1008.460 2917.600 1010.460 ;
        RECT 1.230 963.540 2917.600 1008.460 ;
        RECT 1.230 961.540 2917.200 963.540 ;
        RECT 1.230 945.180 2917.600 961.540 ;
        RECT 2.800 943.180 2917.600 945.180 ;
        RECT 1.230 896.900 2917.600 943.180 ;
        RECT 1.230 894.900 2917.200 896.900 ;
        RECT 1.230 880.580 2917.600 894.900 ;
        RECT 2.800 878.580 2917.600 880.580 ;
        RECT 1.230 830.260 2917.600 878.580 ;
        RECT 1.230 828.260 2917.200 830.260 ;
        RECT 1.230 815.300 2917.600 828.260 ;
        RECT 2.800 813.300 2917.600 815.300 ;
        RECT 1.230 764.300 2917.600 813.300 ;
        RECT 1.230 762.300 2917.200 764.300 ;
        RECT 1.230 750.020 2917.600 762.300 ;
        RECT 2.800 748.020 2917.600 750.020 ;
        RECT 1.230 697.660 2917.600 748.020 ;
        RECT 1.230 695.660 2917.200 697.660 ;
        RECT 1.230 684.740 2917.600 695.660 ;
        RECT 2.800 682.740 2917.600 684.740 ;
        RECT 1.230 631.020 2917.600 682.740 ;
        RECT 1.230 629.020 2917.200 631.020 ;
        RECT 1.230 619.460 2917.600 629.020 ;
        RECT 2.800 617.460 2917.600 619.460 ;
        RECT 1.230 565.060 2917.600 617.460 ;
        RECT 1.230 563.060 2917.200 565.060 ;
        RECT 1.230 554.180 2917.600 563.060 ;
        RECT 2.800 552.180 2917.600 554.180 ;
        RECT 1.230 498.420 2917.600 552.180 ;
        RECT 1.230 496.420 2917.200 498.420 ;
        RECT 1.230 488.900 2917.600 496.420 ;
        RECT 2.800 486.900 2917.600 488.900 ;
        RECT 1.230 431.780 2917.600 486.900 ;
        RECT 1.230 429.780 2917.200 431.780 ;
        RECT 1.230 424.300 2917.600 429.780 ;
        RECT 2.800 422.300 2917.600 424.300 ;
        RECT 1.230 365.820 2917.600 422.300 ;
        RECT 1.230 363.820 2917.200 365.820 ;
        RECT 1.230 359.020 2917.600 363.820 ;
        RECT 2.800 357.020 2917.600 359.020 ;
        RECT 1.230 299.180 2917.600 357.020 ;
        RECT 1.230 297.180 2917.200 299.180 ;
        RECT 1.230 293.740 2917.600 297.180 ;
        RECT 2.800 291.740 2917.600 293.740 ;
        RECT 1.230 232.540 2917.600 291.740 ;
        RECT 1.230 230.540 2917.200 232.540 ;
        RECT 1.230 228.460 2917.600 230.540 ;
        RECT 2.800 226.460 2917.600 228.460 ;
        RECT 1.230 166.580 2917.600 226.460 ;
        RECT 1.230 164.580 2917.200 166.580 ;
        RECT 1.230 163.180 2917.600 164.580 ;
        RECT 2.800 161.180 2917.600 163.180 ;
        RECT 1.230 99.940 2917.600 161.180 ;
        RECT 1.230 97.940 2917.200 99.940 ;
        RECT 1.230 97.900 2917.600 97.940 ;
        RECT 2.800 95.900 2917.600 97.900 ;
        RECT 1.230 33.980 2917.600 95.900 ;
        RECT 1.230 33.300 2917.200 33.980 ;
        RECT 2.800 32.135 2917.200 33.300 ;
      LAYER met4 ;
        RECT 150.620 3376.140 158.570 3501.825 ;
        RECT 162.470 3376.140 164.370 3501.825 ;
        RECT 168.270 3376.140 177.170 3501.825 ;
        RECT 181.070 3376.140 195.770 3501.825 ;
        RECT 199.670 3376.140 208.570 3501.825 ;
        RECT 212.470 3376.140 214.370 3501.825 ;
        RECT 218.270 3376.140 227.170 3501.825 ;
        RECT 231.070 3376.140 245.770 3501.825 ;
        RECT 249.670 3376.140 258.570 3501.825 ;
        RECT 262.470 3376.140 264.370 3501.825 ;
        RECT 268.270 3376.140 277.170 3501.825 ;
        RECT 281.070 3376.140 295.770 3501.825 ;
        RECT 299.670 3376.140 308.570 3501.825 ;
        RECT 312.470 3376.140 314.370 3501.825 ;
        RECT 318.270 3376.140 327.170 3501.825 ;
        RECT 331.070 3376.140 345.770 3501.825 ;
        RECT 349.670 3376.140 358.570 3501.825 ;
        RECT 362.470 3376.140 364.370 3501.825 ;
        RECT 368.270 3376.140 377.170 3501.825 ;
        RECT 381.070 3376.140 395.770 3501.825 ;
        RECT 399.670 3376.140 408.570 3501.825 ;
        RECT 412.470 3376.140 414.370 3501.825 ;
        RECT 418.270 3376.140 427.170 3501.825 ;
        RECT 431.070 3376.140 445.770 3501.825 ;
        RECT 449.670 3376.140 458.570 3501.825 ;
        RECT 462.470 3376.140 464.370 3501.825 ;
        RECT 468.270 3376.140 477.170 3501.825 ;
        RECT 481.070 3376.140 495.770 3501.825 ;
        RECT 499.670 3376.140 508.570 3501.825 ;
        RECT 512.470 3376.140 514.370 3501.825 ;
        RECT 518.270 3376.140 527.170 3501.825 ;
        RECT 531.070 3376.140 545.770 3501.825 ;
        RECT 549.670 3376.140 558.570 3501.825 ;
        RECT 562.470 3376.140 564.370 3501.825 ;
        RECT 568.270 3376.140 577.170 3501.825 ;
        RECT 581.070 3376.140 595.770 3501.825 ;
        RECT 599.670 3376.140 608.570 3501.825 ;
        RECT 612.470 3376.140 614.370 3501.825 ;
        RECT 618.270 3376.140 627.170 3501.825 ;
        RECT 631.070 3376.140 645.770 3501.825 ;
        RECT 649.670 3376.140 658.570 3501.825 ;
        RECT 662.470 3376.140 664.370 3501.825 ;
        RECT 668.270 3376.140 677.170 3501.825 ;
        RECT 681.070 3376.140 695.770 3501.825 ;
        RECT 699.670 3376.140 708.570 3501.825 ;
        RECT 712.470 3376.140 714.370 3501.825 ;
        RECT 718.270 3376.140 727.170 3501.825 ;
        RECT 731.070 3376.140 745.770 3501.825 ;
        RECT 749.670 3376.140 758.570 3501.825 ;
        RECT 762.470 3376.140 764.370 3501.825 ;
        RECT 768.270 3376.140 777.170 3501.825 ;
        RECT 781.070 3376.140 795.770 3501.825 ;
        RECT 799.670 3376.140 808.570 3501.825 ;
        RECT 812.470 3376.140 814.370 3501.825 ;
        RECT 818.270 3376.140 827.170 3501.825 ;
        RECT 831.070 3376.140 845.770 3501.825 ;
        RECT 150.620 2940.400 845.770 3376.140 ;
        RECT 150.620 2816.140 158.570 2940.400 ;
        RECT 162.470 2816.140 164.370 2940.400 ;
        RECT 168.270 2816.140 177.170 2940.400 ;
        RECT 181.070 2816.140 195.770 2940.400 ;
        RECT 199.670 2816.140 208.570 2940.400 ;
        RECT 212.470 2816.140 214.370 2940.400 ;
        RECT 218.270 2816.140 227.170 2940.400 ;
        RECT 231.070 2816.140 245.770 2940.400 ;
        RECT 249.670 2816.140 258.570 2940.400 ;
        RECT 262.470 2816.140 264.370 2940.400 ;
        RECT 268.270 2816.140 277.170 2940.400 ;
        RECT 281.070 2816.140 295.770 2940.400 ;
        RECT 299.670 2816.140 308.570 2940.400 ;
        RECT 312.470 2816.140 314.370 2940.400 ;
        RECT 318.270 2816.140 327.170 2940.400 ;
        RECT 331.070 2816.140 345.770 2940.400 ;
        RECT 349.670 2816.140 358.570 2940.400 ;
        RECT 362.470 2816.140 364.370 2940.400 ;
        RECT 368.270 2816.140 377.170 2940.400 ;
        RECT 381.070 2816.140 395.770 2940.400 ;
        RECT 399.670 2816.140 408.570 2940.400 ;
        RECT 412.470 2816.140 414.370 2940.400 ;
        RECT 418.270 2816.140 427.170 2940.400 ;
        RECT 431.070 2816.140 445.770 2940.400 ;
        RECT 449.670 2816.140 458.570 2940.400 ;
        RECT 462.470 2816.140 464.370 2940.400 ;
        RECT 468.270 2816.140 477.170 2940.400 ;
        RECT 481.070 2816.140 495.770 2940.400 ;
        RECT 499.670 2816.140 508.570 2940.400 ;
        RECT 512.470 2816.140 514.370 2940.400 ;
        RECT 518.270 2816.140 527.170 2940.400 ;
        RECT 531.070 2816.140 545.770 2940.400 ;
        RECT 549.670 2816.140 558.570 2940.400 ;
        RECT 562.470 2816.140 564.370 2940.400 ;
        RECT 568.270 2816.140 577.170 2940.400 ;
        RECT 581.070 2816.140 595.770 2940.400 ;
        RECT 599.670 2816.140 608.570 2940.400 ;
        RECT 612.470 2816.140 614.370 2940.400 ;
        RECT 618.270 2816.140 627.170 2940.400 ;
        RECT 631.070 2816.140 645.770 2940.400 ;
        RECT 649.670 2816.140 658.570 2940.400 ;
        RECT 662.470 2816.140 664.370 2940.400 ;
        RECT 668.270 2816.140 677.170 2940.400 ;
        RECT 681.070 2816.140 695.770 2940.400 ;
        RECT 699.670 2816.140 708.570 2940.400 ;
        RECT 712.470 2816.140 714.370 2940.400 ;
        RECT 718.270 2816.140 727.170 2940.400 ;
        RECT 731.070 2816.140 745.770 2940.400 ;
        RECT 749.670 2816.140 758.570 2940.400 ;
        RECT 762.470 2816.140 764.370 2940.400 ;
        RECT 768.270 2816.140 777.170 2940.400 ;
        RECT 781.070 2816.140 795.770 2940.400 ;
        RECT 799.670 2816.140 808.570 2940.400 ;
        RECT 812.470 2816.140 814.370 2940.400 ;
        RECT 818.270 2816.140 827.170 2940.400 ;
        RECT 831.070 2816.140 845.770 2940.400 ;
        RECT 150.620 2380.400 845.770 2816.140 ;
        RECT 150.620 2256.140 158.570 2380.400 ;
        RECT 162.470 2256.140 164.370 2380.400 ;
        RECT 168.270 2256.140 177.170 2380.400 ;
        RECT 181.070 2256.140 195.770 2380.400 ;
        RECT 199.670 2256.140 208.570 2380.400 ;
        RECT 212.470 2256.140 214.370 2380.400 ;
        RECT 218.270 2256.140 227.170 2380.400 ;
        RECT 231.070 2256.140 245.770 2380.400 ;
        RECT 249.670 2256.140 258.570 2380.400 ;
        RECT 262.470 2256.140 264.370 2380.400 ;
        RECT 268.270 2256.140 277.170 2380.400 ;
        RECT 281.070 2256.140 295.770 2380.400 ;
        RECT 299.670 2256.140 308.570 2380.400 ;
        RECT 312.470 2256.140 314.370 2380.400 ;
        RECT 318.270 2256.140 327.170 2380.400 ;
        RECT 331.070 2256.140 345.770 2380.400 ;
        RECT 349.670 2256.140 358.570 2380.400 ;
        RECT 362.470 2256.140 364.370 2380.400 ;
        RECT 368.270 2256.140 377.170 2380.400 ;
        RECT 381.070 2256.140 395.770 2380.400 ;
        RECT 399.670 2256.140 408.570 2380.400 ;
        RECT 412.470 2256.140 414.370 2380.400 ;
        RECT 418.270 2256.140 427.170 2380.400 ;
        RECT 431.070 2256.140 445.770 2380.400 ;
        RECT 449.670 2256.140 458.570 2380.400 ;
        RECT 462.470 2256.140 464.370 2380.400 ;
        RECT 468.270 2256.140 477.170 2380.400 ;
        RECT 481.070 2256.140 495.770 2380.400 ;
        RECT 499.670 2256.140 508.570 2380.400 ;
        RECT 512.470 2256.140 514.370 2380.400 ;
        RECT 518.270 2256.140 527.170 2380.400 ;
        RECT 531.070 2256.140 545.770 2380.400 ;
        RECT 549.670 2256.140 558.570 2380.400 ;
        RECT 562.470 2256.140 564.370 2380.400 ;
        RECT 568.270 2256.140 577.170 2380.400 ;
        RECT 581.070 2256.140 595.770 2380.400 ;
        RECT 599.670 2256.140 608.570 2380.400 ;
        RECT 612.470 2256.140 614.370 2380.400 ;
        RECT 618.270 2256.140 627.170 2380.400 ;
        RECT 631.070 2256.140 645.770 2380.400 ;
        RECT 649.670 2256.140 658.570 2380.400 ;
        RECT 662.470 2256.140 664.370 2380.400 ;
        RECT 668.270 2256.140 677.170 2380.400 ;
        RECT 681.070 2256.140 695.770 2380.400 ;
        RECT 699.670 2256.140 708.570 2380.400 ;
        RECT 712.470 2256.140 714.370 2380.400 ;
        RECT 718.270 2256.140 727.170 2380.400 ;
        RECT 731.070 2256.140 745.770 2380.400 ;
        RECT 749.670 2256.140 758.570 2380.400 ;
        RECT 762.470 2256.140 764.370 2380.400 ;
        RECT 768.270 2256.140 777.170 2380.400 ;
        RECT 781.070 2256.140 795.770 2380.400 ;
        RECT 799.670 2256.140 808.570 2380.400 ;
        RECT 812.470 2256.140 814.370 2380.400 ;
        RECT 818.270 2256.140 827.170 2380.400 ;
        RECT 831.070 2256.140 845.770 2380.400 ;
        RECT 150.620 1820.400 845.770 2256.140 ;
        RECT 150.620 1696.140 158.570 1820.400 ;
        RECT 162.470 1696.140 164.370 1820.400 ;
        RECT 168.270 1696.140 177.170 1820.400 ;
        RECT 181.070 1696.140 195.770 1820.400 ;
        RECT 199.670 1696.140 208.570 1820.400 ;
        RECT 212.470 1696.140 214.370 1820.400 ;
        RECT 218.270 1696.140 227.170 1820.400 ;
        RECT 231.070 1696.140 245.770 1820.400 ;
        RECT 249.670 1696.140 258.570 1820.400 ;
        RECT 262.470 1696.140 264.370 1820.400 ;
        RECT 268.270 1696.140 277.170 1820.400 ;
        RECT 281.070 1696.140 295.770 1820.400 ;
        RECT 299.670 1696.140 308.570 1820.400 ;
        RECT 312.470 1696.140 314.370 1820.400 ;
        RECT 318.270 1696.140 327.170 1820.400 ;
        RECT 331.070 1696.140 345.770 1820.400 ;
        RECT 349.670 1696.140 358.570 1820.400 ;
        RECT 362.470 1696.140 364.370 1820.400 ;
        RECT 368.270 1696.140 377.170 1820.400 ;
        RECT 381.070 1696.140 395.770 1820.400 ;
        RECT 399.670 1696.140 408.570 1820.400 ;
        RECT 412.470 1696.140 414.370 1820.400 ;
        RECT 418.270 1696.140 427.170 1820.400 ;
        RECT 431.070 1696.140 445.770 1820.400 ;
        RECT 449.670 1696.140 458.570 1820.400 ;
        RECT 462.470 1696.140 464.370 1820.400 ;
        RECT 468.270 1696.140 477.170 1820.400 ;
        RECT 481.070 1696.140 495.770 1820.400 ;
        RECT 499.670 1696.140 508.570 1820.400 ;
        RECT 512.470 1696.140 514.370 1820.400 ;
        RECT 518.270 1696.140 527.170 1820.400 ;
        RECT 531.070 1696.140 545.770 1820.400 ;
        RECT 549.670 1696.140 558.570 1820.400 ;
        RECT 562.470 1696.140 564.370 1820.400 ;
        RECT 568.270 1696.140 577.170 1820.400 ;
        RECT 581.070 1696.140 595.770 1820.400 ;
        RECT 599.670 1696.140 608.570 1820.400 ;
        RECT 612.470 1696.140 614.370 1820.400 ;
        RECT 618.270 1696.140 627.170 1820.400 ;
        RECT 631.070 1696.140 645.770 1820.400 ;
        RECT 649.670 1696.140 658.570 1820.400 ;
        RECT 662.470 1696.140 664.370 1820.400 ;
        RECT 668.270 1696.140 677.170 1820.400 ;
        RECT 681.070 1696.140 695.770 1820.400 ;
        RECT 699.670 1696.140 708.570 1820.400 ;
        RECT 712.470 1696.140 714.370 1820.400 ;
        RECT 718.270 1696.140 727.170 1820.400 ;
        RECT 731.070 1696.140 745.770 1820.400 ;
        RECT 749.670 1696.140 758.570 1820.400 ;
        RECT 762.470 1696.140 764.370 1820.400 ;
        RECT 768.270 1696.140 777.170 1820.400 ;
        RECT 781.070 1696.140 795.770 1820.400 ;
        RECT 799.670 1696.140 808.570 1820.400 ;
        RECT 812.470 1696.140 814.370 1820.400 ;
        RECT 818.270 1696.140 827.170 1820.400 ;
        RECT 831.070 1696.140 845.770 1820.400 ;
        RECT 150.620 1260.400 845.770 1696.140 ;
        RECT 150.620 1136.140 158.570 1260.400 ;
        RECT 162.470 1136.140 164.370 1260.400 ;
        RECT 168.270 1136.140 177.170 1260.400 ;
        RECT 181.070 1136.140 195.770 1260.400 ;
        RECT 199.670 1136.140 208.570 1260.400 ;
        RECT 212.470 1136.140 214.370 1260.400 ;
        RECT 218.270 1136.140 227.170 1260.400 ;
        RECT 231.070 1136.140 245.770 1260.400 ;
        RECT 249.670 1136.140 258.570 1260.400 ;
        RECT 262.470 1136.140 264.370 1260.400 ;
        RECT 268.270 1136.140 277.170 1260.400 ;
        RECT 281.070 1136.140 295.770 1260.400 ;
        RECT 299.670 1136.140 308.570 1260.400 ;
        RECT 312.470 1136.140 314.370 1260.400 ;
        RECT 318.270 1136.140 327.170 1260.400 ;
        RECT 331.070 1136.140 345.770 1260.400 ;
        RECT 349.670 1136.140 358.570 1260.400 ;
        RECT 362.470 1136.140 364.370 1260.400 ;
        RECT 368.270 1136.140 377.170 1260.400 ;
        RECT 381.070 1136.140 395.770 1260.400 ;
        RECT 399.670 1136.140 408.570 1260.400 ;
        RECT 412.470 1136.140 414.370 1260.400 ;
        RECT 418.270 1136.140 427.170 1260.400 ;
        RECT 431.070 1136.140 445.770 1260.400 ;
        RECT 449.670 1136.140 458.570 1260.400 ;
        RECT 462.470 1136.140 464.370 1260.400 ;
        RECT 468.270 1136.140 477.170 1260.400 ;
        RECT 481.070 1136.140 495.770 1260.400 ;
        RECT 499.670 1136.140 508.570 1260.400 ;
        RECT 512.470 1136.140 514.370 1260.400 ;
        RECT 518.270 1136.140 527.170 1260.400 ;
        RECT 531.070 1136.140 545.770 1260.400 ;
        RECT 549.670 1136.140 558.570 1260.400 ;
        RECT 562.470 1136.140 564.370 1260.400 ;
        RECT 568.270 1136.140 577.170 1260.400 ;
        RECT 581.070 1136.140 595.770 1260.400 ;
        RECT 599.670 1136.140 608.570 1260.400 ;
        RECT 612.470 1136.140 614.370 1260.400 ;
        RECT 618.270 1136.140 627.170 1260.400 ;
        RECT 631.070 1136.140 645.770 1260.400 ;
        RECT 649.670 1136.140 658.570 1260.400 ;
        RECT 662.470 1136.140 664.370 1260.400 ;
        RECT 668.270 1136.140 677.170 1260.400 ;
        RECT 681.070 1136.140 695.770 1260.400 ;
        RECT 699.670 1136.140 708.570 1260.400 ;
        RECT 712.470 1136.140 714.370 1260.400 ;
        RECT 718.270 1136.140 727.170 1260.400 ;
        RECT 731.070 1136.140 745.770 1260.400 ;
        RECT 749.670 1136.140 758.570 1260.400 ;
        RECT 762.470 1136.140 764.370 1260.400 ;
        RECT 768.270 1136.140 777.170 1260.400 ;
        RECT 781.070 1136.140 795.770 1260.400 ;
        RECT 799.670 1136.140 808.570 1260.400 ;
        RECT 812.470 1136.140 814.370 1260.400 ;
        RECT 818.270 1136.140 827.170 1260.400 ;
        RECT 831.070 1136.140 845.770 1260.400 ;
        RECT 150.620 700.400 845.770 1136.140 ;
        RECT 150.620 576.140 158.570 700.400 ;
        RECT 162.470 576.140 164.370 700.400 ;
        RECT 168.270 576.140 177.170 700.400 ;
        RECT 181.070 576.140 195.770 700.400 ;
        RECT 199.670 576.140 208.570 700.400 ;
        RECT 212.470 576.140 214.370 700.400 ;
        RECT 218.270 576.140 227.170 700.400 ;
        RECT 231.070 576.140 245.770 700.400 ;
        RECT 249.670 576.140 258.570 700.400 ;
        RECT 262.470 576.140 264.370 700.400 ;
        RECT 268.270 576.140 277.170 700.400 ;
        RECT 281.070 576.140 295.770 700.400 ;
        RECT 299.670 576.140 308.570 700.400 ;
        RECT 312.470 576.140 314.370 700.400 ;
        RECT 318.270 576.140 327.170 700.400 ;
        RECT 331.070 576.140 345.770 700.400 ;
        RECT 349.670 576.140 358.570 700.400 ;
        RECT 362.470 576.140 364.370 700.400 ;
        RECT 368.270 576.140 377.170 700.400 ;
        RECT 381.070 576.140 395.770 700.400 ;
        RECT 399.670 576.140 408.570 700.400 ;
        RECT 412.470 576.140 414.370 700.400 ;
        RECT 418.270 576.140 427.170 700.400 ;
        RECT 431.070 576.140 445.770 700.400 ;
        RECT 449.670 576.140 458.570 700.400 ;
        RECT 462.470 576.140 464.370 700.400 ;
        RECT 468.270 576.140 477.170 700.400 ;
        RECT 481.070 576.140 495.770 700.400 ;
        RECT 499.670 576.140 508.570 700.400 ;
        RECT 512.470 576.140 514.370 700.400 ;
        RECT 518.270 576.140 527.170 700.400 ;
        RECT 531.070 576.140 545.770 700.400 ;
        RECT 549.670 576.140 558.570 700.400 ;
        RECT 562.470 576.140 564.370 700.400 ;
        RECT 568.270 576.140 577.170 700.400 ;
        RECT 581.070 576.140 595.770 700.400 ;
        RECT 599.670 576.140 608.570 700.400 ;
        RECT 612.470 576.140 614.370 700.400 ;
        RECT 618.270 576.140 627.170 700.400 ;
        RECT 631.070 576.140 645.770 700.400 ;
        RECT 649.670 576.140 658.570 700.400 ;
        RECT 662.470 576.140 664.370 700.400 ;
        RECT 668.270 576.140 677.170 700.400 ;
        RECT 681.070 576.140 695.770 700.400 ;
        RECT 699.670 576.140 708.570 700.400 ;
        RECT 712.470 576.140 714.370 700.400 ;
        RECT 718.270 576.140 727.170 700.400 ;
        RECT 731.070 576.140 745.770 700.400 ;
        RECT 749.670 576.140 758.570 700.400 ;
        RECT 762.470 576.140 764.370 700.400 ;
        RECT 768.270 576.140 777.170 700.400 ;
        RECT 781.070 576.140 795.770 700.400 ;
        RECT 799.670 576.140 808.570 700.400 ;
        RECT 812.470 576.140 814.370 700.400 ;
        RECT 818.270 576.140 827.170 700.400 ;
        RECT 831.070 576.140 845.770 700.400 ;
        RECT 150.620 140.400 845.770 576.140 ;
        RECT 150.620 132.095 158.570 140.400 ;
        RECT 162.470 132.095 164.370 140.400 ;
        RECT 168.270 132.095 177.170 140.400 ;
        RECT 181.070 132.095 195.770 140.400 ;
        RECT 199.670 132.095 208.570 140.400 ;
        RECT 212.470 132.095 214.370 140.400 ;
        RECT 218.270 132.095 227.170 140.400 ;
        RECT 231.070 132.095 245.770 140.400 ;
        RECT 249.670 132.095 258.570 140.400 ;
        RECT 262.470 132.095 264.370 140.400 ;
        RECT 268.270 132.095 277.170 140.400 ;
        RECT 281.070 132.095 295.770 140.400 ;
        RECT 299.670 132.095 308.570 140.400 ;
        RECT 312.470 132.095 314.370 140.400 ;
        RECT 318.270 132.095 327.170 140.400 ;
        RECT 331.070 132.095 345.770 140.400 ;
        RECT 349.670 132.095 358.570 140.400 ;
        RECT 362.470 132.095 364.370 140.400 ;
        RECT 368.270 132.095 377.170 140.400 ;
        RECT 381.070 132.095 395.770 140.400 ;
        RECT 399.670 132.095 408.570 140.400 ;
        RECT 412.470 132.095 414.370 140.400 ;
        RECT 418.270 132.095 427.170 140.400 ;
        RECT 431.070 132.095 445.770 140.400 ;
        RECT 449.670 132.095 458.570 140.400 ;
        RECT 462.470 132.095 464.370 140.400 ;
        RECT 468.270 132.095 477.170 140.400 ;
        RECT 481.070 132.095 495.770 140.400 ;
        RECT 499.670 132.095 508.570 140.400 ;
        RECT 512.470 132.095 514.370 140.400 ;
        RECT 518.270 132.095 527.170 140.400 ;
        RECT 531.070 132.095 545.770 140.400 ;
        RECT 549.670 132.095 558.570 140.400 ;
        RECT 562.470 132.095 564.370 140.400 ;
        RECT 568.270 132.095 577.170 140.400 ;
        RECT 581.070 132.095 595.770 140.400 ;
        RECT 599.670 132.095 608.570 140.400 ;
        RECT 612.470 132.095 614.370 140.400 ;
        RECT 618.270 132.095 627.170 140.400 ;
        RECT 631.070 132.095 645.770 140.400 ;
        RECT 649.670 132.095 658.570 140.400 ;
        RECT 662.470 132.095 664.370 140.400 ;
        RECT 668.270 132.095 677.170 140.400 ;
        RECT 681.070 132.095 695.770 140.400 ;
        RECT 699.670 132.095 708.570 140.400 ;
        RECT 712.470 132.095 714.370 140.400 ;
        RECT 718.270 132.095 727.170 140.400 ;
        RECT 731.070 132.095 745.770 140.400 ;
        RECT 749.670 132.095 758.570 140.400 ;
        RECT 762.470 132.095 764.370 140.400 ;
        RECT 768.270 132.095 777.170 140.400 ;
        RECT 781.070 132.095 795.770 140.400 ;
        RECT 799.670 132.095 808.570 140.400 ;
        RECT 812.470 132.095 814.370 140.400 ;
        RECT 818.270 132.095 827.170 140.400 ;
        RECT 831.070 132.095 845.770 140.400 ;
        RECT 849.670 132.095 858.570 3501.825 ;
        RECT 862.470 132.095 864.370 3501.825 ;
        RECT 868.270 132.095 877.170 3501.825 ;
        RECT 881.070 132.095 895.770 3501.825 ;
        RECT 899.670 132.095 908.570 3501.825 ;
        RECT 912.470 132.095 914.370 3501.825 ;
        RECT 918.270 132.095 927.170 3501.825 ;
        RECT 931.070 132.095 945.770 3501.825 ;
        RECT 949.670 132.095 958.570 3501.825 ;
        RECT 962.470 132.095 964.370 3501.825 ;
        RECT 968.270 132.095 977.170 3501.825 ;
        RECT 981.070 2696.140 995.770 3501.825 ;
        RECT 999.670 2696.140 1008.570 3501.825 ;
        RECT 1012.470 2696.140 1014.370 3501.825 ;
        RECT 1018.270 2696.140 1027.170 3501.825 ;
        RECT 1031.070 2696.140 1045.770 3501.825 ;
        RECT 1049.670 2696.140 1058.570 3501.825 ;
        RECT 1062.470 2696.140 1064.370 3501.825 ;
        RECT 1068.270 2696.140 1077.170 3501.825 ;
        RECT 1081.070 2696.140 1095.770 3501.825 ;
        RECT 1099.670 2696.140 1108.570 3501.825 ;
        RECT 1112.470 2696.140 1114.370 3501.825 ;
        RECT 1118.270 2696.140 1127.170 3501.825 ;
        RECT 1131.070 2696.140 1145.770 3501.825 ;
        RECT 1149.670 2696.140 1158.570 3501.825 ;
        RECT 1162.470 2696.140 1164.370 3501.825 ;
        RECT 1168.270 2696.140 1177.170 3501.825 ;
        RECT 1181.070 3297.100 1195.770 3501.825 ;
        RECT 1199.670 3297.100 1208.570 3501.825 ;
        RECT 1212.470 3297.100 1214.370 3501.825 ;
        RECT 1218.270 3297.100 1227.170 3501.825 ;
        RECT 1231.070 3297.100 1245.770 3501.825 ;
        RECT 1249.670 3297.100 1258.570 3501.825 ;
        RECT 1262.470 3297.100 1264.370 3501.825 ;
        RECT 1268.270 3297.100 1277.170 3501.825 ;
        RECT 1281.070 3297.100 1295.770 3501.825 ;
        RECT 1299.670 3297.100 1308.570 3501.825 ;
        RECT 1312.470 3297.100 1314.370 3501.825 ;
        RECT 1318.270 3297.100 1327.170 3501.825 ;
        RECT 1331.070 3297.100 1345.770 3501.825 ;
        RECT 1349.670 3297.100 1358.570 3501.825 ;
        RECT 1362.470 3297.100 1364.370 3501.825 ;
        RECT 1368.270 3297.100 1377.170 3501.825 ;
        RECT 1381.070 3297.100 1395.770 3501.825 ;
        RECT 1399.670 3297.100 1408.570 3501.825 ;
        RECT 1412.470 3297.100 1414.370 3501.825 ;
        RECT 1418.270 3297.100 1427.170 3501.825 ;
        RECT 1431.070 3297.100 1445.770 3501.825 ;
        RECT 1449.670 3297.100 1458.570 3501.825 ;
        RECT 1462.470 3297.100 1464.370 3501.825 ;
        RECT 1468.270 3297.100 1477.170 3501.825 ;
        RECT 1481.070 3297.100 1495.770 3501.825 ;
        RECT 1499.670 3297.100 1508.570 3501.825 ;
        RECT 1512.470 3297.100 1514.370 3501.825 ;
        RECT 1518.270 3297.100 1527.170 3501.825 ;
        RECT 1531.070 3297.100 1545.770 3501.825 ;
        RECT 1549.670 3297.100 1558.570 3501.825 ;
        RECT 1562.470 3297.100 1564.370 3501.825 ;
        RECT 1568.270 3297.100 1577.170 3501.825 ;
        RECT 1581.070 3297.100 1595.770 3501.825 ;
        RECT 1599.670 3297.100 1608.570 3501.825 ;
        RECT 1612.470 3297.100 1614.370 3501.825 ;
        RECT 1618.270 3297.100 1627.170 3501.825 ;
        RECT 1631.070 3297.100 1645.770 3501.825 ;
        RECT 1649.670 3297.100 1658.570 3501.825 ;
        RECT 1662.470 3297.100 1664.370 3501.825 ;
        RECT 1668.270 3297.100 1677.170 3501.825 ;
        RECT 1681.070 3297.100 1695.770 3501.825 ;
        RECT 1181.070 2880.400 1695.770 3297.100 ;
        RECT 1181.070 2696.140 1195.770 2880.400 ;
        RECT 1199.670 2696.140 1208.570 2880.400 ;
        RECT 1212.470 2696.140 1214.370 2880.400 ;
        RECT 1218.270 2696.140 1227.170 2880.400 ;
        RECT 1231.070 2696.140 1245.770 2880.400 ;
        RECT 1249.670 2696.140 1258.570 2880.400 ;
        RECT 1262.470 2696.140 1264.370 2880.400 ;
        RECT 1268.270 2696.140 1277.170 2880.400 ;
        RECT 1281.070 2696.140 1295.770 2880.400 ;
        RECT 1299.670 2696.140 1308.570 2880.400 ;
        RECT 1312.470 2696.140 1314.370 2880.400 ;
        RECT 1318.270 2696.140 1327.170 2880.400 ;
        RECT 1331.070 2696.140 1345.770 2880.400 ;
        RECT 1349.670 2696.140 1358.570 2880.400 ;
        RECT 1362.470 2696.140 1364.370 2880.400 ;
        RECT 1368.270 2696.140 1377.170 2880.400 ;
        RECT 1381.070 2696.140 1395.770 2880.400 ;
        RECT 1399.670 2696.140 1408.570 2880.400 ;
        RECT 1412.470 2696.140 1414.370 2880.400 ;
        RECT 1418.270 2696.140 1427.170 2880.400 ;
        RECT 1431.070 2696.140 1445.770 2880.400 ;
        RECT 1449.670 2696.140 1458.570 2880.400 ;
        RECT 1462.470 2696.140 1464.370 2880.400 ;
        RECT 1468.270 2696.140 1477.170 2880.400 ;
        RECT 1481.070 2696.140 1495.770 2880.400 ;
        RECT 1499.670 2696.140 1508.570 2880.400 ;
        RECT 1512.470 2696.140 1514.370 2880.400 ;
        RECT 1518.270 2696.140 1527.170 2880.400 ;
        RECT 1531.070 2696.140 1545.770 2880.400 ;
        RECT 1549.670 2696.140 1558.570 2880.400 ;
        RECT 1562.470 2696.140 1564.370 2880.400 ;
        RECT 1568.270 2696.140 1577.170 2880.400 ;
        RECT 1581.070 2696.140 1595.770 2880.400 ;
        RECT 1599.670 2696.140 1608.570 2880.400 ;
        RECT 1612.470 2696.140 1614.370 2880.400 ;
        RECT 1618.270 2696.140 1627.170 2880.400 ;
        RECT 1631.070 2696.140 1645.770 2880.400 ;
        RECT 1649.670 2696.140 1658.570 2880.400 ;
        RECT 1662.470 2696.140 1664.370 2880.400 ;
        RECT 1668.270 2696.140 1677.170 2880.400 ;
        RECT 1681.070 2696.140 1695.770 2880.400 ;
        RECT 981.070 2260.400 1695.770 2696.140 ;
        RECT 981.070 2076.700 995.770 2260.400 ;
        RECT 999.670 2076.700 1008.570 2260.400 ;
        RECT 1012.470 2076.700 1014.370 2260.400 ;
        RECT 1018.270 2076.700 1027.170 2260.400 ;
        RECT 1031.070 2076.700 1045.770 2260.400 ;
        RECT 1049.670 2076.700 1058.570 2260.400 ;
        RECT 1062.470 2076.700 1064.370 2260.400 ;
        RECT 1068.270 2076.700 1077.170 2260.400 ;
        RECT 1081.070 2076.700 1095.770 2260.400 ;
        RECT 1099.670 2076.700 1108.570 2260.400 ;
        RECT 1112.470 2076.700 1114.370 2260.400 ;
        RECT 1118.270 2076.700 1127.170 2260.400 ;
        RECT 1131.070 2076.700 1145.770 2260.400 ;
        RECT 1149.670 2076.700 1158.570 2260.400 ;
        RECT 1162.470 2076.700 1164.370 2260.400 ;
        RECT 1168.270 2076.700 1177.170 2260.400 ;
        RECT 1181.070 2076.700 1195.770 2260.400 ;
        RECT 1199.670 2076.700 1208.570 2260.400 ;
        RECT 1212.470 2076.700 1214.370 2260.400 ;
        RECT 1218.270 2076.700 1227.170 2260.400 ;
        RECT 1231.070 2076.700 1245.770 2260.400 ;
        RECT 1249.670 2076.700 1258.570 2260.400 ;
        RECT 1262.470 2076.700 1264.370 2260.400 ;
        RECT 1268.270 2076.700 1277.170 2260.400 ;
        RECT 1281.070 2076.700 1295.770 2260.400 ;
        RECT 1299.670 2076.700 1308.570 2260.400 ;
        RECT 1312.470 2076.700 1314.370 2260.400 ;
        RECT 1318.270 2076.700 1327.170 2260.400 ;
        RECT 1331.070 2076.700 1345.770 2260.400 ;
        RECT 1349.670 2076.700 1358.570 2260.400 ;
        RECT 1362.470 2076.700 1364.370 2260.400 ;
        RECT 1368.270 2076.700 1377.170 2260.400 ;
        RECT 1381.070 2076.700 1395.770 2260.400 ;
        RECT 1399.670 2076.700 1408.570 2260.400 ;
        RECT 1412.470 2076.700 1414.370 2260.400 ;
        RECT 1418.270 2076.700 1427.170 2260.400 ;
        RECT 1431.070 2076.700 1445.770 2260.400 ;
        RECT 1449.670 2076.700 1458.570 2260.400 ;
        RECT 1462.470 2076.700 1464.370 2260.400 ;
        RECT 1468.270 2076.700 1477.170 2260.400 ;
        RECT 1481.070 2076.700 1495.770 2260.400 ;
        RECT 1499.670 2076.700 1508.570 2260.400 ;
        RECT 1512.470 2076.700 1514.370 2260.400 ;
        RECT 1518.270 2076.700 1527.170 2260.400 ;
        RECT 1531.070 2076.700 1545.770 2260.400 ;
        RECT 1549.670 2076.700 1558.570 2260.400 ;
        RECT 1562.470 2076.700 1564.370 2260.400 ;
        RECT 1568.270 2076.700 1577.170 2260.400 ;
        RECT 1581.070 2076.700 1595.770 2260.400 ;
        RECT 1599.670 2076.700 1608.570 2260.400 ;
        RECT 1612.470 2076.700 1614.370 2260.400 ;
        RECT 1618.270 2076.700 1627.170 2260.400 ;
        RECT 1631.070 2076.700 1645.770 2260.400 ;
        RECT 1649.670 2076.700 1658.570 2260.400 ;
        RECT 1662.470 2076.700 1664.370 2260.400 ;
        RECT 1668.270 2076.700 1677.170 2260.400 ;
        RECT 1681.070 2076.700 1695.770 2260.400 ;
        RECT 1699.670 2076.700 1708.570 3501.825 ;
        RECT 1712.470 2076.700 1714.370 3501.825 ;
        RECT 1718.270 2076.700 1727.170 3501.825 ;
        RECT 1731.070 2076.700 1745.770 3501.825 ;
        RECT 1749.670 2076.700 1758.570 3501.825 ;
        RECT 1762.470 2076.700 1764.370 3501.825 ;
        RECT 1768.270 2076.700 1777.170 3501.825 ;
        RECT 1781.070 2076.700 1795.770 3501.825 ;
        RECT 1799.670 2076.700 1808.570 3501.825 ;
        RECT 1812.470 2076.700 1814.370 3501.825 ;
        RECT 1818.270 2076.700 1827.170 3501.825 ;
        RECT 1831.070 2076.700 1845.770 3501.825 ;
        RECT 1849.670 2076.700 1858.570 3501.825 ;
        RECT 1862.470 2076.700 1864.370 3501.825 ;
        RECT 1868.270 2076.700 1877.170 3501.825 ;
        RECT 1881.070 2076.700 1895.770 3501.825 ;
        RECT 1899.670 2076.700 1908.570 3501.825 ;
        RECT 1912.470 2076.700 1914.370 3501.825 ;
        RECT 1918.270 2076.700 1927.170 3501.825 ;
        RECT 1931.070 2076.700 1945.770 3501.825 ;
        RECT 1949.670 2076.700 1958.570 3501.825 ;
        RECT 1962.470 2076.700 1964.370 3501.825 ;
        RECT 1968.270 2076.700 1977.170 3501.825 ;
        RECT 1981.070 2076.700 1995.770 3501.825 ;
        RECT 1999.670 2076.700 2008.570 3501.825 ;
        RECT 2012.470 2076.700 2014.370 3501.825 ;
        RECT 2018.270 2076.700 2027.170 3501.825 ;
        RECT 2031.070 3297.100 2045.770 3501.825 ;
        RECT 2049.670 3297.100 2058.570 3501.825 ;
        RECT 2062.470 3297.100 2064.370 3501.825 ;
        RECT 2068.270 3297.100 2077.170 3501.825 ;
        RECT 2081.070 3297.100 2095.770 3501.825 ;
        RECT 2099.670 3297.100 2108.570 3501.825 ;
        RECT 2112.470 3297.100 2114.370 3501.825 ;
        RECT 2118.270 3297.100 2127.170 3501.825 ;
        RECT 2131.070 3297.100 2145.770 3501.825 ;
        RECT 2149.670 3297.100 2158.570 3501.825 ;
        RECT 2162.470 3297.100 2164.370 3501.825 ;
        RECT 2168.270 3297.100 2177.170 3501.825 ;
        RECT 2181.070 3297.100 2195.770 3501.825 ;
        RECT 2199.670 3297.100 2208.570 3501.825 ;
        RECT 2212.470 3297.100 2214.370 3501.825 ;
        RECT 2218.270 3297.100 2227.170 3501.825 ;
        RECT 2231.070 3297.100 2245.770 3501.825 ;
        RECT 2249.670 3297.100 2258.570 3501.825 ;
        RECT 2262.470 3297.100 2264.370 3501.825 ;
        RECT 2268.270 3297.100 2277.170 3501.825 ;
        RECT 2281.070 3297.100 2295.770 3501.825 ;
        RECT 2299.670 3297.100 2308.570 3501.825 ;
        RECT 2312.470 3297.100 2314.370 3501.825 ;
        RECT 2318.270 3297.100 2327.170 3501.825 ;
        RECT 2331.070 3297.100 2345.770 3501.825 ;
        RECT 2349.670 3297.100 2358.570 3501.825 ;
        RECT 2362.470 3297.100 2364.370 3501.825 ;
        RECT 2368.270 3297.100 2377.170 3501.825 ;
        RECT 2381.070 3297.100 2395.770 3501.825 ;
        RECT 2399.670 3297.100 2408.570 3501.825 ;
        RECT 2412.470 3297.100 2414.370 3501.825 ;
        RECT 2418.270 3297.100 2427.170 3501.825 ;
        RECT 2431.070 3297.100 2445.770 3501.825 ;
        RECT 2449.670 3297.100 2458.570 3501.825 ;
        RECT 2462.470 3297.100 2464.370 3501.825 ;
        RECT 2468.270 3297.100 2477.170 3501.825 ;
        RECT 2481.070 3297.100 2495.770 3501.825 ;
        RECT 2499.670 3297.100 2508.570 3501.825 ;
        RECT 2512.470 3297.100 2514.370 3501.825 ;
        RECT 2518.270 3297.100 2527.170 3501.825 ;
        RECT 2531.070 3297.100 2545.770 3501.825 ;
        RECT 2031.070 2880.400 2545.770 3297.100 ;
        RECT 2031.070 2696.140 2045.770 2880.400 ;
        RECT 2049.670 2696.140 2058.570 2880.400 ;
        RECT 2062.470 2696.140 2064.370 2880.400 ;
        RECT 2068.270 2696.140 2077.170 2880.400 ;
        RECT 2081.070 2696.140 2095.770 2880.400 ;
        RECT 2099.670 2696.140 2108.570 2880.400 ;
        RECT 2112.470 2696.140 2114.370 2880.400 ;
        RECT 2118.270 2696.140 2127.170 2880.400 ;
        RECT 2131.070 2696.140 2145.770 2880.400 ;
        RECT 2149.670 2696.140 2158.570 2880.400 ;
        RECT 2162.470 2696.140 2164.370 2880.400 ;
        RECT 2168.270 2696.140 2177.170 2880.400 ;
        RECT 2181.070 2696.140 2195.770 2880.400 ;
        RECT 2199.670 2696.140 2208.570 2880.400 ;
        RECT 2212.470 2696.140 2214.370 2880.400 ;
        RECT 2218.270 2696.140 2227.170 2880.400 ;
        RECT 2231.070 2696.140 2245.770 2880.400 ;
        RECT 2249.670 2696.140 2258.570 2880.400 ;
        RECT 2262.470 2696.140 2264.370 2880.400 ;
        RECT 2268.270 2696.140 2277.170 2880.400 ;
        RECT 2281.070 2696.140 2295.770 2880.400 ;
        RECT 2299.670 2696.140 2308.570 2880.400 ;
        RECT 2312.470 2696.140 2314.370 2880.400 ;
        RECT 2318.270 2696.140 2327.170 2880.400 ;
        RECT 2331.070 2696.140 2345.770 2880.400 ;
        RECT 2349.670 2696.140 2358.570 2880.400 ;
        RECT 2362.470 2696.140 2364.370 2880.400 ;
        RECT 2368.270 2696.140 2377.170 2880.400 ;
        RECT 2381.070 2696.140 2395.770 2880.400 ;
        RECT 2399.670 2696.140 2408.570 2880.400 ;
        RECT 2412.470 2696.140 2414.370 2880.400 ;
        RECT 2418.270 2696.140 2427.170 2880.400 ;
        RECT 2431.070 2696.140 2445.770 2880.400 ;
        RECT 2449.670 2696.140 2458.570 2880.400 ;
        RECT 2462.470 2696.140 2464.370 2880.400 ;
        RECT 2468.270 2696.140 2477.170 2880.400 ;
        RECT 2481.070 2696.140 2495.770 2880.400 ;
        RECT 2499.670 2696.140 2508.570 2880.400 ;
        RECT 2512.470 2696.140 2514.370 2880.400 ;
        RECT 2518.270 2696.140 2527.170 2880.400 ;
        RECT 2531.070 2696.140 2545.770 2880.400 ;
        RECT 2549.670 2696.140 2558.570 3501.825 ;
        RECT 2562.470 2696.140 2564.370 3501.825 ;
        RECT 2568.270 2696.140 2577.170 3501.825 ;
        RECT 2581.070 2696.140 2595.770 3501.825 ;
        RECT 2599.670 2696.140 2608.570 3501.825 ;
        RECT 2612.470 2696.140 2614.370 3501.825 ;
        RECT 2618.270 2696.140 2627.170 3501.825 ;
        RECT 2631.070 2696.140 2645.770 3501.825 ;
        RECT 2649.670 2696.140 2658.570 3501.825 ;
        RECT 2662.470 2696.140 2664.370 3501.825 ;
        RECT 2668.270 2696.140 2677.170 3501.825 ;
        RECT 2681.070 2696.140 2695.770 3501.825 ;
        RECT 2699.670 2696.140 2708.570 3501.825 ;
        RECT 2712.470 2696.140 2714.370 3501.825 ;
        RECT 2718.270 2696.140 2727.170 3501.825 ;
        RECT 2731.070 2696.140 2732.480 3501.825 ;
        RECT 2031.070 2260.400 2732.480 2696.140 ;
        RECT 2031.070 2076.700 2045.770 2260.400 ;
        RECT 2049.670 2076.700 2058.570 2260.400 ;
        RECT 2062.470 2076.700 2064.370 2260.400 ;
        RECT 2068.270 2076.700 2077.170 2260.400 ;
        RECT 2081.070 2076.700 2095.770 2260.400 ;
        RECT 2099.670 2076.700 2108.570 2260.400 ;
        RECT 2112.470 2076.700 2114.370 2260.400 ;
        RECT 2118.270 2076.700 2127.170 2260.400 ;
        RECT 2131.070 2076.700 2145.770 2260.400 ;
        RECT 2149.670 2076.700 2158.570 2260.400 ;
        RECT 2162.470 2076.700 2164.370 2260.400 ;
        RECT 2168.270 2076.700 2177.170 2260.400 ;
        RECT 2181.070 2076.700 2195.770 2260.400 ;
        RECT 2199.670 2076.700 2208.570 2260.400 ;
        RECT 2212.470 2076.700 2214.370 2260.400 ;
        RECT 2218.270 2076.700 2227.170 2260.400 ;
        RECT 2231.070 2076.700 2245.770 2260.400 ;
        RECT 2249.670 2076.700 2258.570 2260.400 ;
        RECT 2262.470 2076.700 2264.370 2260.400 ;
        RECT 2268.270 2076.700 2277.170 2260.400 ;
        RECT 2281.070 2076.700 2295.770 2260.400 ;
        RECT 2299.670 2076.700 2308.570 2260.400 ;
        RECT 2312.470 2076.700 2314.370 2260.400 ;
        RECT 2318.270 2076.700 2327.170 2260.400 ;
        RECT 2331.070 2076.700 2345.770 2260.400 ;
        RECT 2349.670 2076.700 2358.570 2260.400 ;
        RECT 2362.470 2076.700 2364.370 2260.400 ;
        RECT 2368.270 2076.700 2377.170 2260.400 ;
        RECT 2381.070 2076.700 2395.770 2260.400 ;
        RECT 2399.670 2076.700 2408.570 2260.400 ;
        RECT 2412.470 2076.700 2414.370 2260.400 ;
        RECT 2418.270 2076.700 2427.170 2260.400 ;
        RECT 2431.070 2076.700 2445.770 2260.400 ;
        RECT 2449.670 2076.700 2458.570 2260.400 ;
        RECT 2462.470 2076.700 2464.370 2260.400 ;
        RECT 2468.270 2076.700 2477.170 2260.400 ;
        RECT 2481.070 2076.700 2495.770 2260.400 ;
        RECT 2499.670 2076.700 2508.570 2260.400 ;
        RECT 2512.470 2076.700 2514.370 2260.400 ;
        RECT 2518.270 2076.700 2527.170 2260.400 ;
        RECT 2531.070 2076.700 2545.770 2260.400 ;
        RECT 2549.670 2076.700 2558.570 2260.400 ;
        RECT 2562.470 2076.700 2564.370 2260.400 ;
        RECT 2568.270 2076.700 2577.170 2260.400 ;
        RECT 2581.070 2076.700 2595.770 2260.400 ;
        RECT 2599.670 2076.700 2608.570 2260.400 ;
        RECT 2612.470 2076.700 2614.370 2260.400 ;
        RECT 2618.270 2076.700 2627.170 2260.400 ;
        RECT 2631.070 2076.700 2645.770 2260.400 ;
        RECT 2649.670 2076.700 2658.570 2260.400 ;
        RECT 2662.470 2076.700 2664.370 2260.400 ;
        RECT 2668.270 2076.700 2677.170 2260.400 ;
        RECT 2681.070 2076.700 2695.770 2260.400 ;
        RECT 2699.670 2076.700 2708.570 2260.400 ;
        RECT 2712.470 2076.700 2714.370 2260.400 ;
        RECT 2718.270 2076.700 2727.170 2260.400 ;
        RECT 2731.070 2076.700 2732.480 2260.400 ;
        RECT 981.070 290.400 2732.480 2076.700 ;
        RECT 981.070 132.095 995.770 290.400 ;
        RECT 999.670 132.095 1008.570 290.400 ;
        RECT 1012.470 132.095 1014.370 290.400 ;
        RECT 1018.270 132.095 1027.170 290.400 ;
        RECT 1031.070 132.095 1045.770 290.400 ;
        RECT 1049.670 132.095 1058.570 290.400 ;
        RECT 1062.470 132.095 1064.370 290.400 ;
        RECT 1068.270 132.095 1077.170 290.400 ;
        RECT 1081.070 132.095 1095.770 290.400 ;
        RECT 1099.670 132.095 1108.570 290.400 ;
        RECT 1112.470 132.095 1114.370 290.400 ;
        RECT 1118.270 132.095 1127.170 290.400 ;
        RECT 1131.070 132.095 1145.770 290.400 ;
        RECT 1149.670 132.095 1158.570 290.400 ;
        RECT 1162.470 132.095 1164.370 290.400 ;
        RECT 1168.270 132.095 1177.170 290.400 ;
        RECT 1181.070 132.095 1195.770 290.400 ;
        RECT 1199.670 132.095 1208.570 290.400 ;
        RECT 1212.470 132.095 1214.370 290.400 ;
        RECT 1218.270 132.095 1227.170 290.400 ;
        RECT 1231.070 132.095 1245.770 290.400 ;
        RECT 1249.670 132.095 1258.570 290.400 ;
        RECT 1262.470 132.095 1264.370 290.400 ;
        RECT 1268.270 132.095 1277.170 290.400 ;
        RECT 1281.070 132.095 1295.770 290.400 ;
        RECT 1299.670 132.095 1308.570 290.400 ;
        RECT 1312.470 132.095 1314.370 290.400 ;
        RECT 1318.270 132.095 1327.170 290.400 ;
        RECT 1331.070 132.095 1345.770 290.400 ;
        RECT 1349.670 132.095 1358.570 290.400 ;
        RECT 1362.470 132.095 1364.370 290.400 ;
        RECT 1368.270 132.095 1377.170 290.400 ;
        RECT 1381.070 132.095 1395.770 290.400 ;
        RECT 1399.670 132.095 1408.570 290.400 ;
        RECT 1412.470 132.095 1414.370 290.400 ;
        RECT 1418.270 132.095 1427.170 290.400 ;
        RECT 1431.070 132.095 1445.770 290.400 ;
        RECT 1449.670 132.095 1458.570 290.400 ;
        RECT 1462.470 132.095 1464.370 290.400 ;
        RECT 1468.270 132.095 1477.170 290.400 ;
        RECT 1481.070 132.095 1495.770 290.400 ;
        RECT 1499.670 132.095 1508.570 290.400 ;
        RECT 1512.470 132.095 1514.370 290.400 ;
        RECT 1518.270 132.095 1527.170 290.400 ;
        RECT 1531.070 132.095 1545.770 290.400 ;
        RECT 1549.670 132.095 1558.570 290.400 ;
        RECT 1562.470 132.095 1564.370 290.400 ;
        RECT 1568.270 132.095 1577.170 290.400 ;
        RECT 1581.070 132.095 1595.770 290.400 ;
        RECT 1599.670 132.095 1608.570 290.400 ;
        RECT 1612.470 132.095 1614.370 290.400 ;
        RECT 1618.270 132.095 1627.170 290.400 ;
        RECT 1631.070 132.095 1645.770 290.400 ;
        RECT 1649.670 132.095 1658.570 290.400 ;
        RECT 1662.470 132.095 1664.370 290.400 ;
        RECT 1668.270 132.095 1677.170 290.400 ;
        RECT 1681.070 132.095 1695.770 290.400 ;
        RECT 1699.670 132.095 1708.570 290.400 ;
        RECT 1712.470 132.095 1714.370 290.400 ;
        RECT 1718.270 132.095 1727.170 290.400 ;
        RECT 1731.070 132.095 1745.770 290.400 ;
        RECT 1749.670 132.095 1758.570 290.400 ;
        RECT 1762.470 132.095 1764.370 290.400 ;
        RECT 1768.270 132.095 1777.170 290.400 ;
        RECT 1781.070 132.095 1795.770 290.400 ;
        RECT 1799.670 132.095 1808.570 290.400 ;
        RECT 1812.470 132.095 1814.370 290.400 ;
        RECT 1818.270 132.095 1827.170 290.400 ;
        RECT 1831.070 132.095 1845.770 290.400 ;
        RECT 1849.670 132.095 1858.570 290.400 ;
        RECT 1862.470 132.095 1864.370 290.400 ;
        RECT 1868.270 132.095 1877.170 290.400 ;
        RECT 1881.070 132.095 1895.770 290.400 ;
        RECT 1899.670 132.095 1908.570 290.400 ;
        RECT 1912.470 132.095 1914.370 290.400 ;
        RECT 1918.270 132.095 1927.170 290.400 ;
        RECT 1931.070 132.095 1945.770 290.400 ;
        RECT 1949.670 132.095 1958.570 290.400 ;
        RECT 1962.470 132.095 1964.370 290.400 ;
        RECT 1968.270 132.095 1977.170 290.400 ;
        RECT 1981.070 132.095 1995.770 290.400 ;
        RECT 1999.670 132.095 2008.570 290.400 ;
        RECT 2012.470 132.095 2014.370 290.400 ;
        RECT 2018.270 132.095 2027.170 290.400 ;
        RECT 2031.070 132.095 2045.770 290.400 ;
        RECT 2049.670 132.095 2058.570 290.400 ;
        RECT 2062.470 132.095 2064.370 290.400 ;
        RECT 2068.270 132.095 2077.170 290.400 ;
        RECT 2081.070 132.095 2095.770 290.400 ;
        RECT 2099.670 132.095 2108.570 290.400 ;
        RECT 2112.470 132.095 2114.370 290.400 ;
        RECT 2118.270 132.095 2127.170 290.400 ;
        RECT 2131.070 132.095 2145.770 290.400 ;
        RECT 2149.670 132.095 2158.570 290.400 ;
        RECT 2162.470 132.095 2164.370 290.400 ;
        RECT 2168.270 132.095 2177.170 290.400 ;
        RECT 2181.070 132.095 2195.770 290.400 ;
        RECT 2199.670 132.095 2208.570 290.400 ;
        RECT 2212.470 132.095 2214.370 290.400 ;
        RECT 2218.270 132.095 2227.170 290.400 ;
        RECT 2231.070 132.095 2245.770 290.400 ;
        RECT 2249.670 132.095 2258.570 290.400 ;
        RECT 2262.470 132.095 2264.370 290.400 ;
        RECT 2268.270 132.095 2277.170 290.400 ;
        RECT 2281.070 132.095 2295.770 290.400 ;
        RECT 2299.670 132.095 2308.570 290.400 ;
        RECT 2312.470 132.095 2314.370 290.400 ;
        RECT 2318.270 132.095 2327.170 290.400 ;
        RECT 2331.070 132.095 2345.770 290.400 ;
        RECT 2349.670 132.095 2358.570 290.400 ;
        RECT 2362.470 132.095 2364.370 290.400 ;
        RECT 2368.270 132.095 2377.170 290.400 ;
        RECT 2381.070 132.095 2395.770 290.400 ;
        RECT 2399.670 132.095 2408.570 290.400 ;
        RECT 2412.470 132.095 2414.370 290.400 ;
        RECT 2418.270 132.095 2427.170 290.400 ;
        RECT 2431.070 132.095 2445.770 290.400 ;
        RECT 2449.670 132.095 2458.570 290.400 ;
        RECT 2462.470 132.095 2464.370 290.400 ;
        RECT 2468.270 132.095 2477.170 290.400 ;
        RECT 2481.070 132.095 2495.770 290.400 ;
        RECT 2499.670 132.095 2508.570 290.400 ;
        RECT 2512.470 132.095 2514.370 290.400 ;
        RECT 2518.270 132.095 2527.170 290.400 ;
        RECT 2531.070 132.095 2545.770 290.400 ;
        RECT 2549.670 132.095 2558.570 290.400 ;
        RECT 2562.470 132.095 2564.370 290.400 ;
        RECT 2568.270 132.095 2577.170 290.400 ;
        RECT 2581.070 132.095 2595.770 290.400 ;
        RECT 2599.670 132.095 2608.570 290.400 ;
        RECT 2612.470 132.095 2614.370 290.400 ;
        RECT 2618.270 132.095 2627.170 290.400 ;
        RECT 2631.070 132.095 2645.770 290.400 ;
        RECT 2649.670 132.095 2658.570 290.400 ;
        RECT 2662.470 132.095 2664.370 290.400 ;
        RECT 2668.270 132.095 2677.170 290.400 ;
        RECT 2681.070 132.095 2695.770 290.400 ;
        RECT 2699.670 132.095 2708.570 290.400 ;
        RECT 2712.470 132.095 2714.370 290.400 ;
        RECT 2718.270 132.095 2727.170 290.400 ;
        RECT 2731.070 132.095 2732.480 290.400 ;
  END
END user_project_wrapper
END LIBRARY

