VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Marmot
  CLASS BLOCK ;
  FOREIGN Marmot ;
  ORIGIN 0.000 0.000 ;
  SIZE 1767.600 BY 1778.320 ;
  PIN data_arrays_0_0_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END data_arrays_0_0_ext_ram_addr1[0]
  PIN data_arrays_0_0_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END data_arrays_0_0_ext_ram_addr1[1]
  PIN data_arrays_0_0_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 772.520 4.000 773.120 ;
    END
  END data_arrays_0_0_ext_ram_addr1[2]
  PIN data_arrays_0_0_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.920 4.000 776.520 ;
    END
  END data_arrays_0_0_ext_ram_addr1[3]
  PIN data_arrays_0_0_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END data_arrays_0_0_ext_ram_addr1[4]
  PIN data_arrays_0_0_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END data_arrays_0_0_ext_ram_addr1[5]
  PIN data_arrays_0_0_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END data_arrays_0_0_ext_ram_addr1[6]
  PIN data_arrays_0_0_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 789.520 4.000 790.120 ;
    END
  END data_arrays_0_0_ext_ram_addr1[7]
  PIN data_arrays_0_0_ext_ram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 793.600 4.000 794.200 ;
    END
  END data_arrays_0_0_ext_ram_addr1[8]
  PIN data_arrays_0_0_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END data_arrays_0_0_ext_ram_addr[0]
  PIN data_arrays_0_0_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END data_arrays_0_0_ext_ram_addr[1]
  PIN data_arrays_0_0_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END data_arrays_0_0_ext_ram_addr[2]
  PIN data_arrays_0_0_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END data_arrays_0_0_ext_ram_addr[3]
  PIN data_arrays_0_0_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END data_arrays_0_0_ext_ram_addr[4]
  PIN data_arrays_0_0_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END data_arrays_0_0_ext_ram_addr[5]
  PIN data_arrays_0_0_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END data_arrays_0_0_ext_ram_addr[6]
  PIN data_arrays_0_0_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END data_arrays_0_0_ext_ram_addr[7]
  PIN data_arrays_0_0_ext_ram_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END data_arrays_0_0_ext_ram_addr[8]
  PIN data_arrays_0_0_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 483.520 4.000 484.120 ;
    END
  END data_arrays_0_0_ext_ram_clk
  PIN data_arrays_0_0_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END data_arrays_0_0_ext_ram_csb1[0]
  PIN data_arrays_0_0_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 740.560 4.000 741.160 ;
    END
  END data_arrays_0_0_ext_ram_csb1[1]
  PIN data_arrays_0_0_ext_ram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END data_arrays_0_0_ext_ram_csb1[2]
  PIN data_arrays_0_0_ext_ram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 747.360 4.000 747.960 ;
    END
  END data_arrays_0_0_ext_ram_csb1[3]
  PIN data_arrays_0_0_ext_ram_csb1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.760 4.000 751.360 ;
    END
  END data_arrays_0_0_ext_ram_csb1[4]
  PIN data_arrays_0_0_ext_ram_csb1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END data_arrays_0_0_ext_ram_csb1[5]
  PIN data_arrays_0_0_ext_ram_csb1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END data_arrays_0_0_ext_ram_csb1[6]
  PIN data_arrays_0_0_ext_ram_csb1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END data_arrays_0_0_ext_ram_csb1[7]
  PIN data_arrays_0_0_ext_ram_csb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END data_arrays_0_0_ext_ram_csb[0]
  PIN data_arrays_0_0_ext_ram_csb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END data_arrays_0_0_ext_ram_csb[1]
  PIN data_arrays_0_0_ext_ram_csb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END data_arrays_0_0_ext_ram_csb[2]
  PIN data_arrays_0_0_ext_ram_csb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END data_arrays_0_0_ext_ram_csb[3]
  PIN data_arrays_0_0_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[0]
  PIN data_arrays_0_0_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[10]
  PIN data_arrays_0_0_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[11]
  PIN data_arrays_0_0_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[12]
  PIN data_arrays_0_0_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[13]
  PIN data_arrays_0_0_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[14]
  PIN data_arrays_0_0_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[15]
  PIN data_arrays_0_0_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[16]
  PIN data_arrays_0_0_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[17]
  PIN data_arrays_0_0_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[18]
  PIN data_arrays_0_0_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[19]
  PIN data_arrays_0_0_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[1]
  PIN data_arrays_0_0_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[20]
  PIN data_arrays_0_0_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[21]
  PIN data_arrays_0_0_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[22]
  PIN data_arrays_0_0_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[23]
  PIN data_arrays_0_0_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[24]
  PIN data_arrays_0_0_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[25]
  PIN data_arrays_0_0_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[26]
  PIN data_arrays_0_0_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[27]
  PIN data_arrays_0_0_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[28]
  PIN data_arrays_0_0_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[29]
  PIN data_arrays_0_0_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[2]
  PIN data_arrays_0_0_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[30]
  PIN data_arrays_0_0_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[31]
  PIN data_arrays_0_0_ext_ram_rdata0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[32]
  PIN data_arrays_0_0_ext_ram_rdata0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[33]
  PIN data_arrays_0_0_ext_ram_rdata0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[34]
  PIN data_arrays_0_0_ext_ram_rdata0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[35]
  PIN data_arrays_0_0_ext_ram_rdata0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[36]
  PIN data_arrays_0_0_ext_ram_rdata0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[37]
  PIN data_arrays_0_0_ext_ram_rdata0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[38]
  PIN data_arrays_0_0_ext_ram_rdata0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[39]
  PIN data_arrays_0_0_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[3]
  PIN data_arrays_0_0_ext_ram_rdata0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[40]
  PIN data_arrays_0_0_ext_ram_rdata0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[41]
  PIN data_arrays_0_0_ext_ram_rdata0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[42]
  PIN data_arrays_0_0_ext_ram_rdata0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[43]
  PIN data_arrays_0_0_ext_ram_rdata0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[44]
  PIN data_arrays_0_0_ext_ram_rdata0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[45]
  PIN data_arrays_0_0_ext_ram_rdata0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[46]
  PIN data_arrays_0_0_ext_ram_rdata0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[47]
  PIN data_arrays_0_0_ext_ram_rdata0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[48]
  PIN data_arrays_0_0_ext_ram_rdata0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[49]
  PIN data_arrays_0_0_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[4]
  PIN data_arrays_0_0_ext_ram_rdata0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[50]
  PIN data_arrays_0_0_ext_ram_rdata0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[51]
  PIN data_arrays_0_0_ext_ram_rdata0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[52]
  PIN data_arrays_0_0_ext_ram_rdata0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[53]
  PIN data_arrays_0_0_ext_ram_rdata0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[54]
  PIN data_arrays_0_0_ext_ram_rdata0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[55]
  PIN data_arrays_0_0_ext_ram_rdata0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[56]
  PIN data_arrays_0_0_ext_ram_rdata0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[57]
  PIN data_arrays_0_0_ext_ram_rdata0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[58]
  PIN data_arrays_0_0_ext_ram_rdata0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[59]
  PIN data_arrays_0_0_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[5]
  PIN data_arrays_0_0_ext_ram_rdata0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[60]
  PIN data_arrays_0_0_ext_ram_rdata0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[61]
  PIN data_arrays_0_0_ext_ram_rdata0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[62]
  PIN data_arrays_0_0_ext_ram_rdata0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[63]
  PIN data_arrays_0_0_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[6]
  PIN data_arrays_0_0_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[7]
  PIN data_arrays_0_0_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[8]
  PIN data_arrays_0_0_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[9]
  PIN data_arrays_0_0_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[0]
  PIN data_arrays_0_0_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[10]
  PIN data_arrays_0_0_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[11]
  PIN data_arrays_0_0_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[12]
  PIN data_arrays_0_0_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[13]
  PIN data_arrays_0_0_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[14]
  PIN data_arrays_0_0_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[15]
  PIN data_arrays_0_0_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[16]
  PIN data_arrays_0_0_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[17]
  PIN data_arrays_0_0_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[18]
  PIN data_arrays_0_0_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[19]
  PIN data_arrays_0_0_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[1]
  PIN data_arrays_0_0_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[20]
  PIN data_arrays_0_0_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[21]
  PIN data_arrays_0_0_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[22]
  PIN data_arrays_0_0_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[23]
  PIN data_arrays_0_0_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[24]
  PIN data_arrays_0_0_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[25]
  PIN data_arrays_0_0_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[26]
  PIN data_arrays_0_0_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[27]
  PIN data_arrays_0_0_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[28]
  PIN data_arrays_0_0_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[29]
  PIN data_arrays_0_0_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[2]
  PIN data_arrays_0_0_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[30]
  PIN data_arrays_0_0_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[31]
  PIN data_arrays_0_0_ext_ram_rdata1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[32]
  PIN data_arrays_0_0_ext_ram_rdata1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[33]
  PIN data_arrays_0_0_ext_ram_rdata1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[34]
  PIN data_arrays_0_0_ext_ram_rdata1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[35]
  PIN data_arrays_0_0_ext_ram_rdata1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[36]
  PIN data_arrays_0_0_ext_ram_rdata1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[37]
  PIN data_arrays_0_0_ext_ram_rdata1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[38]
  PIN data_arrays_0_0_ext_ram_rdata1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[39]
  PIN data_arrays_0_0_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[3]
  PIN data_arrays_0_0_ext_ram_rdata1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[40]
  PIN data_arrays_0_0_ext_ram_rdata1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[41]
  PIN data_arrays_0_0_ext_ram_rdata1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[42]
  PIN data_arrays_0_0_ext_ram_rdata1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[43]
  PIN data_arrays_0_0_ext_ram_rdata1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[44]
  PIN data_arrays_0_0_ext_ram_rdata1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[45]
  PIN data_arrays_0_0_ext_ram_rdata1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[46]
  PIN data_arrays_0_0_ext_ram_rdata1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[47]
  PIN data_arrays_0_0_ext_ram_rdata1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[48]
  PIN data_arrays_0_0_ext_ram_rdata1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[49]
  PIN data_arrays_0_0_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[4]
  PIN data_arrays_0_0_ext_ram_rdata1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[50]
  PIN data_arrays_0_0_ext_ram_rdata1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[51]
  PIN data_arrays_0_0_ext_ram_rdata1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[52]
  PIN data_arrays_0_0_ext_ram_rdata1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[53]
  PIN data_arrays_0_0_ext_ram_rdata1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 4.000 417.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[54]
  PIN data_arrays_0_0_ext_ram_rdata1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[55]
  PIN data_arrays_0_0_ext_ram_rdata1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[56]
  PIN data_arrays_0_0_ext_ram_rdata1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[57]
  PIN data_arrays_0_0_ext_ram_rdata1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[58]
  PIN data_arrays_0_0_ext_ram_rdata1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[59]
  PIN data_arrays_0_0_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[5]
  PIN data_arrays_0_0_ext_ram_rdata1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[60]
  PIN data_arrays_0_0_ext_ram_rdata1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[61]
  PIN data_arrays_0_0_ext_ram_rdata1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[62]
  PIN data_arrays_0_0_ext_ram_rdata1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.160 4.000 448.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[63]
  PIN data_arrays_0_0_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[6]
  PIN data_arrays_0_0_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[7]
  PIN data_arrays_0_0_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[8]
  PIN data_arrays_0_0_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[9]
  PIN data_arrays_0_0_ext_ram_rdata2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[0]
  PIN data_arrays_0_0_ext_ram_rdata2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[10]
  PIN data_arrays_0_0_ext_ram_rdata2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.760 4.000 836.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[11]
  PIN data_arrays_0_0_ext_ram_rdata2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[12]
  PIN data_arrays_0_0_ext_ram_rdata2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 842.560 4.000 843.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[13]
  PIN data_arrays_0_0_ext_ram_rdata2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.960 4.000 846.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[14]
  PIN data_arrays_0_0_ext_ram_rdata2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 849.360 4.000 849.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[15]
  PIN data_arrays_0_0_ext_ram_rdata2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[16]
  PIN data_arrays_0_0_ext_ram_rdata2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[17]
  PIN data_arrays_0_0_ext_ram_rdata2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[18]
  PIN data_arrays_0_0_ext_ram_rdata2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[19]
  PIN data_arrays_0_0_ext_ram_rdata2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 800.400 4.000 801.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[1]
  PIN data_arrays_0_0_ext_ram_rdata2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[20]
  PIN data_arrays_0_0_ext_ram_rdata2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.120 4.000 871.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[21]
  PIN data_arrays_0_0_ext_ram_rdata2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 874.520 4.000 875.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[22]
  PIN data_arrays_0_0_ext_ram_rdata2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.920 4.000 878.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[23]
  PIN data_arrays_0_0_ext_ram_rdata2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[24]
  PIN data_arrays_0_0_ext_ram_rdata2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.720 4.000 885.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[25]
  PIN data_arrays_0_0_ext_ram_rdata2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[26]
  PIN data_arrays_0_0_ext_ram_rdata2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[27]
  PIN data_arrays_0_0_ext_ram_rdata2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 895.600 4.000 896.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[28]
  PIN data_arrays_0_0_ext_ram_rdata2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[29]
  PIN data_arrays_0_0_ext_ram_rdata2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.800 4.000 804.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[2]
  PIN data_arrays_0_0_ext_ram_rdata2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 902.400 4.000 903.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[30]
  PIN data_arrays_0_0_ext_ram_rdata2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[31]
  PIN data_arrays_0_0_ext_ram_rdata2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.200 4.000 909.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[32]
  PIN data_arrays_0_0_ext_ram_rdata2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.280 4.000 913.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[33]
  PIN data_arrays_0_0_ext_ram_rdata2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[34]
  PIN data_arrays_0_0_ext_ram_rdata2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[35]
  PIN data_arrays_0_0_ext_ram_rdata2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 923.480 4.000 924.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[36]
  PIN data_arrays_0_0_ext_ram_rdata2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.880 4.000 927.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[37]
  PIN data_arrays_0_0_ext_ram_rdata2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[38]
  PIN data_arrays_0_0_ext_ram_rdata2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 4.000 934.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[39]
  PIN data_arrays_0_0_ext_ram_rdata2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.200 4.000 807.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[3]
  PIN data_arrays_0_0_ext_ram_rdata2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.760 4.000 938.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[40]
  PIN data_arrays_0_0_ext_ram_rdata2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[41]
  PIN data_arrays_0_0_ext_ram_rdata2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 944.560 4.000 945.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[42]
  PIN data_arrays_0_0_ext_ram_rdata2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[43]
  PIN data_arrays_0_0_ext_ram_rdata2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[44]
  PIN data_arrays_0_0_ext_ram_rdata2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[45]
  PIN data_arrays_0_0_ext_ram_rdata2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[46]
  PIN data_arrays_0_0_ext_ram_rdata2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[47]
  PIN data_arrays_0_0_ext_ram_rdata2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[48]
  PIN data_arrays_0_0_ext_ram_rdata2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.720 4.000 970.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[49]
  PIN data_arrays_0_0_ext_ram_rdata2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[4]
  PIN data_arrays_0_0_ext_ram_rdata2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.120 4.000 973.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[50]
  PIN data_arrays_0_0_ext_ram_rdata2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 976.520 4.000 977.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[51]
  PIN data_arrays_0_0_ext_ram_rdata2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.920 4.000 980.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[52]
  PIN data_arrays_0_0_ext_ram_rdata2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[53]
  PIN data_arrays_0_0_ext_ram_rdata2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.720 4.000 987.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[54]
  PIN data_arrays_0_0_ext_ram_rdata2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.800 4.000 991.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[55]
  PIN data_arrays_0_0_ext_ram_rdata2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[56]
  PIN data_arrays_0_0_ext_ram_rdata2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 997.600 4.000 998.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[57]
  PIN data_arrays_0_0_ext_ram_rdata2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.000 4.000 1001.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[58]
  PIN data_arrays_0_0_ext_ram_rdata2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1004.400 4.000 1005.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[59]
  PIN data_arrays_0_0_ext_ram_rdata2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[5]
  PIN data_arrays_0_0_ext_ram_rdata2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[60]
  PIN data_arrays_0_0_ext_ram_rdata2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[61]
  PIN data_arrays_0_0_ext_ram_rdata2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1015.280 4.000 1015.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[62]
  PIN data_arrays_0_0_ext_ram_rdata2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.680 4.000 1019.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[63]
  PIN data_arrays_0_0_ext_ram_rdata2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[6]
  PIN data_arrays_0_0_ext_ram_rdata2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 821.480 4.000 822.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[7]
  PIN data_arrays_0_0_ext_ram_rdata2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.880 4.000 825.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[8]
  PIN data_arrays_0_0_ext_ram_rdata2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[9]
  PIN data_arrays_0_0_ext_ram_rdata3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1022.080 4.000 1022.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[0]
  PIN data_arrays_0_0_ext_ram_rdata3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[10]
  PIN data_arrays_0_0_ext_ram_rdata3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[11]
  PIN data_arrays_0_0_ext_ram_rdata3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[12]
  PIN data_arrays_0_0_ext_ram_rdata3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1068.320 4.000 1068.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[13]
  PIN data_arrays_0_0_ext_ram_rdata3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.720 4.000 1072.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[14]
  PIN data_arrays_0_0_ext_ram_rdata3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.120 4.000 1075.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[15]
  PIN data_arrays_0_0_ext_ram_rdata3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1078.520 4.000 1079.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[16]
  PIN data_arrays_0_0_ext_ram_rdata3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.920 4.000 1082.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[17]
  PIN data_arrays_0_0_ext_ram_rdata3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1085.320 4.000 1085.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[18]
  PIN data_arrays_0_0_ext_ram_rdata3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1089.400 4.000 1090.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[19]
  PIN data_arrays_0_0_ext_ram_rdata3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[1]
  PIN data_arrays_0_0_ext_ram_rdata3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1092.800 4.000 1093.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[20]
  PIN data_arrays_0_0_ext_ram_rdata3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.200 4.000 1096.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[21]
  PIN data_arrays_0_0_ext_ram_rdata3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[22]
  PIN data_arrays_0_0_ext_ram_rdata3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1103.000 4.000 1103.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[23]
  PIN data_arrays_0_0_ext_ram_rdata3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1106.400 4.000 1107.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[24]
  PIN data_arrays_0_0_ext_ram_rdata3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1110.480 4.000 1111.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[25]
  PIN data_arrays_0_0_ext_ram_rdata3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1113.880 4.000 1114.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[26]
  PIN data_arrays_0_0_ext_ram_rdata3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.280 4.000 1117.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[27]
  PIN data_arrays_0_0_ext_ram_rdata3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.680 4.000 1121.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[28]
  PIN data_arrays_0_0_ext_ram_rdata3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.080 4.000 1124.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[29]
  PIN data_arrays_0_0_ext_ram_rdata3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[2]
  PIN data_arrays_0_0_ext_ram_rdata3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.160 4.000 1128.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[30]
  PIN data_arrays_0_0_ext_ram_rdata3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1131.560 4.000 1132.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[31]
  PIN data_arrays_0_0_ext_ram_rdata3[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1134.960 4.000 1135.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[32]
  PIN data_arrays_0_0_ext_ram_rdata3[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1138.360 4.000 1138.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[33]
  PIN data_arrays_0_0_ext_ram_rdata3[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.760 4.000 1142.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[34]
  PIN data_arrays_0_0_ext_ram_rdata3[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.160 4.000 1145.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[35]
  PIN data_arrays_0_0_ext_ram_rdata3[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[36]
  PIN data_arrays_0_0_ext_ram_rdata3[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[37]
  PIN data_arrays_0_0_ext_ram_rdata3[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[38]
  PIN data_arrays_0_0_ext_ram_rdata3[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[39]
  PIN data_arrays_0_0_ext_ram_rdata3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.960 4.000 1033.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[3]
  PIN data_arrays_0_0_ext_ram_rdata3[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[40]
  PIN data_arrays_0_0_ext_ram_rdata3[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[41]
  PIN data_arrays_0_0_ext_ram_rdata3[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1170.320 4.000 1170.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[42]
  PIN data_arrays_0_0_ext_ram_rdata3[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.720 4.000 1174.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[43]
  PIN data_arrays_0_0_ext_ram_rdata3[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.120 4.000 1177.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[44]
  PIN data_arrays_0_0_ext_ram_rdata3[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1180.520 4.000 1181.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[45]
  PIN data_arrays_0_0_ext_ram_rdata3[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.920 4.000 1184.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[46]
  PIN data_arrays_0_0_ext_ram_rdata3[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1188.000 4.000 1188.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[47]
  PIN data_arrays_0_0_ext_ram_rdata3[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1191.400 4.000 1192.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[48]
  PIN data_arrays_0_0_ext_ram_rdata3[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.800 4.000 1195.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[49]
  PIN data_arrays_0_0_ext_ram_rdata3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[4]
  PIN data_arrays_0_0_ext_ram_rdata3[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1198.200 4.000 1198.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[50]
  PIN data_arrays_0_0_ext_ram_rdata3[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1201.600 4.000 1202.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[51]
  PIN data_arrays_0_0_ext_ram_rdata3[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1205.000 4.000 1205.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[52]
  PIN data_arrays_0_0_ext_ram_rdata3[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1209.080 4.000 1209.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[53]
  PIN data_arrays_0_0_ext_ram_rdata3[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1212.480 4.000 1213.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[54]
  PIN data_arrays_0_0_ext_ram_rdata3[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1215.880 4.000 1216.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[55]
  PIN data_arrays_0_0_ext_ram_rdata3[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1219.280 4.000 1219.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[56]
  PIN data_arrays_0_0_ext_ram_rdata3[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1222.680 4.000 1223.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[57]
  PIN data_arrays_0_0_ext_ram_rdata3[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1226.760 4.000 1227.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[58]
  PIN data_arrays_0_0_ext_ram_rdata3[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.160 4.000 1230.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[59]
  PIN data_arrays_0_0_ext_ram_rdata3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1039.760 4.000 1040.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[5]
  PIN data_arrays_0_0_ext_ram_rdata3[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1233.560 4.000 1234.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[60]
  PIN data_arrays_0_0_ext_ram_rdata3[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.960 4.000 1237.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[61]
  PIN data_arrays_0_0_ext_ram_rdata3[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1240.360 4.000 1240.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[62]
  PIN data_arrays_0_0_ext_ram_rdata3[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.760 4.000 1244.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[63]
  PIN data_arrays_0_0_ext_ram_rdata3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.160 4.000 1043.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[6]
  PIN data_arrays_0_0_ext_ram_rdata3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1046.560 4.000 1047.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[7]
  PIN data_arrays_0_0_ext_ram_rdata3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[8]
  PIN data_arrays_0_0_ext_ram_rdata3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[9]
  PIN data_arrays_0_0_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[0]
  PIN data_arrays_0_0_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata[10]
  PIN data_arrays_0_0_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata[11]
  PIN data_arrays_0_0_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[12]
  PIN data_arrays_0_0_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 532.480 4.000 533.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[13]
  PIN data_arrays_0_0_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[14]
  PIN data_arrays_0_0_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata[15]
  PIN data_arrays_0_0_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata[16]
  PIN data_arrays_0_0_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata[17]
  PIN data_arrays_0_0_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[18]
  PIN data_arrays_0_0_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[19]
  PIN data_arrays_0_0_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 490.320 4.000 490.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[1]
  PIN data_arrays_0_0_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[20]
  PIN data_arrays_0_0_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata[21]
  PIN data_arrays_0_0_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata[22]
  PIN data_arrays_0_0_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata[23]
  PIN data_arrays_0_0_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata[24]
  PIN data_arrays_0_0_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[25]
  PIN data_arrays_0_0_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[26]
  PIN data_arrays_0_0_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata[27]
  PIN data_arrays_0_0_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[28]
  PIN data_arrays_0_0_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[29]
  PIN data_arrays_0_0_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[2]
  PIN data_arrays_0_0_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[30]
  PIN data_arrays_0_0_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[31]
  PIN data_arrays_0_0_ext_ram_wdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[32]
  PIN data_arrays_0_0_ext_ram_wdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[33]
  PIN data_arrays_0_0_ext_ram_wdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[34]
  PIN data_arrays_0_0_ext_ram_wdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.000 4.000 610.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[35]
  PIN data_arrays_0_0_ext_ram_wdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.080 4.000 614.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[36]
  PIN data_arrays_0_0_ext_ram_wdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[37]
  PIN data_arrays_0_0_ext_ram_wdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.880 4.000 621.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[38]
  PIN data_arrays_0_0_ext_ram_wdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata[39]
  PIN data_arrays_0_0_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[3]
  PIN data_arrays_0_0_ext_ram_wdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata[40]
  PIN data_arrays_0_0_ext_ram_wdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[41]
  PIN data_arrays_0_0_ext_ram_wdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[42]
  PIN data_arrays_0_0_ext_ram_wdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[43]
  PIN data_arrays_0_0_ext_ram_wdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata[44]
  PIN data_arrays_0_0_ext_ram_wdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 645.360 4.000 645.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata[45]
  PIN data_arrays_0_0_ext_ram_wdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata[46]
  PIN data_arrays_0_0_ext_ram_wdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[47]
  PIN data_arrays_0_0_ext_ram_wdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata[48]
  PIN data_arrays_0_0_ext_ram_wdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[49]
  PIN data_arrays_0_0_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[4]
  PIN data_arrays_0_0_ext_ram_wdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata[50]
  PIN data_arrays_0_0_ext_ram_wdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata[51]
  PIN data_arrays_0_0_ext_ram_wdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata[52]
  PIN data_arrays_0_0_ext_ram_wdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[53]
  PIN data_arrays_0_0_ext_ram_wdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[54]
  PIN data_arrays_0_0_ext_ram_wdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[55]
  PIN data_arrays_0_0_ext_ram_wdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata[56]
  PIN data_arrays_0_0_ext_ram_wdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.520 4.000 688.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[57]
  PIN data_arrays_0_0_ext_ram_wdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[58]
  PIN data_arrays_0_0_ext_ram_wdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[59]
  PIN data_arrays_0_0_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[5]
  PIN data_arrays_0_0_ext_ram_wdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 698.400 4.000 699.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[60]
  PIN data_arrays_0_0_ext_ram_wdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[61]
  PIN data_arrays_0_0_ext_ram_wdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 4.000 705.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[62]
  PIN data_arrays_0_0_ext_ram_wdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[63]
  PIN data_arrays_0_0_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[6]
  PIN data_arrays_0_0_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[7]
  PIN data_arrays_0_0_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[8]
  PIN data_arrays_0_0_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[9]
  PIN data_arrays_0_0_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.760 4.000 734.360 ;
    END
  END data_arrays_0_0_ext_ram_web
  PIN data_arrays_0_0_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END data_arrays_0_0_ext_ram_wmask[0]
  PIN data_arrays_0_0_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END data_arrays_0_0_ext_ram_wmask[1]
  PIN data_arrays_0_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1037.040 1767.600 1037.640 ;
    END
  END data_arrays_0_ext_ram_addr1[0]
  PIN data_arrays_0_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1042.480 1767.600 1043.080 ;
    END
  END data_arrays_0_ext_ram_addr1[1]
  PIN data_arrays_0_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1047.920 1767.600 1048.520 ;
    END
  END data_arrays_0_ext_ram_addr1[2]
  PIN data_arrays_0_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1053.360 1767.600 1053.960 ;
    END
  END data_arrays_0_ext_ram_addr1[3]
  PIN data_arrays_0_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1058.800 1767.600 1059.400 ;
    END
  END data_arrays_0_ext_ram_addr1[4]
  PIN data_arrays_0_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1064.240 1767.600 1064.840 ;
    END
  END data_arrays_0_ext_ram_addr1[5]
  PIN data_arrays_0_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1069.680 1767.600 1070.280 ;
    END
  END data_arrays_0_ext_ram_addr1[6]
  PIN data_arrays_0_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1075.120 1767.600 1075.720 ;
    END
  END data_arrays_0_ext_ram_addr1[7]
  PIN data_arrays_0_ext_ram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1080.560 1767.600 1081.160 ;
    END
  END data_arrays_0_ext_ram_addr1[8]
  PIN data_arrays_0_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 695.680 1767.600 696.280 ;
    END
  END data_arrays_0_ext_ram_addr[0]
  PIN data_arrays_0_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 701.120 1767.600 701.720 ;
    END
  END data_arrays_0_ext_ram_addr[1]
  PIN data_arrays_0_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 706.560 1767.600 707.160 ;
    END
  END data_arrays_0_ext_ram_addr[2]
  PIN data_arrays_0_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 712.000 1767.600 712.600 ;
    END
  END data_arrays_0_ext_ram_addr[3]
  PIN data_arrays_0_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 717.440 1767.600 718.040 ;
    END
  END data_arrays_0_ext_ram_addr[4]
  PIN data_arrays_0_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 722.880 1767.600 723.480 ;
    END
  END data_arrays_0_ext_ram_addr[5]
  PIN data_arrays_0_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 728.320 1767.600 728.920 ;
    END
  END data_arrays_0_ext_ram_addr[6]
  PIN data_arrays_0_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 733.760 1767.600 734.360 ;
    END
  END data_arrays_0_ext_ram_addr[7]
  PIN data_arrays_0_ext_ram_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 739.200 1767.600 739.800 ;
    END
  END data_arrays_0_ext_ram_addr[8]
  PIN data_arrays_0_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 744.640 1767.600 745.240 ;
    END
  END data_arrays_0_ext_ram_clk
  PIN data_arrays_0_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 993.520 1767.600 994.120 ;
    END
  END data_arrays_0_ext_ram_csb1[0]
  PIN data_arrays_0_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 998.960 1767.600 999.560 ;
    END
  END data_arrays_0_ext_ram_csb1[1]
  PIN data_arrays_0_ext_ram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1004.400 1767.600 1005.000 ;
    END
  END data_arrays_0_ext_ram_csb1[2]
  PIN data_arrays_0_ext_ram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1009.840 1767.600 1010.440 ;
    END
  END data_arrays_0_ext_ram_csb1[3]
  PIN data_arrays_0_ext_ram_csb1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1015.280 1767.600 1015.880 ;
    END
  END data_arrays_0_ext_ram_csb1[4]
  PIN data_arrays_0_ext_ram_csb1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1020.720 1767.600 1021.320 ;
    END
  END data_arrays_0_ext_ram_csb1[5]
  PIN data_arrays_0_ext_ram_csb1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1026.160 1767.600 1026.760 ;
    END
  END data_arrays_0_ext_ram_csb1[6]
  PIN data_arrays_0_ext_ram_csb1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1031.600 1767.600 1032.200 ;
    END
  END data_arrays_0_ext_ram_csb1[7]
  PIN data_arrays_0_ext_ram_csb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 945.240 1767.600 945.840 ;
    END
  END data_arrays_0_ext_ram_csb[0]
  PIN data_arrays_0_ext_ram_csb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 950.680 1767.600 951.280 ;
    END
  END data_arrays_0_ext_ram_csb[1]
  PIN data_arrays_0_ext_ram_csb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 956.120 1767.600 956.720 ;
    END
  END data_arrays_0_ext_ram_csb[2]
  PIN data_arrays_0_ext_ram_csb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 961.560 1767.600 962.160 ;
    END
  END data_arrays_0_ext_ram_csb[3]
  PIN data_arrays_0_ext_ram_csb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 967.000 1767.600 967.600 ;
    END
  END data_arrays_0_ext_ram_csb[4]
  PIN data_arrays_0_ext_ram_csb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 972.440 1767.600 973.040 ;
    END
  END data_arrays_0_ext_ram_csb[5]
  PIN data_arrays_0_ext_ram_csb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 977.880 1767.600 978.480 ;
    END
  END data_arrays_0_ext_ram_csb[6]
  PIN data_arrays_0_ext_ram_csb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 983.320 1767.600 983.920 ;
    END
  END data_arrays_0_ext_ram_csb[7]
  PIN data_arrays_0_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 2.080 1767.600 2.680 ;
    END
  END data_arrays_0_ext_ram_rdata0[0]
  PIN data_arrays_0_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 55.800 1767.600 56.400 ;
    END
  END data_arrays_0_ext_ram_rdata0[10]
  PIN data_arrays_0_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 61.240 1767.600 61.840 ;
    END
  END data_arrays_0_ext_ram_rdata0[11]
  PIN data_arrays_0_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 66.680 1767.600 67.280 ;
    END
  END data_arrays_0_ext_ram_rdata0[12]
  PIN data_arrays_0_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 72.120 1767.600 72.720 ;
    END
  END data_arrays_0_ext_ram_rdata0[13]
  PIN data_arrays_0_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 77.560 1767.600 78.160 ;
    END
  END data_arrays_0_ext_ram_rdata0[14]
  PIN data_arrays_0_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 83.000 1767.600 83.600 ;
    END
  END data_arrays_0_ext_ram_rdata0[15]
  PIN data_arrays_0_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 88.440 1767.600 89.040 ;
    END
  END data_arrays_0_ext_ram_rdata0[16]
  PIN data_arrays_0_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 93.880 1767.600 94.480 ;
    END
  END data_arrays_0_ext_ram_rdata0[17]
  PIN data_arrays_0_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 99.320 1767.600 99.920 ;
    END
  END data_arrays_0_ext_ram_rdata0[18]
  PIN data_arrays_0_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 104.760 1767.600 105.360 ;
    END
  END data_arrays_0_ext_ram_rdata0[19]
  PIN data_arrays_0_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 6.840 1767.600 7.440 ;
    END
  END data_arrays_0_ext_ram_rdata0[1]
  PIN data_arrays_0_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 110.200 1767.600 110.800 ;
    END
  END data_arrays_0_ext_ram_rdata0[20]
  PIN data_arrays_0_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 115.640 1767.600 116.240 ;
    END
  END data_arrays_0_ext_ram_rdata0[21]
  PIN data_arrays_0_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 121.080 1767.600 121.680 ;
    END
  END data_arrays_0_ext_ram_rdata0[22]
  PIN data_arrays_0_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 126.520 1767.600 127.120 ;
    END
  END data_arrays_0_ext_ram_rdata0[23]
  PIN data_arrays_0_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 131.960 1767.600 132.560 ;
    END
  END data_arrays_0_ext_ram_rdata0[24]
  PIN data_arrays_0_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 137.400 1767.600 138.000 ;
    END
  END data_arrays_0_ext_ram_rdata0[25]
  PIN data_arrays_0_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 142.840 1767.600 143.440 ;
    END
  END data_arrays_0_ext_ram_rdata0[26]
  PIN data_arrays_0_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 148.280 1767.600 148.880 ;
    END
  END data_arrays_0_ext_ram_rdata0[27]
  PIN data_arrays_0_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 153.720 1767.600 154.320 ;
    END
  END data_arrays_0_ext_ram_rdata0[28]
  PIN data_arrays_0_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 159.160 1767.600 159.760 ;
    END
  END data_arrays_0_ext_ram_rdata0[29]
  PIN data_arrays_0_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 12.280 1767.600 12.880 ;
    END
  END data_arrays_0_ext_ram_rdata0[2]
  PIN data_arrays_0_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 164.600 1767.600 165.200 ;
    END
  END data_arrays_0_ext_ram_rdata0[30]
  PIN data_arrays_0_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 170.040 1767.600 170.640 ;
    END
  END data_arrays_0_ext_ram_rdata0[31]
  PIN data_arrays_0_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 17.720 1767.600 18.320 ;
    END
  END data_arrays_0_ext_ram_rdata0[3]
  PIN data_arrays_0_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 23.160 1767.600 23.760 ;
    END
  END data_arrays_0_ext_ram_rdata0[4]
  PIN data_arrays_0_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 28.600 1767.600 29.200 ;
    END
  END data_arrays_0_ext_ram_rdata0[5]
  PIN data_arrays_0_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 34.040 1767.600 34.640 ;
    END
  END data_arrays_0_ext_ram_rdata0[6]
  PIN data_arrays_0_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 39.480 1767.600 40.080 ;
    END
  END data_arrays_0_ext_ram_rdata0[7]
  PIN data_arrays_0_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 44.920 1767.600 45.520 ;
    END
  END data_arrays_0_ext_ram_rdata0[8]
  PIN data_arrays_0_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 50.360 1767.600 50.960 ;
    END
  END data_arrays_0_ext_ram_rdata0[9]
  PIN data_arrays_0_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 175.480 1767.600 176.080 ;
    END
  END data_arrays_0_ext_ram_rdata1[0]
  PIN data_arrays_0_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 229.200 1767.600 229.800 ;
    END
  END data_arrays_0_ext_ram_rdata1[10]
  PIN data_arrays_0_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 234.640 1767.600 235.240 ;
    END
  END data_arrays_0_ext_ram_rdata1[11]
  PIN data_arrays_0_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 240.080 1767.600 240.680 ;
    END
  END data_arrays_0_ext_ram_rdata1[12]
  PIN data_arrays_0_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 245.520 1767.600 246.120 ;
    END
  END data_arrays_0_ext_ram_rdata1[13]
  PIN data_arrays_0_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 250.960 1767.600 251.560 ;
    END
  END data_arrays_0_ext_ram_rdata1[14]
  PIN data_arrays_0_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 256.400 1767.600 257.000 ;
    END
  END data_arrays_0_ext_ram_rdata1[15]
  PIN data_arrays_0_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 261.840 1767.600 262.440 ;
    END
  END data_arrays_0_ext_ram_rdata1[16]
  PIN data_arrays_0_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 267.280 1767.600 267.880 ;
    END
  END data_arrays_0_ext_ram_rdata1[17]
  PIN data_arrays_0_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 272.720 1767.600 273.320 ;
    END
  END data_arrays_0_ext_ram_rdata1[18]
  PIN data_arrays_0_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 278.160 1767.600 278.760 ;
    END
  END data_arrays_0_ext_ram_rdata1[19]
  PIN data_arrays_0_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 180.920 1767.600 181.520 ;
    END
  END data_arrays_0_ext_ram_rdata1[1]
  PIN data_arrays_0_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 283.600 1767.600 284.200 ;
    END
  END data_arrays_0_ext_ram_rdata1[20]
  PIN data_arrays_0_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 289.040 1767.600 289.640 ;
    END
  END data_arrays_0_ext_ram_rdata1[21]
  PIN data_arrays_0_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 294.480 1767.600 295.080 ;
    END
  END data_arrays_0_ext_ram_rdata1[22]
  PIN data_arrays_0_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 299.920 1767.600 300.520 ;
    END
  END data_arrays_0_ext_ram_rdata1[23]
  PIN data_arrays_0_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 305.360 1767.600 305.960 ;
    END
  END data_arrays_0_ext_ram_rdata1[24]
  PIN data_arrays_0_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 310.800 1767.600 311.400 ;
    END
  END data_arrays_0_ext_ram_rdata1[25]
  PIN data_arrays_0_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 316.240 1767.600 316.840 ;
    END
  END data_arrays_0_ext_ram_rdata1[26]
  PIN data_arrays_0_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 321.680 1767.600 322.280 ;
    END
  END data_arrays_0_ext_ram_rdata1[27]
  PIN data_arrays_0_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 327.120 1767.600 327.720 ;
    END
  END data_arrays_0_ext_ram_rdata1[28]
  PIN data_arrays_0_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 332.560 1767.600 333.160 ;
    END
  END data_arrays_0_ext_ram_rdata1[29]
  PIN data_arrays_0_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 186.360 1767.600 186.960 ;
    END
  END data_arrays_0_ext_ram_rdata1[2]
  PIN data_arrays_0_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 338.000 1767.600 338.600 ;
    END
  END data_arrays_0_ext_ram_rdata1[30]
  PIN data_arrays_0_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 343.440 1767.600 344.040 ;
    END
  END data_arrays_0_ext_ram_rdata1[31]
  PIN data_arrays_0_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 191.800 1767.600 192.400 ;
    END
  END data_arrays_0_ext_ram_rdata1[3]
  PIN data_arrays_0_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 197.240 1767.600 197.840 ;
    END
  END data_arrays_0_ext_ram_rdata1[4]
  PIN data_arrays_0_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 202.000 1767.600 202.600 ;
    END
  END data_arrays_0_ext_ram_rdata1[5]
  PIN data_arrays_0_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 207.440 1767.600 208.040 ;
    END
  END data_arrays_0_ext_ram_rdata1[6]
  PIN data_arrays_0_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 212.880 1767.600 213.480 ;
    END
  END data_arrays_0_ext_ram_rdata1[7]
  PIN data_arrays_0_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 218.320 1767.600 218.920 ;
    END
  END data_arrays_0_ext_ram_rdata1[8]
  PIN data_arrays_0_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 223.760 1767.600 224.360 ;
    END
  END data_arrays_0_ext_ram_rdata1[9]
  PIN data_arrays_0_ext_ram_rdata2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 348.880 1767.600 349.480 ;
    END
  END data_arrays_0_ext_ram_rdata2[0]
  PIN data_arrays_0_ext_ram_rdata2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 402.600 1767.600 403.200 ;
    END
  END data_arrays_0_ext_ram_rdata2[10]
  PIN data_arrays_0_ext_ram_rdata2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 408.040 1767.600 408.640 ;
    END
  END data_arrays_0_ext_ram_rdata2[11]
  PIN data_arrays_0_ext_ram_rdata2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 413.480 1767.600 414.080 ;
    END
  END data_arrays_0_ext_ram_rdata2[12]
  PIN data_arrays_0_ext_ram_rdata2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 418.920 1767.600 419.520 ;
    END
  END data_arrays_0_ext_ram_rdata2[13]
  PIN data_arrays_0_ext_ram_rdata2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 424.360 1767.600 424.960 ;
    END
  END data_arrays_0_ext_ram_rdata2[14]
  PIN data_arrays_0_ext_ram_rdata2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 429.800 1767.600 430.400 ;
    END
  END data_arrays_0_ext_ram_rdata2[15]
  PIN data_arrays_0_ext_ram_rdata2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 435.240 1767.600 435.840 ;
    END
  END data_arrays_0_ext_ram_rdata2[16]
  PIN data_arrays_0_ext_ram_rdata2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 440.680 1767.600 441.280 ;
    END
  END data_arrays_0_ext_ram_rdata2[17]
  PIN data_arrays_0_ext_ram_rdata2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 446.120 1767.600 446.720 ;
    END
  END data_arrays_0_ext_ram_rdata2[18]
  PIN data_arrays_0_ext_ram_rdata2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 451.560 1767.600 452.160 ;
    END
  END data_arrays_0_ext_ram_rdata2[19]
  PIN data_arrays_0_ext_ram_rdata2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 354.320 1767.600 354.920 ;
    END
  END data_arrays_0_ext_ram_rdata2[1]
  PIN data_arrays_0_ext_ram_rdata2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 457.000 1767.600 457.600 ;
    END
  END data_arrays_0_ext_ram_rdata2[20]
  PIN data_arrays_0_ext_ram_rdata2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 462.440 1767.600 463.040 ;
    END
  END data_arrays_0_ext_ram_rdata2[21]
  PIN data_arrays_0_ext_ram_rdata2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 467.880 1767.600 468.480 ;
    END
  END data_arrays_0_ext_ram_rdata2[22]
  PIN data_arrays_0_ext_ram_rdata2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 473.320 1767.600 473.920 ;
    END
  END data_arrays_0_ext_ram_rdata2[23]
  PIN data_arrays_0_ext_ram_rdata2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 478.760 1767.600 479.360 ;
    END
  END data_arrays_0_ext_ram_rdata2[24]
  PIN data_arrays_0_ext_ram_rdata2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 484.200 1767.600 484.800 ;
    END
  END data_arrays_0_ext_ram_rdata2[25]
  PIN data_arrays_0_ext_ram_rdata2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 489.640 1767.600 490.240 ;
    END
  END data_arrays_0_ext_ram_rdata2[26]
  PIN data_arrays_0_ext_ram_rdata2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 495.080 1767.600 495.680 ;
    END
  END data_arrays_0_ext_ram_rdata2[27]
  PIN data_arrays_0_ext_ram_rdata2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 500.520 1767.600 501.120 ;
    END
  END data_arrays_0_ext_ram_rdata2[28]
  PIN data_arrays_0_ext_ram_rdata2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 505.960 1767.600 506.560 ;
    END
  END data_arrays_0_ext_ram_rdata2[29]
  PIN data_arrays_0_ext_ram_rdata2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 359.760 1767.600 360.360 ;
    END
  END data_arrays_0_ext_ram_rdata2[2]
  PIN data_arrays_0_ext_ram_rdata2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 511.400 1767.600 512.000 ;
    END
  END data_arrays_0_ext_ram_rdata2[30]
  PIN data_arrays_0_ext_ram_rdata2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 516.840 1767.600 517.440 ;
    END
  END data_arrays_0_ext_ram_rdata2[31]
  PIN data_arrays_0_ext_ram_rdata2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 365.200 1767.600 365.800 ;
    END
  END data_arrays_0_ext_ram_rdata2[3]
  PIN data_arrays_0_ext_ram_rdata2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 370.640 1767.600 371.240 ;
    END
  END data_arrays_0_ext_ram_rdata2[4]
  PIN data_arrays_0_ext_ram_rdata2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 376.080 1767.600 376.680 ;
    END
  END data_arrays_0_ext_ram_rdata2[5]
  PIN data_arrays_0_ext_ram_rdata2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 381.520 1767.600 382.120 ;
    END
  END data_arrays_0_ext_ram_rdata2[6]
  PIN data_arrays_0_ext_ram_rdata2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 386.960 1767.600 387.560 ;
    END
  END data_arrays_0_ext_ram_rdata2[7]
  PIN data_arrays_0_ext_ram_rdata2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 392.400 1767.600 393.000 ;
    END
  END data_arrays_0_ext_ram_rdata2[8]
  PIN data_arrays_0_ext_ram_rdata2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 397.160 1767.600 397.760 ;
    END
  END data_arrays_0_ext_ram_rdata2[9]
  PIN data_arrays_0_ext_ram_rdata3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 522.280 1767.600 522.880 ;
    END
  END data_arrays_0_ext_ram_rdata3[0]
  PIN data_arrays_0_ext_ram_rdata3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 576.680 1767.600 577.280 ;
    END
  END data_arrays_0_ext_ram_rdata3[10]
  PIN data_arrays_0_ext_ram_rdata3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 582.120 1767.600 582.720 ;
    END
  END data_arrays_0_ext_ram_rdata3[11]
  PIN data_arrays_0_ext_ram_rdata3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 587.560 1767.600 588.160 ;
    END
  END data_arrays_0_ext_ram_rdata3[12]
  PIN data_arrays_0_ext_ram_rdata3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 593.000 1767.600 593.600 ;
    END
  END data_arrays_0_ext_ram_rdata3[13]
  PIN data_arrays_0_ext_ram_rdata3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 597.760 1767.600 598.360 ;
    END
  END data_arrays_0_ext_ram_rdata3[14]
  PIN data_arrays_0_ext_ram_rdata3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 603.200 1767.600 603.800 ;
    END
  END data_arrays_0_ext_ram_rdata3[15]
  PIN data_arrays_0_ext_ram_rdata3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 608.640 1767.600 609.240 ;
    END
  END data_arrays_0_ext_ram_rdata3[16]
  PIN data_arrays_0_ext_ram_rdata3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 614.080 1767.600 614.680 ;
    END
  END data_arrays_0_ext_ram_rdata3[17]
  PIN data_arrays_0_ext_ram_rdata3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 619.520 1767.600 620.120 ;
    END
  END data_arrays_0_ext_ram_rdata3[18]
  PIN data_arrays_0_ext_ram_rdata3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 624.960 1767.600 625.560 ;
    END
  END data_arrays_0_ext_ram_rdata3[19]
  PIN data_arrays_0_ext_ram_rdata3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 527.720 1767.600 528.320 ;
    END
  END data_arrays_0_ext_ram_rdata3[1]
  PIN data_arrays_0_ext_ram_rdata3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 630.400 1767.600 631.000 ;
    END
  END data_arrays_0_ext_ram_rdata3[20]
  PIN data_arrays_0_ext_ram_rdata3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 635.840 1767.600 636.440 ;
    END
  END data_arrays_0_ext_ram_rdata3[21]
  PIN data_arrays_0_ext_ram_rdata3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 641.280 1767.600 641.880 ;
    END
  END data_arrays_0_ext_ram_rdata3[22]
  PIN data_arrays_0_ext_ram_rdata3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 646.720 1767.600 647.320 ;
    END
  END data_arrays_0_ext_ram_rdata3[23]
  PIN data_arrays_0_ext_ram_rdata3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 652.160 1767.600 652.760 ;
    END
  END data_arrays_0_ext_ram_rdata3[24]
  PIN data_arrays_0_ext_ram_rdata3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 657.600 1767.600 658.200 ;
    END
  END data_arrays_0_ext_ram_rdata3[25]
  PIN data_arrays_0_ext_ram_rdata3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 663.040 1767.600 663.640 ;
    END
  END data_arrays_0_ext_ram_rdata3[26]
  PIN data_arrays_0_ext_ram_rdata3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 668.480 1767.600 669.080 ;
    END
  END data_arrays_0_ext_ram_rdata3[27]
  PIN data_arrays_0_ext_ram_rdata3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 673.920 1767.600 674.520 ;
    END
  END data_arrays_0_ext_ram_rdata3[28]
  PIN data_arrays_0_ext_ram_rdata3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 679.360 1767.600 679.960 ;
    END
  END data_arrays_0_ext_ram_rdata3[29]
  PIN data_arrays_0_ext_ram_rdata3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 533.160 1767.600 533.760 ;
    END
  END data_arrays_0_ext_ram_rdata3[2]
  PIN data_arrays_0_ext_ram_rdata3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 684.800 1767.600 685.400 ;
    END
  END data_arrays_0_ext_ram_rdata3[30]
  PIN data_arrays_0_ext_ram_rdata3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 690.240 1767.600 690.840 ;
    END
  END data_arrays_0_ext_ram_rdata3[31]
  PIN data_arrays_0_ext_ram_rdata3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 538.600 1767.600 539.200 ;
    END
  END data_arrays_0_ext_ram_rdata3[3]
  PIN data_arrays_0_ext_ram_rdata3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 544.040 1767.600 544.640 ;
    END
  END data_arrays_0_ext_ram_rdata3[4]
  PIN data_arrays_0_ext_ram_rdata3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 549.480 1767.600 550.080 ;
    END
  END data_arrays_0_ext_ram_rdata3[5]
  PIN data_arrays_0_ext_ram_rdata3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 554.920 1767.600 555.520 ;
    END
  END data_arrays_0_ext_ram_rdata3[6]
  PIN data_arrays_0_ext_ram_rdata3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 560.360 1767.600 560.960 ;
    END
  END data_arrays_0_ext_ram_rdata3[7]
  PIN data_arrays_0_ext_ram_rdata3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 565.800 1767.600 566.400 ;
    END
  END data_arrays_0_ext_ram_rdata3[8]
  PIN data_arrays_0_ext_ram_rdata3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 571.240 1767.600 571.840 ;
    END
  END data_arrays_0_ext_ram_rdata3[9]
  PIN data_arrays_0_ext_ram_rdata4[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1086.000 1767.600 1086.600 ;
    END
  END data_arrays_0_ext_ram_rdata4[0]
  PIN data_arrays_0_ext_ram_rdata4[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1140.400 1767.600 1141.000 ;
    END
  END data_arrays_0_ext_ram_rdata4[10]
  PIN data_arrays_0_ext_ram_rdata4[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1145.840 1767.600 1146.440 ;
    END
  END data_arrays_0_ext_ram_rdata4[11]
  PIN data_arrays_0_ext_ram_rdata4[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1151.280 1767.600 1151.880 ;
    END
  END data_arrays_0_ext_ram_rdata4[12]
  PIN data_arrays_0_ext_ram_rdata4[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1156.720 1767.600 1157.320 ;
    END
  END data_arrays_0_ext_ram_rdata4[13]
  PIN data_arrays_0_ext_ram_rdata4[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1162.160 1767.600 1162.760 ;
    END
  END data_arrays_0_ext_ram_rdata4[14]
  PIN data_arrays_0_ext_ram_rdata4[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1167.600 1767.600 1168.200 ;
    END
  END data_arrays_0_ext_ram_rdata4[15]
  PIN data_arrays_0_ext_ram_rdata4[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1173.040 1767.600 1173.640 ;
    END
  END data_arrays_0_ext_ram_rdata4[16]
  PIN data_arrays_0_ext_ram_rdata4[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1178.480 1767.600 1179.080 ;
    END
  END data_arrays_0_ext_ram_rdata4[17]
  PIN data_arrays_0_ext_ram_rdata4[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1183.920 1767.600 1184.520 ;
    END
  END data_arrays_0_ext_ram_rdata4[18]
  PIN data_arrays_0_ext_ram_rdata4[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1188.680 1767.600 1189.280 ;
    END
  END data_arrays_0_ext_ram_rdata4[19]
  PIN data_arrays_0_ext_ram_rdata4[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1091.440 1767.600 1092.040 ;
    END
  END data_arrays_0_ext_ram_rdata4[1]
  PIN data_arrays_0_ext_ram_rdata4[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1194.120 1767.600 1194.720 ;
    END
  END data_arrays_0_ext_ram_rdata4[20]
  PIN data_arrays_0_ext_ram_rdata4[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1199.560 1767.600 1200.160 ;
    END
  END data_arrays_0_ext_ram_rdata4[21]
  PIN data_arrays_0_ext_ram_rdata4[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1205.000 1767.600 1205.600 ;
    END
  END data_arrays_0_ext_ram_rdata4[22]
  PIN data_arrays_0_ext_ram_rdata4[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1210.440 1767.600 1211.040 ;
    END
  END data_arrays_0_ext_ram_rdata4[23]
  PIN data_arrays_0_ext_ram_rdata4[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1215.880 1767.600 1216.480 ;
    END
  END data_arrays_0_ext_ram_rdata4[24]
  PIN data_arrays_0_ext_ram_rdata4[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1221.320 1767.600 1221.920 ;
    END
  END data_arrays_0_ext_ram_rdata4[25]
  PIN data_arrays_0_ext_ram_rdata4[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1226.760 1767.600 1227.360 ;
    END
  END data_arrays_0_ext_ram_rdata4[26]
  PIN data_arrays_0_ext_ram_rdata4[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1232.200 1767.600 1232.800 ;
    END
  END data_arrays_0_ext_ram_rdata4[27]
  PIN data_arrays_0_ext_ram_rdata4[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1237.640 1767.600 1238.240 ;
    END
  END data_arrays_0_ext_ram_rdata4[28]
  PIN data_arrays_0_ext_ram_rdata4[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1243.080 1767.600 1243.680 ;
    END
  END data_arrays_0_ext_ram_rdata4[29]
  PIN data_arrays_0_ext_ram_rdata4[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1096.880 1767.600 1097.480 ;
    END
  END data_arrays_0_ext_ram_rdata4[2]
  PIN data_arrays_0_ext_ram_rdata4[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1248.520 1767.600 1249.120 ;
    END
  END data_arrays_0_ext_ram_rdata4[30]
  PIN data_arrays_0_ext_ram_rdata4[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1253.960 1767.600 1254.560 ;
    END
  END data_arrays_0_ext_ram_rdata4[31]
  PIN data_arrays_0_ext_ram_rdata4[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1102.320 1767.600 1102.920 ;
    END
  END data_arrays_0_ext_ram_rdata4[3]
  PIN data_arrays_0_ext_ram_rdata4[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1107.760 1767.600 1108.360 ;
    END
  END data_arrays_0_ext_ram_rdata4[4]
  PIN data_arrays_0_ext_ram_rdata4[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1113.200 1767.600 1113.800 ;
    END
  END data_arrays_0_ext_ram_rdata4[5]
  PIN data_arrays_0_ext_ram_rdata4[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1118.640 1767.600 1119.240 ;
    END
  END data_arrays_0_ext_ram_rdata4[6]
  PIN data_arrays_0_ext_ram_rdata4[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1124.080 1767.600 1124.680 ;
    END
  END data_arrays_0_ext_ram_rdata4[7]
  PIN data_arrays_0_ext_ram_rdata4[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1129.520 1767.600 1130.120 ;
    END
  END data_arrays_0_ext_ram_rdata4[8]
  PIN data_arrays_0_ext_ram_rdata4[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1134.960 1767.600 1135.560 ;
    END
  END data_arrays_0_ext_ram_rdata4[9]
  PIN data_arrays_0_ext_ram_rdata5[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1259.400 1767.600 1260.000 ;
    END
  END data_arrays_0_ext_ram_rdata5[0]
  PIN data_arrays_0_ext_ram_rdata5[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1313.800 1767.600 1314.400 ;
    END
  END data_arrays_0_ext_ram_rdata5[10]
  PIN data_arrays_0_ext_ram_rdata5[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1319.240 1767.600 1319.840 ;
    END
  END data_arrays_0_ext_ram_rdata5[11]
  PIN data_arrays_0_ext_ram_rdata5[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1324.680 1767.600 1325.280 ;
    END
  END data_arrays_0_ext_ram_rdata5[12]
  PIN data_arrays_0_ext_ram_rdata5[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1330.120 1767.600 1330.720 ;
    END
  END data_arrays_0_ext_ram_rdata5[13]
  PIN data_arrays_0_ext_ram_rdata5[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1335.560 1767.600 1336.160 ;
    END
  END data_arrays_0_ext_ram_rdata5[14]
  PIN data_arrays_0_ext_ram_rdata5[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1341.000 1767.600 1341.600 ;
    END
  END data_arrays_0_ext_ram_rdata5[15]
  PIN data_arrays_0_ext_ram_rdata5[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1346.440 1767.600 1347.040 ;
    END
  END data_arrays_0_ext_ram_rdata5[16]
  PIN data_arrays_0_ext_ram_rdata5[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1351.880 1767.600 1352.480 ;
    END
  END data_arrays_0_ext_ram_rdata5[17]
  PIN data_arrays_0_ext_ram_rdata5[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1357.320 1767.600 1357.920 ;
    END
  END data_arrays_0_ext_ram_rdata5[18]
  PIN data_arrays_0_ext_ram_rdata5[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1362.760 1767.600 1363.360 ;
    END
  END data_arrays_0_ext_ram_rdata5[19]
  PIN data_arrays_0_ext_ram_rdata5[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1264.840 1767.600 1265.440 ;
    END
  END data_arrays_0_ext_ram_rdata5[1]
  PIN data_arrays_0_ext_ram_rdata5[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1368.200 1767.600 1368.800 ;
    END
  END data_arrays_0_ext_ram_rdata5[20]
  PIN data_arrays_0_ext_ram_rdata5[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1373.640 1767.600 1374.240 ;
    END
  END data_arrays_0_ext_ram_rdata5[21]
  PIN data_arrays_0_ext_ram_rdata5[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1379.080 1767.600 1379.680 ;
    END
  END data_arrays_0_ext_ram_rdata5[22]
  PIN data_arrays_0_ext_ram_rdata5[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1384.520 1767.600 1385.120 ;
    END
  END data_arrays_0_ext_ram_rdata5[23]
  PIN data_arrays_0_ext_ram_rdata5[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1389.280 1767.600 1389.880 ;
    END
  END data_arrays_0_ext_ram_rdata5[24]
  PIN data_arrays_0_ext_ram_rdata5[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1394.720 1767.600 1395.320 ;
    END
  END data_arrays_0_ext_ram_rdata5[25]
  PIN data_arrays_0_ext_ram_rdata5[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1400.160 1767.600 1400.760 ;
    END
  END data_arrays_0_ext_ram_rdata5[26]
  PIN data_arrays_0_ext_ram_rdata5[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1405.600 1767.600 1406.200 ;
    END
  END data_arrays_0_ext_ram_rdata5[27]
  PIN data_arrays_0_ext_ram_rdata5[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1411.040 1767.600 1411.640 ;
    END
  END data_arrays_0_ext_ram_rdata5[28]
  PIN data_arrays_0_ext_ram_rdata5[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1416.480 1767.600 1417.080 ;
    END
  END data_arrays_0_ext_ram_rdata5[29]
  PIN data_arrays_0_ext_ram_rdata5[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1270.280 1767.600 1270.880 ;
    END
  END data_arrays_0_ext_ram_rdata5[2]
  PIN data_arrays_0_ext_ram_rdata5[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1421.920 1767.600 1422.520 ;
    END
  END data_arrays_0_ext_ram_rdata5[30]
  PIN data_arrays_0_ext_ram_rdata5[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1427.360 1767.600 1427.960 ;
    END
  END data_arrays_0_ext_ram_rdata5[31]
  PIN data_arrays_0_ext_ram_rdata5[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1275.720 1767.600 1276.320 ;
    END
  END data_arrays_0_ext_ram_rdata5[3]
  PIN data_arrays_0_ext_ram_rdata5[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1281.160 1767.600 1281.760 ;
    END
  END data_arrays_0_ext_ram_rdata5[4]
  PIN data_arrays_0_ext_ram_rdata5[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1286.600 1767.600 1287.200 ;
    END
  END data_arrays_0_ext_ram_rdata5[5]
  PIN data_arrays_0_ext_ram_rdata5[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1292.040 1767.600 1292.640 ;
    END
  END data_arrays_0_ext_ram_rdata5[6]
  PIN data_arrays_0_ext_ram_rdata5[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1297.480 1767.600 1298.080 ;
    END
  END data_arrays_0_ext_ram_rdata5[7]
  PIN data_arrays_0_ext_ram_rdata5[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1302.920 1767.600 1303.520 ;
    END
  END data_arrays_0_ext_ram_rdata5[8]
  PIN data_arrays_0_ext_ram_rdata5[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1308.360 1767.600 1308.960 ;
    END
  END data_arrays_0_ext_ram_rdata5[9]
  PIN data_arrays_0_ext_ram_rdata6[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1432.800 1767.600 1433.400 ;
    END
  END data_arrays_0_ext_ram_rdata6[0]
  PIN data_arrays_0_ext_ram_rdata6[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1487.200 1767.600 1487.800 ;
    END
  END data_arrays_0_ext_ram_rdata6[10]
  PIN data_arrays_0_ext_ram_rdata6[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1492.640 1767.600 1493.240 ;
    END
  END data_arrays_0_ext_ram_rdata6[11]
  PIN data_arrays_0_ext_ram_rdata6[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1498.080 1767.600 1498.680 ;
    END
  END data_arrays_0_ext_ram_rdata6[12]
  PIN data_arrays_0_ext_ram_rdata6[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1503.520 1767.600 1504.120 ;
    END
  END data_arrays_0_ext_ram_rdata6[13]
  PIN data_arrays_0_ext_ram_rdata6[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1508.960 1767.600 1509.560 ;
    END
  END data_arrays_0_ext_ram_rdata6[14]
  PIN data_arrays_0_ext_ram_rdata6[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1514.400 1767.600 1515.000 ;
    END
  END data_arrays_0_ext_ram_rdata6[15]
  PIN data_arrays_0_ext_ram_rdata6[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1519.840 1767.600 1520.440 ;
    END
  END data_arrays_0_ext_ram_rdata6[16]
  PIN data_arrays_0_ext_ram_rdata6[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1525.280 1767.600 1525.880 ;
    END
  END data_arrays_0_ext_ram_rdata6[17]
  PIN data_arrays_0_ext_ram_rdata6[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1530.720 1767.600 1531.320 ;
    END
  END data_arrays_0_ext_ram_rdata6[18]
  PIN data_arrays_0_ext_ram_rdata6[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1536.160 1767.600 1536.760 ;
    END
  END data_arrays_0_ext_ram_rdata6[19]
  PIN data_arrays_0_ext_ram_rdata6[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1438.240 1767.600 1438.840 ;
    END
  END data_arrays_0_ext_ram_rdata6[1]
  PIN data_arrays_0_ext_ram_rdata6[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1541.600 1767.600 1542.200 ;
    END
  END data_arrays_0_ext_ram_rdata6[20]
  PIN data_arrays_0_ext_ram_rdata6[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1547.040 1767.600 1547.640 ;
    END
  END data_arrays_0_ext_ram_rdata6[21]
  PIN data_arrays_0_ext_ram_rdata6[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1552.480 1767.600 1553.080 ;
    END
  END data_arrays_0_ext_ram_rdata6[22]
  PIN data_arrays_0_ext_ram_rdata6[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1557.920 1767.600 1558.520 ;
    END
  END data_arrays_0_ext_ram_rdata6[23]
  PIN data_arrays_0_ext_ram_rdata6[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1563.360 1767.600 1563.960 ;
    END
  END data_arrays_0_ext_ram_rdata6[24]
  PIN data_arrays_0_ext_ram_rdata6[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1568.800 1767.600 1569.400 ;
    END
  END data_arrays_0_ext_ram_rdata6[25]
  PIN data_arrays_0_ext_ram_rdata6[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1574.240 1767.600 1574.840 ;
    END
  END data_arrays_0_ext_ram_rdata6[26]
  PIN data_arrays_0_ext_ram_rdata6[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1579.680 1767.600 1580.280 ;
    END
  END data_arrays_0_ext_ram_rdata6[27]
  PIN data_arrays_0_ext_ram_rdata6[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1584.440 1767.600 1585.040 ;
    END
  END data_arrays_0_ext_ram_rdata6[28]
  PIN data_arrays_0_ext_ram_rdata6[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1589.880 1767.600 1590.480 ;
    END
  END data_arrays_0_ext_ram_rdata6[29]
  PIN data_arrays_0_ext_ram_rdata6[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1443.680 1767.600 1444.280 ;
    END
  END data_arrays_0_ext_ram_rdata6[2]
  PIN data_arrays_0_ext_ram_rdata6[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1595.320 1767.600 1595.920 ;
    END
  END data_arrays_0_ext_ram_rdata6[30]
  PIN data_arrays_0_ext_ram_rdata6[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1600.760 1767.600 1601.360 ;
    END
  END data_arrays_0_ext_ram_rdata6[31]
  PIN data_arrays_0_ext_ram_rdata6[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1449.120 1767.600 1449.720 ;
    END
  END data_arrays_0_ext_ram_rdata6[3]
  PIN data_arrays_0_ext_ram_rdata6[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1454.560 1767.600 1455.160 ;
    END
  END data_arrays_0_ext_ram_rdata6[4]
  PIN data_arrays_0_ext_ram_rdata6[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1460.000 1767.600 1460.600 ;
    END
  END data_arrays_0_ext_ram_rdata6[5]
  PIN data_arrays_0_ext_ram_rdata6[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1465.440 1767.600 1466.040 ;
    END
  END data_arrays_0_ext_ram_rdata6[6]
  PIN data_arrays_0_ext_ram_rdata6[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1470.880 1767.600 1471.480 ;
    END
  END data_arrays_0_ext_ram_rdata6[7]
  PIN data_arrays_0_ext_ram_rdata6[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1476.320 1767.600 1476.920 ;
    END
  END data_arrays_0_ext_ram_rdata6[8]
  PIN data_arrays_0_ext_ram_rdata6[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1481.760 1767.600 1482.360 ;
    END
  END data_arrays_0_ext_ram_rdata6[9]
  PIN data_arrays_0_ext_ram_rdata7[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1606.200 1767.600 1606.800 ;
    END
  END data_arrays_0_ext_ram_rdata7[0]
  PIN data_arrays_0_ext_ram_rdata7[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1660.600 1767.600 1661.200 ;
    END
  END data_arrays_0_ext_ram_rdata7[10]
  PIN data_arrays_0_ext_ram_rdata7[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1666.040 1767.600 1666.640 ;
    END
  END data_arrays_0_ext_ram_rdata7[11]
  PIN data_arrays_0_ext_ram_rdata7[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1671.480 1767.600 1672.080 ;
    END
  END data_arrays_0_ext_ram_rdata7[12]
  PIN data_arrays_0_ext_ram_rdata7[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1676.920 1767.600 1677.520 ;
    END
  END data_arrays_0_ext_ram_rdata7[13]
  PIN data_arrays_0_ext_ram_rdata7[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1682.360 1767.600 1682.960 ;
    END
  END data_arrays_0_ext_ram_rdata7[14]
  PIN data_arrays_0_ext_ram_rdata7[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1687.800 1767.600 1688.400 ;
    END
  END data_arrays_0_ext_ram_rdata7[15]
  PIN data_arrays_0_ext_ram_rdata7[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1693.240 1767.600 1693.840 ;
    END
  END data_arrays_0_ext_ram_rdata7[16]
  PIN data_arrays_0_ext_ram_rdata7[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1698.680 1767.600 1699.280 ;
    END
  END data_arrays_0_ext_ram_rdata7[17]
  PIN data_arrays_0_ext_ram_rdata7[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1704.120 1767.600 1704.720 ;
    END
  END data_arrays_0_ext_ram_rdata7[18]
  PIN data_arrays_0_ext_ram_rdata7[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1709.560 1767.600 1710.160 ;
    END
  END data_arrays_0_ext_ram_rdata7[19]
  PIN data_arrays_0_ext_ram_rdata7[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1611.640 1767.600 1612.240 ;
    END
  END data_arrays_0_ext_ram_rdata7[1]
  PIN data_arrays_0_ext_ram_rdata7[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1715.000 1767.600 1715.600 ;
    END
  END data_arrays_0_ext_ram_rdata7[20]
  PIN data_arrays_0_ext_ram_rdata7[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1720.440 1767.600 1721.040 ;
    END
  END data_arrays_0_ext_ram_rdata7[21]
  PIN data_arrays_0_ext_ram_rdata7[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1725.880 1767.600 1726.480 ;
    END
  END data_arrays_0_ext_ram_rdata7[22]
  PIN data_arrays_0_ext_ram_rdata7[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1731.320 1767.600 1731.920 ;
    END
  END data_arrays_0_ext_ram_rdata7[23]
  PIN data_arrays_0_ext_ram_rdata7[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1736.760 1767.600 1737.360 ;
    END
  END data_arrays_0_ext_ram_rdata7[24]
  PIN data_arrays_0_ext_ram_rdata7[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1742.200 1767.600 1742.800 ;
    END
  END data_arrays_0_ext_ram_rdata7[25]
  PIN data_arrays_0_ext_ram_rdata7[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1747.640 1767.600 1748.240 ;
    END
  END data_arrays_0_ext_ram_rdata7[26]
  PIN data_arrays_0_ext_ram_rdata7[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1753.080 1767.600 1753.680 ;
    END
  END data_arrays_0_ext_ram_rdata7[27]
  PIN data_arrays_0_ext_ram_rdata7[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1758.520 1767.600 1759.120 ;
    END
  END data_arrays_0_ext_ram_rdata7[28]
  PIN data_arrays_0_ext_ram_rdata7[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1763.960 1767.600 1764.560 ;
    END
  END data_arrays_0_ext_ram_rdata7[29]
  PIN data_arrays_0_ext_ram_rdata7[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1617.080 1767.600 1617.680 ;
    END
  END data_arrays_0_ext_ram_rdata7[2]
  PIN data_arrays_0_ext_ram_rdata7[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1769.400 1767.600 1770.000 ;
    END
  END data_arrays_0_ext_ram_rdata7[30]
  PIN data_arrays_0_ext_ram_rdata7[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1774.840 1767.600 1775.440 ;
    END
  END data_arrays_0_ext_ram_rdata7[31]
  PIN data_arrays_0_ext_ram_rdata7[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1622.520 1767.600 1623.120 ;
    END
  END data_arrays_0_ext_ram_rdata7[3]
  PIN data_arrays_0_ext_ram_rdata7[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1627.960 1767.600 1628.560 ;
    END
  END data_arrays_0_ext_ram_rdata7[4]
  PIN data_arrays_0_ext_ram_rdata7[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1633.400 1767.600 1634.000 ;
    END
  END data_arrays_0_ext_ram_rdata7[5]
  PIN data_arrays_0_ext_ram_rdata7[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1638.840 1767.600 1639.440 ;
    END
  END data_arrays_0_ext_ram_rdata7[6]
  PIN data_arrays_0_ext_ram_rdata7[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1644.280 1767.600 1644.880 ;
    END
  END data_arrays_0_ext_ram_rdata7[7]
  PIN data_arrays_0_ext_ram_rdata7[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1649.720 1767.600 1650.320 ;
    END
  END data_arrays_0_ext_ram_rdata7[8]
  PIN data_arrays_0_ext_ram_rdata7[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 1655.160 1767.600 1655.760 ;
    END
  END data_arrays_0_ext_ram_rdata7[9]
  PIN data_arrays_0_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 750.080 1767.600 750.680 ;
    END
  END data_arrays_0_ext_ram_wdata[0]
  PIN data_arrays_0_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 803.800 1767.600 804.400 ;
    END
  END data_arrays_0_ext_ram_wdata[10]
  PIN data_arrays_0_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 809.240 1767.600 809.840 ;
    END
  END data_arrays_0_ext_ram_wdata[11]
  PIN data_arrays_0_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 814.680 1767.600 815.280 ;
    END
  END data_arrays_0_ext_ram_wdata[12]
  PIN data_arrays_0_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 820.120 1767.600 820.720 ;
    END
  END data_arrays_0_ext_ram_wdata[13]
  PIN data_arrays_0_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 825.560 1767.600 826.160 ;
    END
  END data_arrays_0_ext_ram_wdata[14]
  PIN data_arrays_0_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 831.000 1767.600 831.600 ;
    END
  END data_arrays_0_ext_ram_wdata[15]
  PIN data_arrays_0_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 836.440 1767.600 837.040 ;
    END
  END data_arrays_0_ext_ram_wdata[16]
  PIN data_arrays_0_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 841.880 1767.600 842.480 ;
    END
  END data_arrays_0_ext_ram_wdata[17]
  PIN data_arrays_0_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 847.320 1767.600 847.920 ;
    END
  END data_arrays_0_ext_ram_wdata[18]
  PIN data_arrays_0_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 852.760 1767.600 853.360 ;
    END
  END data_arrays_0_ext_ram_wdata[19]
  PIN data_arrays_0_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 755.520 1767.600 756.120 ;
    END
  END data_arrays_0_ext_ram_wdata[1]
  PIN data_arrays_0_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 858.200 1767.600 858.800 ;
    END
  END data_arrays_0_ext_ram_wdata[20]
  PIN data_arrays_0_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 863.640 1767.600 864.240 ;
    END
  END data_arrays_0_ext_ram_wdata[21]
  PIN data_arrays_0_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 869.080 1767.600 869.680 ;
    END
  END data_arrays_0_ext_ram_wdata[22]
  PIN data_arrays_0_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 874.520 1767.600 875.120 ;
    END
  END data_arrays_0_ext_ram_wdata[23]
  PIN data_arrays_0_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 879.960 1767.600 880.560 ;
    END
  END data_arrays_0_ext_ram_wdata[24]
  PIN data_arrays_0_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 885.400 1767.600 886.000 ;
    END
  END data_arrays_0_ext_ram_wdata[25]
  PIN data_arrays_0_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 890.840 1767.600 891.440 ;
    END
  END data_arrays_0_ext_ram_wdata[26]
  PIN data_arrays_0_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 896.280 1767.600 896.880 ;
    END
  END data_arrays_0_ext_ram_wdata[27]
  PIN data_arrays_0_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 901.720 1767.600 902.320 ;
    END
  END data_arrays_0_ext_ram_wdata[28]
  PIN data_arrays_0_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 907.160 1767.600 907.760 ;
    END
  END data_arrays_0_ext_ram_wdata[29]
  PIN data_arrays_0_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 760.960 1767.600 761.560 ;
    END
  END data_arrays_0_ext_ram_wdata[2]
  PIN data_arrays_0_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 912.600 1767.600 913.200 ;
    END
  END data_arrays_0_ext_ram_wdata[30]
  PIN data_arrays_0_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 918.040 1767.600 918.640 ;
    END
  END data_arrays_0_ext_ram_wdata[31]
  PIN data_arrays_0_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 766.400 1767.600 767.000 ;
    END
  END data_arrays_0_ext_ram_wdata[3]
  PIN data_arrays_0_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 771.840 1767.600 772.440 ;
    END
  END data_arrays_0_ext_ram_wdata[4]
  PIN data_arrays_0_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 777.280 1767.600 777.880 ;
    END
  END data_arrays_0_ext_ram_wdata[5]
  PIN data_arrays_0_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 782.720 1767.600 783.320 ;
    END
  END data_arrays_0_ext_ram_wdata[6]
  PIN data_arrays_0_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 788.160 1767.600 788.760 ;
    END
  END data_arrays_0_ext_ram_wdata[7]
  PIN data_arrays_0_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 792.920 1767.600 793.520 ;
    END
  END data_arrays_0_ext_ram_wdata[8]
  PIN data_arrays_0_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 798.360 1767.600 798.960 ;
    END
  END data_arrays_0_ext_ram_wdata[9]
  PIN data_arrays_0_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 988.760 1767.600 989.360 ;
    END
  END data_arrays_0_ext_ram_web
  PIN data_arrays_0_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 923.480 1767.600 924.080 ;
    END
  END data_arrays_0_ext_ram_wmask[0]
  PIN data_arrays_0_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 928.920 1767.600 929.520 ;
    END
  END data_arrays_0_ext_ram_wmask[1]
  PIN data_arrays_0_ext_ram_wmask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 934.360 1767.600 934.960 ;
    END
  END data_arrays_0_ext_ram_wmask[2]
  PIN data_arrays_0_ext_ram_wmask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.600 939.800 1767.600 940.400 ;
    END
  END data_arrays_0_ext_ram_wmask[3]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 1774.320 7.730 1778.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 1774.320 472.790 1778.320 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 1774.320 519.250 1778.320 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 1774.320 565.710 1778.320 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1774.320 612.170 1778.320 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 1774.320 658.630 1778.320 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 1774.320 705.090 1778.320 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 1774.320 752.010 1778.320 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 1774.320 798.470 1778.320 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 1774.320 844.930 1778.320 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 1774.320 891.390 1778.320 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 1774.320 54.190 1778.320 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 1774.320 937.850 1778.320 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 1774.320 984.310 1778.320 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 1774.320 1030.770 1778.320 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.410 1774.320 1077.690 1778.320 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 1774.320 1124.150 1778.320 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.330 1774.320 1170.610 1778.320 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.790 1774.320 1217.070 1778.320 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.250 1774.320 1263.530 1778.320 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 1774.320 1309.990 1778.320 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.170 1774.320 1356.450 1778.320 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 1774.320 100.650 1778.320 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.630 1774.320 1402.910 1778.320 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.550 1774.320 1449.830 1778.320 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.010 1774.320 1496.290 1778.320 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 1774.320 1542.750 1778.320 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.930 1774.320 1589.210 1778.320 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.390 1774.320 1635.670 1778.320 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.850 1774.320 1682.130 1778.320 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.310 1774.320 1728.590 1778.320 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 1774.320 147.110 1778.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1774.320 193.570 1778.320 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 1774.320 240.030 1778.320 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 1774.320 286.490 1778.320 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 1774.320 332.950 1778.320 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 1774.320 379.870 1778.320 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 1774.320 426.330 1778.320 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1774.320 22.910 1778.320 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 1774.320 488.430 1778.320 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 1774.320 534.890 1778.320 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 1774.320 581.350 1778.320 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 1774.320 627.810 1778.320 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 1774.320 674.270 1778.320 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 1774.320 720.730 1778.320 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 1774.320 767.190 1778.320 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 1774.320 813.650 1778.320 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 1774.320 860.570 1778.320 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 1774.320 907.030 1778.320 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 1774.320 69.370 1778.320 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 1774.320 953.490 1778.320 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 1774.320 999.950 1778.320 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 1774.320 1046.410 1778.320 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 1774.320 1092.870 1778.320 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.050 1774.320 1139.330 1778.320 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.970 1774.320 1186.250 1778.320 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.430 1774.320 1232.710 1778.320 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.890 1774.320 1279.170 1778.320 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.350 1774.320 1325.630 1778.320 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 1774.320 1372.090 1778.320 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 1774.320 115.830 1778.320 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.270 1774.320 1418.550 1778.320 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.730 1774.320 1465.010 1778.320 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.190 1774.320 1511.470 1778.320 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.110 1774.320 1558.390 1778.320 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.570 1774.320 1604.850 1778.320 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.030 1774.320 1651.310 1778.320 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.490 1774.320 1697.770 1778.320 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.950 1774.320 1744.230 1778.320 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 1774.320 162.750 1778.320 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 1774.320 209.210 1778.320 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 1774.320 255.670 1778.320 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 1774.320 302.130 1778.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 1774.320 348.590 1778.320 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 1774.320 395.050 1778.320 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 1774.320 441.510 1778.320 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 1774.320 38.550 1778.320 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 1774.320 503.610 1778.320 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 1774.320 550.070 1778.320 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 1774.320 596.990 1778.320 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 1774.320 643.450 1778.320 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 1774.320 689.910 1778.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 1774.320 736.370 1778.320 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 1774.320 782.830 1778.320 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 1774.320 829.290 1778.320 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.470 1774.320 875.750 1778.320 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 1774.320 922.210 1778.320 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 1774.320 85.010 1778.320 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 1774.320 969.130 1778.320 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.310 1774.320 1015.590 1778.320 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.770 1774.320 1062.050 1778.320 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.230 1774.320 1108.510 1778.320 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 1774.320 1154.970 1778.320 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 1774.320 1201.430 1778.320 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 1774.320 1247.890 1778.320 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.070 1774.320 1294.350 1778.320 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 1774.320 1341.270 1778.320 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.450 1774.320 1387.730 1778.320 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 1774.320 131.470 1778.320 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.910 1774.320 1434.190 1778.320 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.370 1774.320 1480.650 1778.320 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.830 1774.320 1527.110 1778.320 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.290 1774.320 1573.570 1778.320 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.750 1774.320 1620.030 1778.320 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.670 1774.320 1666.950 1778.320 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 1774.320 1713.410 1778.320 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1759.590 1774.320 1759.870 1778.320 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 1774.320 177.930 1778.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 1774.320 224.390 1778.320 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 1774.320 271.310 1778.320 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 1774.320 317.770 1778.320 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1774.320 364.230 1778.320 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 1774.320 410.690 1778.320 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 1774.320 457.150 1778.320 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.890 0.000 1762.170 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.570 0.000 1765.850 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.910 0.000 1457.190 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.950 0.000 1468.230 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.530 0.000 1478.810 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 0.000 1489.390 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.150 0.000 1500.430 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 0.000 1511.010 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.770 0.000 1522.050 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.350 0.000 1532.630 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 0.000 1543.210 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.970 0.000 1554.250 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.550 0.000 1564.830 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.590 0.000 1575.870 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.170 0.000 1586.450 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.750 0.000 1597.030 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.790 0.000 1608.070 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.370 0.000 1618.650 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.950 0.000 1629.230 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.990 0.000 1640.270 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.570 0.000 1650.850 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 0.000 1661.890 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 0.000 1672.470 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.770 0.000 1683.050 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.390 0.000 1704.670 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.430 0.000 1715.710 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 0.000 1726.290 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.590 0.000 1736.870 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.630 0.000 1747.910 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 0.000 510.510 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 0.000 725.790 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 0.000 757.990 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 0.000 865.630 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 0.000 887.250 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 0.000 908.870 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.170 0.000 919.450 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 0.000 930.030 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.790 0.000 941.070 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 0.000 951.650 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.990 0.000 973.270 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 0.000 983.850 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 0.000 1016.510 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.810 0.000 1027.090 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 0.000 1059.290 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 0.000 1080.910 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.830 0.000 1113.110 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.410 0.000 1123.690 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.650 0.000 1166.930 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 0.000 1177.510 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.850 0.000 1199.130 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.430 0.000 1209.710 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 0.000 1220.750 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 0.000 1231.330 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.090 0.000 1242.370 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.250 0.000 1263.530 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.290 0.000 1274.570 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 0.000 1285.150 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.910 0.000 1296.190 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.490 0.000 1306.770 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.110 0.000 1328.390 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.690 0.000 1338.970 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.310 0.000 1360.590 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.890 0.000 1371.170 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 0.000 1382.210 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.510 0.000 1392.790 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 0.000 1403.370 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.130 0.000 1414.410 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.710 0.000 1424.990 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.750 0.000 1436.030 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 0.000 1446.610 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.590 0.000 1460.870 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.210 0.000 1482.490 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 0.000 1493.070 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 0.000 1504.110 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.410 0.000 1514.690 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.990 0.000 1525.270 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 0.000 1536.310 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.610 0.000 1546.890 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.650 0.000 1557.930 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 0.000 1568.510 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.810 0.000 1579.090 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.850 0.000 1590.130 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.430 0.000 1600.710 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.050 0.000 1622.330 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 0.000 1632.910 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.670 0.000 1643.950 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.250 0.000 1654.530 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.830 0.000 1665.110 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.870 0.000 1676.150 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.450 0.000 1686.730 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.490 0.000 1697.770 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.070 0.000 1708.350 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.650 0.000 1718.930 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.690 0.000 1729.970 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.270 0.000 1740.550 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.310 0.000 1751.590 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 0.000 665.070 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 0.000 675.650 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 0.000 751.090 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 0.000 826.070 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.830 0.000 837.110 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 0.000 847.690 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 0.000 858.730 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 0.000 869.310 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.650 0.000 890.930 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 0.000 912.090 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.850 0.000 923.130 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 0.000 933.710 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.470 0.000 944.750 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.630 0.000 965.910 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 0.000 976.950 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.870 0.000 1009.150 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.450 0.000 1019.730 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.070 0.000 1041.350 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 0.000 1051.930 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 0.000 1073.550 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 0.000 1084.590 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.470 0.000 1105.750 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 0.000 1116.790 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.710 0.000 1148.990 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.330 0.000 1170.610 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 0.000 1191.770 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.530 0.000 1202.810 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.110 0.000 1213.390 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 0.000 1224.430 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.730 0.000 1235.010 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.310 0.000 1245.590 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.350 0.000 1256.630 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 0.000 1267.210 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.970 0.000 1278.250 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.550 0.000 1288.830 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.170 0.000 1310.450 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 0.000 1321.030 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.330 0.000 1331.610 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 0.000 1364.270 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.570 0.000 1374.850 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.190 0.000 1396.470 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.770 0.000 1407.050 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.810 0.000 1418.090 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.390 0.000 1428.670 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.970 0.000 1439.250 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.010 0.000 1450.290 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 0.000 1464.550 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.890 0.000 1486.170 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.470 0.000 1496.750 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 0.000 1507.330 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.090 0.000 1518.370 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.670 0.000 1528.950 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.710 0.000 1539.990 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.290 0.000 1550.570 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.870 0.000 1561.150 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.910 0.000 1572.190 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.490 0.000 1582.770 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.530 0.000 1593.810 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.110 0.000 1604.390 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.690 0.000 1614.970 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 0.000 1626.010 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.310 0.000 1636.590 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.890 0.000 1647.170 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.930 0.000 1658.210 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.510 0.000 1668.790 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.550 0.000 1679.830 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.130 0.000 1690.410 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.710 0.000 1700.990 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.750 0.000 1712.030 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.330 0.000 1722.610 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.370 0.000 1733.650 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.950 0.000 1744.230 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.530 0.000 1754.810 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 0.000 625.510 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 0.000 722.110 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 0.000 743.730 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.070 0.000 765.350 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 0.000 819.170 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 0.000 883.570 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 0.000 894.150 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 0.000 915.770 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.530 0.000 926.810 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.690 0.000 947.970 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.930 0.000 991.210 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 0.000 1012.830 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 0.000 1023.410 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 0.000 1045.030 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.330 0.000 1055.610 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 0.000 1066.650 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 0.000 1077.230 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 0.000 1087.810 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 0.000 1109.430 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.770 0.000 1131.050 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 0.000 1141.630 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.390 0.000 1152.670 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.970 0.000 1163.250 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 0.000 1174.290 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.590 0.000 1184.870 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.210 0.000 1206.490 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.790 0.000 1217.070 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 0.000 1227.650 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 0.000 1238.690 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990 0.000 1249.270 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.030 0.000 1260.310 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1270.610 0.000 1270.890 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.190 0.000 1281.470 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.230 0.000 1292.510 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.810 0.000 1303.090 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 0.000 1314.130 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.430 0.000 1324.710 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.010 0.000 1335.290 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.630 0.000 1356.910 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.210 0.000 1367.490 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 0.000 1378.530 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.830 0.000 1389.110 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.870 0.000 1400.150 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 0.000 1421.310 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.070 0.000 1432.350 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 0.000 1442.930 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 0.000 1453.970 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END la_oenb[9]
  PIN tag_array_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.160 4.000 1638.760 ;
    END
  END tag_array_ext_ram_addr1[0]
  PIN tag_array_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1642.240 4.000 1642.840 ;
    END
  END tag_array_ext_ram_addr1[1]
  PIN tag_array_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1645.640 4.000 1646.240 ;
    END
  END tag_array_ext_ram_addr1[2]
  PIN tag_array_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1649.040 4.000 1649.640 ;
    END
  END tag_array_ext_ram_addr1[3]
  PIN tag_array_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1652.440 4.000 1653.040 ;
    END
  END tag_array_ext_ram_addr1[4]
  PIN tag_array_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1655.840 4.000 1656.440 ;
    END
  END tag_array_ext_ram_addr1[5]
  PIN tag_array_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END tag_array_ext_ram_addr1[6]
  PIN tag_array_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1663.320 4.000 1663.920 ;
    END
  END tag_array_ext_ram_addr1[7]
  PIN tag_array_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END tag_array_ext_ram_addr[0]
  PIN tag_array_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1363.440 4.000 1364.040 ;
    END
  END tag_array_ext_ram_addr[1]
  PIN tag_array_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1367.520 4.000 1368.120 ;
    END
  END tag_array_ext_ram_addr[2]
  PIN tag_array_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.920 4.000 1371.520 ;
    END
  END tag_array_ext_ram_addr[3]
  PIN tag_array_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1374.320 4.000 1374.920 ;
    END
  END tag_array_ext_ram_addr[4]
  PIN tag_array_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.720 4.000 1378.320 ;
    END
  END tag_array_ext_ram_addr[5]
  PIN tag_array_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1381.120 4.000 1381.720 ;
    END
  END tag_array_ext_ram_addr[6]
  PIN tag_array_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1385.200 4.000 1385.800 ;
    END
  END tag_array_ext_ram_addr[7]
  PIN tag_array_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1388.600 4.000 1389.200 ;
    END
  END tag_array_ext_ram_clk
  PIN tag_array_ext_ram_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1624.560 4.000 1625.160 ;
    END
  END tag_array_ext_ram_csb
  PIN tag_array_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1631.360 4.000 1631.960 ;
    END
  END tag_array_ext_ram_csb1[0]
  PIN tag_array_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1634.760 4.000 1635.360 ;
    END
  END tag_array_ext_ram_csb1[1]
  PIN tag_array_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END tag_array_ext_ram_rdata0[0]
  PIN tag_array_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1282.520 4.000 1283.120 ;
    END
  END tag_array_ext_ram_rdata0[10]
  PIN tag_array_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1286.600 4.000 1287.200 ;
    END
  END tag_array_ext_ram_rdata0[11]
  PIN tag_array_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1290.000 4.000 1290.600 ;
    END
  END tag_array_ext_ram_rdata0[12]
  PIN tag_array_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END tag_array_ext_ram_rdata0[13]
  PIN tag_array_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1296.800 4.000 1297.400 ;
    END
  END tag_array_ext_ram_rdata0[14]
  PIN tag_array_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.200 4.000 1300.800 ;
    END
  END tag_array_ext_ram_rdata0[15]
  PIN tag_array_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1303.600 4.000 1304.200 ;
    END
  END tag_array_ext_ram_rdata0[16]
  PIN tag_array_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1307.680 4.000 1308.280 ;
    END
  END tag_array_ext_ram_rdata0[17]
  PIN tag_array_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1311.080 4.000 1311.680 ;
    END
  END tag_array_ext_ram_rdata0[18]
  PIN tag_array_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1314.480 4.000 1315.080 ;
    END
  END tag_array_ext_ram_rdata0[19]
  PIN tag_array_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.240 4.000 1251.840 ;
    END
  END tag_array_ext_ram_rdata0[1]
  PIN tag_array_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1317.880 4.000 1318.480 ;
    END
  END tag_array_ext_ram_rdata0[20]
  PIN tag_array_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1321.280 4.000 1321.880 ;
    END
  END tag_array_ext_ram_rdata0[21]
  PIN tag_array_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1325.360 4.000 1325.960 ;
    END
  END tag_array_ext_ram_rdata0[22]
  PIN tag_array_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1328.760 4.000 1329.360 ;
    END
  END tag_array_ext_ram_rdata0[23]
  PIN tag_array_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.160 4.000 1332.760 ;
    END
  END tag_array_ext_ram_rdata0[24]
  PIN tag_array_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1335.560 4.000 1336.160 ;
    END
  END tag_array_ext_ram_rdata0[25]
  PIN tag_array_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1338.960 4.000 1339.560 ;
    END
  END tag_array_ext_ram_rdata0[26]
  PIN tag_array_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1342.360 4.000 1342.960 ;
    END
  END tag_array_ext_ram_rdata0[27]
  PIN tag_array_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1346.440 4.000 1347.040 ;
    END
  END tag_array_ext_ram_rdata0[28]
  PIN tag_array_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.840 4.000 1350.440 ;
    END
  END tag_array_ext_ram_rdata0[29]
  PIN tag_array_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END tag_array_ext_ram_rdata0[2]
  PIN tag_array_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END tag_array_ext_ram_rdata0[30]
  PIN tag_array_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1356.640 4.000 1357.240 ;
    END
  END tag_array_ext_ram_rdata0[31]
  PIN tag_array_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END tag_array_ext_ram_rdata0[3]
  PIN tag_array_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END tag_array_ext_ram_rdata0[4]
  PIN tag_array_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END tag_array_ext_ram_rdata0[5]
  PIN tag_array_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.920 4.000 1269.520 ;
    END
  END tag_array_ext_ram_rdata0[6]
  PIN tag_array_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1272.320 4.000 1272.920 ;
    END
  END tag_array_ext_ram_rdata0[7]
  PIN tag_array_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.720 4.000 1276.320 ;
    END
  END tag_array_ext_ram_rdata0[8]
  PIN tag_array_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.120 4.000 1279.720 ;
    END
  END tag_array_ext_ram_rdata0[9]
  PIN tag_array_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.720 4.000 1667.320 ;
    END
  END tag_array_ext_ram_rdata1[0]
  PIN tag_array_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1702.080 4.000 1702.680 ;
    END
  END tag_array_ext_ram_rdata1[10]
  PIN tag_array_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1705.480 4.000 1706.080 ;
    END
  END tag_array_ext_ram_rdata1[11]
  PIN tag_array_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1708.880 4.000 1709.480 ;
    END
  END tag_array_ext_ram_rdata1[12]
  PIN tag_array_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1712.280 4.000 1712.880 ;
    END
  END tag_array_ext_ram_rdata1[13]
  PIN tag_array_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.680 4.000 1716.280 ;
    END
  END tag_array_ext_ram_rdata1[14]
  PIN tag_array_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1719.080 4.000 1719.680 ;
    END
  END tag_array_ext_ram_rdata1[15]
  PIN tag_array_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.160 4.000 1723.760 ;
    END
  END tag_array_ext_ram_rdata1[16]
  PIN tag_array_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1726.560 4.000 1727.160 ;
    END
  END tag_array_ext_ram_rdata1[17]
  PIN tag_array_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1729.960 4.000 1730.560 ;
    END
  END tag_array_ext_ram_rdata1[18]
  PIN tag_array_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1733.360 4.000 1733.960 ;
    END
  END tag_array_ext_ram_rdata1[19]
  PIN tag_array_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1670.120 4.000 1670.720 ;
    END
  END tag_array_ext_ram_rdata1[1]
  PIN tag_array_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1736.760 4.000 1737.360 ;
    END
  END tag_array_ext_ram_rdata1[20]
  PIN tag_array_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1740.840 4.000 1741.440 ;
    END
  END tag_array_ext_ram_rdata1[21]
  PIN tag_array_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1744.240 4.000 1744.840 ;
    END
  END tag_array_ext_ram_rdata1[22]
  PIN tag_array_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END tag_array_ext_ram_rdata1[23]
  PIN tag_array_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.040 4.000 1751.640 ;
    END
  END tag_array_ext_ram_rdata1[24]
  PIN tag_array_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1754.440 4.000 1755.040 ;
    END
  END tag_array_ext_ram_rdata1[25]
  PIN tag_array_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.840 4.000 1758.440 ;
    END
  END tag_array_ext_ram_rdata1[26]
  PIN tag_array_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1761.920 4.000 1762.520 ;
    END
  END tag_array_ext_ram_rdata1[27]
  PIN tag_array_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1765.320 4.000 1765.920 ;
    END
  END tag_array_ext_ram_rdata1[28]
  PIN tag_array_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.720 4.000 1769.320 ;
    END
  END tag_array_ext_ram_rdata1[29]
  PIN tag_array_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1673.520 4.000 1674.120 ;
    END
  END tag_array_ext_ram_rdata1[2]
  PIN tag_array_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1772.120 4.000 1772.720 ;
    END
  END tag_array_ext_ram_rdata1[30]
  PIN tag_array_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1775.520 4.000 1776.120 ;
    END
  END tag_array_ext_ram_rdata1[31]
  PIN tag_array_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1676.920 4.000 1677.520 ;
    END
  END tag_array_ext_ram_rdata1[3]
  PIN tag_array_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1681.000 4.000 1681.600 ;
    END
  END tag_array_ext_ram_rdata1[4]
  PIN tag_array_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1684.400 4.000 1685.000 ;
    END
  END tag_array_ext_ram_rdata1[5]
  PIN tag_array_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1687.800 4.000 1688.400 ;
    END
  END tag_array_ext_ram_rdata1[6]
  PIN tag_array_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1691.200 4.000 1691.800 ;
    END
  END tag_array_ext_ram_rdata1[7]
  PIN tag_array_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1694.600 4.000 1695.200 ;
    END
  END tag_array_ext_ram_rdata1[8]
  PIN tag_array_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1698.000 4.000 1698.600 ;
    END
  END tag_array_ext_ram_rdata1[9]
  PIN tag_array_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.000 4.000 1392.600 ;
    END
  END tag_array_ext_ram_wdata[0]
  PIN tag_array_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1427.360 4.000 1427.960 ;
    END
  END tag_array_ext_ram_wdata[10]
  PIN tag_array_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1430.760 4.000 1431.360 ;
    END
  END tag_array_ext_ram_wdata[11]
  PIN tag_array_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.160 4.000 1434.760 ;
    END
  END tag_array_ext_ram_wdata[12]
  PIN tag_array_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1437.560 4.000 1438.160 ;
    END
  END tag_array_ext_ram_wdata[13]
  PIN tag_array_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1440.960 4.000 1441.560 ;
    END
  END tag_array_ext_ram_wdata[14]
  PIN tag_array_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.040 4.000 1445.640 ;
    END
  END tag_array_ext_ram_wdata[15]
  PIN tag_array_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 4.000 1449.040 ;
    END
  END tag_array_ext_ram_wdata[16]
  PIN tag_array_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.840 4.000 1452.440 ;
    END
  END tag_array_ext_ram_wdata[17]
  PIN tag_array_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END tag_array_ext_ram_wdata[18]
  PIN tag_array_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END tag_array_ext_ram_wdata[19]
  PIN tag_array_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1395.400 4.000 1396.000 ;
    END
  END tag_array_ext_ram_wdata[1]
  PIN tag_array_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END tag_array_ext_ram_wdata[20]
  PIN tag_array_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1466.120 4.000 1466.720 ;
    END
  END tag_array_ext_ram_wdata[21]
  PIN tag_array_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1469.520 4.000 1470.120 ;
    END
  END tag_array_ext_ram_wdata[22]
  PIN tag_array_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.920 4.000 1473.520 ;
    END
  END tag_array_ext_ram_wdata[23]
  PIN tag_array_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1476.320 4.000 1476.920 ;
    END
  END tag_array_ext_ram_wdata[24]
  PIN tag_array_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.720 4.000 1480.320 ;
    END
  END tag_array_ext_ram_wdata[25]
  PIN tag_array_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1483.800 4.000 1484.400 ;
    END
  END tag_array_ext_ram_wdata[26]
  PIN tag_array_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1487.200 4.000 1487.800 ;
    END
  END tag_array_ext_ram_wdata[27]
  PIN tag_array_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1490.600 4.000 1491.200 ;
    END
  END tag_array_ext_ram_wdata[28]
  PIN tag_array_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1494.000 4.000 1494.600 ;
    END
  END tag_array_ext_ram_wdata[29]
  PIN tag_array_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1398.800 4.000 1399.400 ;
    END
  END tag_array_ext_ram_wdata[2]
  PIN tag_array_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1497.400 4.000 1498.000 ;
    END
  END tag_array_ext_ram_wdata[30]
  PIN tag_array_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1500.800 4.000 1501.400 ;
    END
  END tag_array_ext_ram_wdata[31]
  PIN tag_array_ext_ram_wdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1504.880 4.000 1505.480 ;
    END
  END tag_array_ext_ram_wdata[32]
  PIN tag_array_ext_ram_wdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1508.280 4.000 1508.880 ;
    END
  END tag_array_ext_ram_wdata[33]
  PIN tag_array_ext_ram_wdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1511.680 4.000 1512.280 ;
    END
  END tag_array_ext_ram_wdata[34]
  PIN tag_array_ext_ram_wdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1515.080 4.000 1515.680 ;
    END
  END tag_array_ext_ram_wdata[35]
  PIN tag_array_ext_ram_wdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1518.480 4.000 1519.080 ;
    END
  END tag_array_ext_ram_wdata[36]
  PIN tag_array_ext_ram_wdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1521.880 4.000 1522.480 ;
    END
  END tag_array_ext_ram_wdata[37]
  PIN tag_array_ext_ram_wdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1525.960 4.000 1526.560 ;
    END
  END tag_array_ext_ram_wdata[38]
  PIN tag_array_ext_ram_wdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1529.360 4.000 1529.960 ;
    END
  END tag_array_ext_ram_wdata[39]
  PIN tag_array_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1402.200 4.000 1402.800 ;
    END
  END tag_array_ext_ram_wdata[3]
  PIN tag_array_ext_ram_wdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1532.760 4.000 1533.360 ;
    END
  END tag_array_ext_ram_wdata[40]
  PIN tag_array_ext_ram_wdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.160 4.000 1536.760 ;
    END
  END tag_array_ext_ram_wdata[41]
  PIN tag_array_ext_ram_wdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1539.560 4.000 1540.160 ;
    END
  END tag_array_ext_ram_wdata[42]
  PIN tag_array_ext_ram_wdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END tag_array_ext_ram_wdata[43]
  PIN tag_array_ext_ram_wdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.040 4.000 1547.640 ;
    END
  END tag_array_ext_ram_wdata[44]
  PIN tag_array_ext_ram_wdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END tag_array_ext_ram_wdata[45]
  PIN tag_array_ext_ram_wdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.840 4.000 1554.440 ;
    END
  END tag_array_ext_ram_wdata[46]
  PIN tag_array_ext_ram_wdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1557.240 4.000 1557.840 ;
    END
  END tag_array_ext_ram_wdata[47]
  PIN tag_array_ext_ram_wdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1560.640 4.000 1561.240 ;
    END
  END tag_array_ext_ram_wdata[48]
  PIN tag_array_ext_ram_wdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.720 4.000 1565.320 ;
    END
  END tag_array_ext_ram_wdata[49]
  PIN tag_array_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1406.280 4.000 1406.880 ;
    END
  END tag_array_ext_ram_wdata[4]
  PIN tag_array_ext_ram_wdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1568.120 4.000 1568.720 ;
    END
  END tag_array_ext_ram_wdata[50]
  PIN tag_array_ext_ram_wdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1571.520 4.000 1572.120 ;
    END
  END tag_array_ext_ram_wdata[51]
  PIN tag_array_ext_ram_wdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.920 4.000 1575.520 ;
    END
  END tag_array_ext_ram_wdata[52]
  PIN tag_array_ext_ram_wdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1578.320 4.000 1578.920 ;
    END
  END tag_array_ext_ram_wdata[53]
  PIN tag_array_ext_ram_wdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1582.400 4.000 1583.000 ;
    END
  END tag_array_ext_ram_wdata[54]
  PIN tag_array_ext_ram_wdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1585.800 4.000 1586.400 ;
    END
  END tag_array_ext_ram_wdata[55]
  PIN tag_array_ext_ram_wdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1589.200 4.000 1589.800 ;
    END
  END tag_array_ext_ram_wdata[56]
  PIN tag_array_ext_ram_wdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1592.600 4.000 1593.200 ;
    END
  END tag_array_ext_ram_wdata[57]
  PIN tag_array_ext_ram_wdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1596.000 4.000 1596.600 ;
    END
  END tag_array_ext_ram_wdata[58]
  PIN tag_array_ext_ram_wdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1599.400 4.000 1600.000 ;
    END
  END tag_array_ext_ram_wdata[59]
  PIN tag_array_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.680 4.000 1410.280 ;
    END
  END tag_array_ext_ram_wdata[5]
  PIN tag_array_ext_ram_wdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1603.480 4.000 1604.080 ;
    END
  END tag_array_ext_ram_wdata[60]
  PIN tag_array_ext_ram_wdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1606.880 4.000 1607.480 ;
    END
  END tag_array_ext_ram_wdata[61]
  PIN tag_array_ext_ram_wdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1610.280 4.000 1610.880 ;
    END
  END tag_array_ext_ram_wdata[62]
  PIN tag_array_ext_ram_wdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1613.680 4.000 1614.280 ;
    END
  END tag_array_ext_ram_wdata[63]
  PIN tag_array_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1413.080 4.000 1413.680 ;
    END
  END tag_array_ext_ram_wdata[6]
  PIN tag_array_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1416.480 4.000 1417.080 ;
    END
  END tag_array_ext_ram_wdata[7]
  PIN tag_array_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1419.880 4.000 1420.480 ;
    END
  END tag_array_ext_ram_wdata[8]
  PIN tag_array_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1423.960 4.000 1424.560 ;
    END
  END tag_array_ext_ram_wdata[9]
  PIN tag_array_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1627.960 4.000 1628.560 ;
    END
  END tag_array_ext_ram_web
  PIN tag_array_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1617.080 4.000 1617.680 ;
    END
  END tag_array_ext_ram_wmask[0]
  PIN tag_array_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1620.480 4.000 1621.080 ;
    END
  END tag_array_ext_ram_wmask[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1765.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1765.520 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1761.800 1765.365 ;
      LAYER met1 ;
        RECT 1.450 1547.240 1767.600 1768.980 ;
        RECT 1.450 1545.740 1767.620 1547.240 ;
        RECT 1.450 1309.240 1767.600 1545.740 ;
        RECT 1.450 1307.400 1767.620 1309.240 ;
        RECT 1.450 4.800 1767.600 1307.400 ;
      LAYER met2 ;
        RECT 1.470 1774.040 7.170 1775.325 ;
        RECT 8.010 1774.040 22.350 1775.325 ;
        RECT 23.190 1774.040 37.990 1775.325 ;
        RECT 38.830 1774.040 53.630 1775.325 ;
        RECT 54.470 1774.040 68.810 1775.325 ;
        RECT 69.650 1774.040 84.450 1775.325 ;
        RECT 85.290 1774.040 100.090 1775.325 ;
        RECT 100.930 1774.040 115.270 1775.325 ;
        RECT 116.110 1774.040 130.910 1775.325 ;
        RECT 131.750 1774.040 146.550 1775.325 ;
        RECT 147.390 1774.040 162.190 1775.325 ;
        RECT 163.030 1774.040 177.370 1775.325 ;
        RECT 178.210 1774.040 193.010 1775.325 ;
        RECT 193.850 1774.040 208.650 1775.325 ;
        RECT 209.490 1774.040 223.830 1775.325 ;
        RECT 224.670 1774.040 239.470 1775.325 ;
        RECT 240.310 1774.040 255.110 1775.325 ;
        RECT 255.950 1774.040 270.750 1775.325 ;
        RECT 271.590 1774.040 285.930 1775.325 ;
        RECT 286.770 1774.040 301.570 1775.325 ;
        RECT 302.410 1774.040 317.210 1775.325 ;
        RECT 318.050 1774.040 332.390 1775.325 ;
        RECT 333.230 1774.040 348.030 1775.325 ;
        RECT 348.870 1774.040 363.670 1775.325 ;
        RECT 364.510 1774.040 379.310 1775.325 ;
        RECT 380.150 1774.040 394.490 1775.325 ;
        RECT 395.330 1774.040 410.130 1775.325 ;
        RECT 410.970 1774.040 425.770 1775.325 ;
        RECT 426.610 1774.040 440.950 1775.325 ;
        RECT 441.790 1774.040 456.590 1775.325 ;
        RECT 457.430 1774.040 472.230 1775.325 ;
        RECT 473.070 1774.040 487.870 1775.325 ;
        RECT 488.710 1774.040 503.050 1775.325 ;
        RECT 503.890 1774.040 518.690 1775.325 ;
        RECT 519.530 1774.040 534.330 1775.325 ;
        RECT 535.170 1774.040 549.510 1775.325 ;
        RECT 550.350 1774.040 565.150 1775.325 ;
        RECT 565.990 1774.040 580.790 1775.325 ;
        RECT 581.630 1774.040 596.430 1775.325 ;
        RECT 597.270 1774.040 611.610 1775.325 ;
        RECT 612.450 1774.040 627.250 1775.325 ;
        RECT 628.090 1774.040 642.890 1775.325 ;
        RECT 643.730 1774.040 658.070 1775.325 ;
        RECT 658.910 1774.040 673.710 1775.325 ;
        RECT 674.550 1774.040 689.350 1775.325 ;
        RECT 690.190 1774.040 704.530 1775.325 ;
        RECT 705.370 1774.040 720.170 1775.325 ;
        RECT 721.010 1774.040 735.810 1775.325 ;
        RECT 736.650 1774.040 751.450 1775.325 ;
        RECT 752.290 1774.040 766.630 1775.325 ;
        RECT 767.470 1774.040 782.270 1775.325 ;
        RECT 783.110 1774.040 797.910 1775.325 ;
        RECT 798.750 1774.040 813.090 1775.325 ;
        RECT 813.930 1774.040 828.730 1775.325 ;
        RECT 829.570 1774.040 844.370 1775.325 ;
        RECT 845.210 1774.040 860.010 1775.325 ;
        RECT 860.850 1774.040 875.190 1775.325 ;
        RECT 876.030 1774.040 890.830 1775.325 ;
        RECT 891.670 1774.040 906.470 1775.325 ;
        RECT 907.310 1774.040 921.650 1775.325 ;
        RECT 922.490 1774.040 937.290 1775.325 ;
        RECT 938.130 1774.040 952.930 1775.325 ;
        RECT 953.770 1774.040 968.570 1775.325 ;
        RECT 969.410 1774.040 983.750 1775.325 ;
        RECT 984.590 1774.040 999.390 1775.325 ;
        RECT 1000.230 1774.040 1015.030 1775.325 ;
        RECT 1015.870 1774.040 1030.210 1775.325 ;
        RECT 1031.050 1774.040 1045.850 1775.325 ;
        RECT 1046.690 1774.040 1061.490 1775.325 ;
        RECT 1062.330 1774.040 1077.130 1775.325 ;
        RECT 1077.970 1774.040 1092.310 1775.325 ;
        RECT 1093.150 1774.040 1107.950 1775.325 ;
        RECT 1108.790 1774.040 1123.590 1775.325 ;
        RECT 1124.430 1774.040 1138.770 1775.325 ;
        RECT 1139.610 1774.040 1154.410 1775.325 ;
        RECT 1155.250 1774.040 1170.050 1775.325 ;
        RECT 1170.890 1774.040 1185.690 1775.325 ;
        RECT 1186.530 1774.040 1200.870 1775.325 ;
        RECT 1201.710 1774.040 1216.510 1775.325 ;
        RECT 1217.350 1774.040 1232.150 1775.325 ;
        RECT 1232.990 1774.040 1247.330 1775.325 ;
        RECT 1248.170 1774.040 1262.970 1775.325 ;
        RECT 1263.810 1774.040 1278.610 1775.325 ;
        RECT 1279.450 1774.040 1293.790 1775.325 ;
        RECT 1294.630 1774.040 1309.430 1775.325 ;
        RECT 1310.270 1774.040 1325.070 1775.325 ;
        RECT 1325.910 1774.040 1340.710 1775.325 ;
        RECT 1341.550 1774.040 1355.890 1775.325 ;
        RECT 1356.730 1774.040 1371.530 1775.325 ;
        RECT 1372.370 1774.040 1387.170 1775.325 ;
        RECT 1388.010 1774.040 1402.350 1775.325 ;
        RECT 1403.190 1774.040 1417.990 1775.325 ;
        RECT 1418.830 1774.040 1433.630 1775.325 ;
        RECT 1434.470 1774.040 1449.270 1775.325 ;
        RECT 1450.110 1774.040 1464.450 1775.325 ;
        RECT 1465.290 1774.040 1480.090 1775.325 ;
        RECT 1480.930 1774.040 1495.730 1775.325 ;
        RECT 1496.570 1774.040 1510.910 1775.325 ;
        RECT 1511.750 1774.040 1526.550 1775.325 ;
        RECT 1527.390 1774.040 1542.190 1775.325 ;
        RECT 1543.030 1774.040 1557.830 1775.325 ;
        RECT 1558.670 1774.040 1573.010 1775.325 ;
        RECT 1573.850 1774.040 1588.650 1775.325 ;
        RECT 1589.490 1774.040 1604.290 1775.325 ;
        RECT 1605.130 1774.040 1619.470 1775.325 ;
        RECT 1620.310 1774.040 1635.110 1775.325 ;
        RECT 1635.950 1774.040 1650.750 1775.325 ;
        RECT 1651.590 1774.040 1666.390 1775.325 ;
        RECT 1667.230 1774.040 1681.570 1775.325 ;
        RECT 1682.410 1774.040 1697.210 1775.325 ;
        RECT 1698.050 1774.040 1712.850 1775.325 ;
        RECT 1713.690 1774.040 1728.030 1775.325 ;
        RECT 1728.870 1774.040 1743.670 1775.325 ;
        RECT 1744.510 1774.040 1759.310 1775.325 ;
        RECT 1760.150 1774.040 1767.600 1775.325 ;
        RECT 1.470 1594.330 1767.600 1774.040 ;
        RECT 1.470 1436.940 1767.620 1594.330 ;
        RECT 1.470 1393.870 1767.600 1436.940 ;
        RECT 1.470 1307.910 1767.620 1393.870 ;
        RECT 1.470 811.820 1767.600 1307.910 ;
        RECT 1.470 742.660 1767.620 811.820 ;
        RECT 1.470 724.570 1767.600 742.660 ;
        RECT 1.470 717.500 1767.620 724.570 ;
        RECT 1.470 716.960 1767.600 717.500 ;
        RECT 1.470 664.800 1767.620 716.960 ;
        RECT 1.470 653.890 1767.600 664.800 ;
        RECT 1.470 596.800 1767.620 653.890 ;
        RECT 1.470 596.090 1767.600 596.800 ;
        RECT 1.470 571.640 1767.620 596.090 ;
        RECT 1.470 541.860 1767.600 571.640 ;
        RECT 1.470 420.830 1767.620 541.860 ;
        RECT 1.470 4.280 1767.600 420.830 ;
        RECT 2.030 1.515 4.410 4.280 ;
        RECT 5.250 1.515 8.090 4.280 ;
        RECT 8.930 1.515 11.770 4.280 ;
        RECT 12.610 1.515 15.450 4.280 ;
        RECT 16.290 1.515 18.670 4.280 ;
        RECT 19.510 1.515 22.350 4.280 ;
        RECT 23.190 1.515 26.030 4.280 ;
        RECT 26.870 1.515 29.710 4.280 ;
        RECT 30.550 1.515 33.390 4.280 ;
        RECT 34.230 1.515 36.610 4.280 ;
        RECT 37.450 1.515 40.290 4.280 ;
        RECT 41.130 1.515 43.970 4.280 ;
        RECT 44.810 1.515 47.650 4.280 ;
        RECT 48.490 1.515 51.330 4.280 ;
        RECT 52.170 1.515 54.550 4.280 ;
        RECT 55.390 1.515 58.230 4.280 ;
        RECT 59.070 1.515 61.910 4.280 ;
        RECT 62.750 1.515 65.590 4.280 ;
        RECT 66.430 1.515 69.270 4.280 ;
        RECT 70.110 1.515 72.490 4.280 ;
        RECT 73.330 1.515 76.170 4.280 ;
        RECT 77.010 1.515 79.850 4.280 ;
        RECT 80.690 1.515 83.530 4.280 ;
        RECT 84.370 1.515 87.210 4.280 ;
        RECT 88.050 1.515 90.430 4.280 ;
        RECT 91.270 1.515 94.110 4.280 ;
        RECT 94.950 1.515 97.790 4.280 ;
        RECT 98.630 1.515 101.470 4.280 ;
        RECT 102.310 1.515 105.150 4.280 ;
        RECT 105.990 1.515 108.370 4.280 ;
        RECT 109.210 1.515 112.050 4.280 ;
        RECT 112.890 1.515 115.730 4.280 ;
        RECT 116.570 1.515 119.410 4.280 ;
        RECT 120.250 1.515 123.090 4.280 ;
        RECT 123.930 1.515 126.310 4.280 ;
        RECT 127.150 1.515 129.990 4.280 ;
        RECT 130.830 1.515 133.670 4.280 ;
        RECT 134.510 1.515 137.350 4.280 ;
        RECT 138.190 1.515 141.030 4.280 ;
        RECT 141.870 1.515 144.250 4.280 ;
        RECT 145.090 1.515 147.930 4.280 ;
        RECT 148.770 1.515 151.610 4.280 ;
        RECT 152.450 1.515 155.290 4.280 ;
        RECT 156.130 1.515 158.510 4.280 ;
        RECT 159.350 1.515 162.190 4.280 ;
        RECT 163.030 1.515 165.870 4.280 ;
        RECT 166.710 1.515 169.550 4.280 ;
        RECT 170.390 1.515 173.230 4.280 ;
        RECT 174.070 1.515 176.450 4.280 ;
        RECT 177.290 1.515 180.130 4.280 ;
        RECT 180.970 1.515 183.810 4.280 ;
        RECT 184.650 1.515 187.490 4.280 ;
        RECT 188.330 1.515 191.170 4.280 ;
        RECT 192.010 1.515 194.390 4.280 ;
        RECT 195.230 1.515 198.070 4.280 ;
        RECT 198.910 1.515 201.750 4.280 ;
        RECT 202.590 1.515 205.430 4.280 ;
        RECT 206.270 1.515 209.110 4.280 ;
        RECT 209.950 1.515 212.330 4.280 ;
        RECT 213.170 1.515 216.010 4.280 ;
        RECT 216.850 1.515 219.690 4.280 ;
        RECT 220.530 1.515 223.370 4.280 ;
        RECT 224.210 1.515 227.050 4.280 ;
        RECT 227.890 1.515 230.270 4.280 ;
        RECT 231.110 1.515 233.950 4.280 ;
        RECT 234.790 1.515 237.630 4.280 ;
        RECT 238.470 1.515 241.310 4.280 ;
        RECT 242.150 1.515 244.990 4.280 ;
        RECT 245.830 1.515 248.210 4.280 ;
        RECT 249.050 1.515 251.890 4.280 ;
        RECT 252.730 1.515 255.570 4.280 ;
        RECT 256.410 1.515 259.250 4.280 ;
        RECT 260.090 1.515 262.930 4.280 ;
        RECT 263.770 1.515 266.150 4.280 ;
        RECT 266.990 1.515 269.830 4.280 ;
        RECT 270.670 1.515 273.510 4.280 ;
        RECT 274.350 1.515 277.190 4.280 ;
        RECT 278.030 1.515 280.870 4.280 ;
        RECT 281.710 1.515 284.090 4.280 ;
        RECT 284.930 1.515 287.770 4.280 ;
        RECT 288.610 1.515 291.450 4.280 ;
        RECT 292.290 1.515 295.130 4.280 ;
        RECT 295.970 1.515 298.350 4.280 ;
        RECT 299.190 1.515 302.030 4.280 ;
        RECT 302.870 1.515 305.710 4.280 ;
        RECT 306.550 1.515 309.390 4.280 ;
        RECT 310.230 1.515 313.070 4.280 ;
        RECT 313.910 1.515 316.290 4.280 ;
        RECT 317.130 1.515 319.970 4.280 ;
        RECT 320.810 1.515 323.650 4.280 ;
        RECT 324.490 1.515 327.330 4.280 ;
        RECT 328.170 1.515 331.010 4.280 ;
        RECT 331.850 1.515 334.230 4.280 ;
        RECT 335.070 1.515 337.910 4.280 ;
        RECT 338.750 1.515 341.590 4.280 ;
        RECT 342.430 1.515 345.270 4.280 ;
        RECT 346.110 1.515 348.950 4.280 ;
        RECT 349.790 1.515 352.170 4.280 ;
        RECT 353.010 1.515 355.850 4.280 ;
        RECT 356.690 1.515 359.530 4.280 ;
        RECT 360.370 1.515 363.210 4.280 ;
        RECT 364.050 1.515 366.890 4.280 ;
        RECT 367.730 1.515 370.110 4.280 ;
        RECT 370.950 1.515 373.790 4.280 ;
        RECT 374.630 1.515 377.470 4.280 ;
        RECT 378.310 1.515 381.150 4.280 ;
        RECT 381.990 1.515 384.830 4.280 ;
        RECT 385.670 1.515 388.050 4.280 ;
        RECT 388.890 1.515 391.730 4.280 ;
        RECT 392.570 1.515 395.410 4.280 ;
        RECT 396.250 1.515 399.090 4.280 ;
        RECT 399.930 1.515 402.770 4.280 ;
        RECT 403.610 1.515 405.990 4.280 ;
        RECT 406.830 1.515 409.670 4.280 ;
        RECT 410.510 1.515 413.350 4.280 ;
        RECT 414.190 1.515 417.030 4.280 ;
        RECT 417.870 1.515 420.710 4.280 ;
        RECT 421.550 1.515 423.930 4.280 ;
        RECT 424.770 1.515 427.610 4.280 ;
        RECT 428.450 1.515 431.290 4.280 ;
        RECT 432.130 1.515 434.970 4.280 ;
        RECT 435.810 1.515 438.650 4.280 ;
        RECT 439.490 1.515 441.870 4.280 ;
        RECT 442.710 1.515 445.550 4.280 ;
        RECT 446.390 1.515 449.230 4.280 ;
        RECT 450.070 1.515 452.910 4.280 ;
        RECT 453.750 1.515 456.130 4.280 ;
        RECT 456.970 1.515 459.810 4.280 ;
        RECT 460.650 1.515 463.490 4.280 ;
        RECT 464.330 1.515 467.170 4.280 ;
        RECT 468.010 1.515 470.850 4.280 ;
        RECT 471.690 1.515 474.070 4.280 ;
        RECT 474.910 1.515 477.750 4.280 ;
        RECT 478.590 1.515 481.430 4.280 ;
        RECT 482.270 1.515 485.110 4.280 ;
        RECT 485.950 1.515 488.790 4.280 ;
        RECT 489.630 1.515 492.010 4.280 ;
        RECT 492.850 1.515 495.690 4.280 ;
        RECT 496.530 1.515 499.370 4.280 ;
        RECT 500.210 1.515 503.050 4.280 ;
        RECT 503.890 1.515 506.730 4.280 ;
        RECT 507.570 1.515 509.950 4.280 ;
        RECT 510.790 1.515 513.630 4.280 ;
        RECT 514.470 1.515 517.310 4.280 ;
        RECT 518.150 1.515 520.990 4.280 ;
        RECT 521.830 1.515 524.670 4.280 ;
        RECT 525.510 1.515 527.890 4.280 ;
        RECT 528.730 1.515 531.570 4.280 ;
        RECT 532.410 1.515 535.250 4.280 ;
        RECT 536.090 1.515 538.930 4.280 ;
        RECT 539.770 1.515 542.610 4.280 ;
        RECT 543.450 1.515 545.830 4.280 ;
        RECT 546.670 1.515 549.510 4.280 ;
        RECT 550.350 1.515 553.190 4.280 ;
        RECT 554.030 1.515 556.870 4.280 ;
        RECT 557.710 1.515 560.550 4.280 ;
        RECT 561.390 1.515 563.770 4.280 ;
        RECT 564.610 1.515 567.450 4.280 ;
        RECT 568.290 1.515 571.130 4.280 ;
        RECT 571.970 1.515 574.810 4.280 ;
        RECT 575.650 1.515 578.490 4.280 ;
        RECT 579.330 1.515 581.710 4.280 ;
        RECT 582.550 1.515 585.390 4.280 ;
        RECT 586.230 1.515 589.070 4.280 ;
        RECT 589.910 1.515 592.750 4.280 ;
        RECT 593.590 1.515 595.970 4.280 ;
        RECT 596.810 1.515 599.650 4.280 ;
        RECT 600.490 1.515 603.330 4.280 ;
        RECT 604.170 1.515 607.010 4.280 ;
        RECT 607.850 1.515 610.690 4.280 ;
        RECT 611.530 1.515 613.910 4.280 ;
        RECT 614.750 1.515 617.590 4.280 ;
        RECT 618.430 1.515 621.270 4.280 ;
        RECT 622.110 1.515 624.950 4.280 ;
        RECT 625.790 1.515 628.630 4.280 ;
        RECT 629.470 1.515 631.850 4.280 ;
        RECT 632.690 1.515 635.530 4.280 ;
        RECT 636.370 1.515 639.210 4.280 ;
        RECT 640.050 1.515 642.890 4.280 ;
        RECT 643.730 1.515 646.570 4.280 ;
        RECT 647.410 1.515 649.790 4.280 ;
        RECT 650.630 1.515 653.470 4.280 ;
        RECT 654.310 1.515 657.150 4.280 ;
        RECT 657.990 1.515 660.830 4.280 ;
        RECT 661.670 1.515 664.510 4.280 ;
        RECT 665.350 1.515 667.730 4.280 ;
        RECT 668.570 1.515 671.410 4.280 ;
        RECT 672.250 1.515 675.090 4.280 ;
        RECT 675.930 1.515 678.770 4.280 ;
        RECT 679.610 1.515 682.450 4.280 ;
        RECT 683.290 1.515 685.670 4.280 ;
        RECT 686.510 1.515 689.350 4.280 ;
        RECT 690.190 1.515 693.030 4.280 ;
        RECT 693.870 1.515 696.710 4.280 ;
        RECT 697.550 1.515 700.390 4.280 ;
        RECT 701.230 1.515 703.610 4.280 ;
        RECT 704.450 1.515 707.290 4.280 ;
        RECT 708.130 1.515 710.970 4.280 ;
        RECT 711.810 1.515 714.650 4.280 ;
        RECT 715.490 1.515 718.330 4.280 ;
        RECT 719.170 1.515 721.550 4.280 ;
        RECT 722.390 1.515 725.230 4.280 ;
        RECT 726.070 1.515 728.910 4.280 ;
        RECT 729.750 1.515 732.590 4.280 ;
        RECT 733.430 1.515 736.270 4.280 ;
        RECT 737.110 1.515 739.490 4.280 ;
        RECT 740.330 1.515 743.170 4.280 ;
        RECT 744.010 1.515 746.850 4.280 ;
        RECT 747.690 1.515 750.530 4.280 ;
        RECT 751.370 1.515 753.750 4.280 ;
        RECT 754.590 1.515 757.430 4.280 ;
        RECT 758.270 1.515 761.110 4.280 ;
        RECT 761.950 1.515 764.790 4.280 ;
        RECT 765.630 1.515 768.470 4.280 ;
        RECT 769.310 1.515 771.690 4.280 ;
        RECT 772.530 1.515 775.370 4.280 ;
        RECT 776.210 1.515 779.050 4.280 ;
        RECT 779.890 1.515 782.730 4.280 ;
        RECT 783.570 1.515 786.410 4.280 ;
        RECT 787.250 1.515 789.630 4.280 ;
        RECT 790.470 1.515 793.310 4.280 ;
        RECT 794.150 1.515 796.990 4.280 ;
        RECT 797.830 1.515 800.670 4.280 ;
        RECT 801.510 1.515 804.350 4.280 ;
        RECT 805.190 1.515 807.570 4.280 ;
        RECT 808.410 1.515 811.250 4.280 ;
        RECT 812.090 1.515 814.930 4.280 ;
        RECT 815.770 1.515 818.610 4.280 ;
        RECT 819.450 1.515 822.290 4.280 ;
        RECT 823.130 1.515 825.510 4.280 ;
        RECT 826.350 1.515 829.190 4.280 ;
        RECT 830.030 1.515 832.870 4.280 ;
        RECT 833.710 1.515 836.550 4.280 ;
        RECT 837.390 1.515 840.230 4.280 ;
        RECT 841.070 1.515 843.450 4.280 ;
        RECT 844.290 1.515 847.130 4.280 ;
        RECT 847.970 1.515 850.810 4.280 ;
        RECT 851.650 1.515 854.490 4.280 ;
        RECT 855.330 1.515 858.170 4.280 ;
        RECT 859.010 1.515 861.390 4.280 ;
        RECT 862.230 1.515 865.070 4.280 ;
        RECT 865.910 1.515 868.750 4.280 ;
        RECT 869.590 1.515 872.430 4.280 ;
        RECT 873.270 1.515 876.110 4.280 ;
        RECT 876.950 1.515 879.330 4.280 ;
        RECT 880.170 1.515 883.010 4.280 ;
        RECT 883.850 1.515 886.690 4.280 ;
        RECT 887.530 1.515 890.370 4.280 ;
        RECT 891.210 1.515 893.590 4.280 ;
        RECT 894.430 1.515 897.270 4.280 ;
        RECT 898.110 1.515 900.950 4.280 ;
        RECT 901.790 1.515 904.630 4.280 ;
        RECT 905.470 1.515 908.310 4.280 ;
        RECT 909.150 1.515 911.530 4.280 ;
        RECT 912.370 1.515 915.210 4.280 ;
        RECT 916.050 1.515 918.890 4.280 ;
        RECT 919.730 1.515 922.570 4.280 ;
        RECT 923.410 1.515 926.250 4.280 ;
        RECT 927.090 1.515 929.470 4.280 ;
        RECT 930.310 1.515 933.150 4.280 ;
        RECT 933.990 1.515 936.830 4.280 ;
        RECT 937.670 1.515 940.510 4.280 ;
        RECT 941.350 1.515 944.190 4.280 ;
        RECT 945.030 1.515 947.410 4.280 ;
        RECT 948.250 1.515 951.090 4.280 ;
        RECT 951.930 1.515 954.770 4.280 ;
        RECT 955.610 1.515 958.450 4.280 ;
        RECT 959.290 1.515 962.130 4.280 ;
        RECT 962.970 1.515 965.350 4.280 ;
        RECT 966.190 1.515 969.030 4.280 ;
        RECT 969.870 1.515 972.710 4.280 ;
        RECT 973.550 1.515 976.390 4.280 ;
        RECT 977.230 1.515 980.070 4.280 ;
        RECT 980.910 1.515 983.290 4.280 ;
        RECT 984.130 1.515 986.970 4.280 ;
        RECT 987.810 1.515 990.650 4.280 ;
        RECT 991.490 1.515 994.330 4.280 ;
        RECT 995.170 1.515 998.010 4.280 ;
        RECT 998.850 1.515 1001.230 4.280 ;
        RECT 1002.070 1.515 1004.910 4.280 ;
        RECT 1005.750 1.515 1008.590 4.280 ;
        RECT 1009.430 1.515 1012.270 4.280 ;
        RECT 1013.110 1.515 1015.950 4.280 ;
        RECT 1016.790 1.515 1019.170 4.280 ;
        RECT 1020.010 1.515 1022.850 4.280 ;
        RECT 1023.690 1.515 1026.530 4.280 ;
        RECT 1027.370 1.515 1030.210 4.280 ;
        RECT 1031.050 1.515 1033.430 4.280 ;
        RECT 1034.270 1.515 1037.110 4.280 ;
        RECT 1037.950 1.515 1040.790 4.280 ;
        RECT 1041.630 1.515 1044.470 4.280 ;
        RECT 1045.310 1.515 1048.150 4.280 ;
        RECT 1048.990 1.515 1051.370 4.280 ;
        RECT 1052.210 1.515 1055.050 4.280 ;
        RECT 1055.890 1.515 1058.730 4.280 ;
        RECT 1059.570 1.515 1062.410 4.280 ;
        RECT 1063.250 1.515 1066.090 4.280 ;
        RECT 1066.930 1.515 1069.310 4.280 ;
        RECT 1070.150 1.515 1072.990 4.280 ;
        RECT 1073.830 1.515 1076.670 4.280 ;
        RECT 1077.510 1.515 1080.350 4.280 ;
        RECT 1081.190 1.515 1084.030 4.280 ;
        RECT 1084.870 1.515 1087.250 4.280 ;
        RECT 1088.090 1.515 1090.930 4.280 ;
        RECT 1091.770 1.515 1094.610 4.280 ;
        RECT 1095.450 1.515 1098.290 4.280 ;
        RECT 1099.130 1.515 1101.970 4.280 ;
        RECT 1102.810 1.515 1105.190 4.280 ;
        RECT 1106.030 1.515 1108.870 4.280 ;
        RECT 1109.710 1.515 1112.550 4.280 ;
        RECT 1113.390 1.515 1116.230 4.280 ;
        RECT 1117.070 1.515 1119.910 4.280 ;
        RECT 1120.750 1.515 1123.130 4.280 ;
        RECT 1123.970 1.515 1126.810 4.280 ;
        RECT 1127.650 1.515 1130.490 4.280 ;
        RECT 1131.330 1.515 1134.170 4.280 ;
        RECT 1135.010 1.515 1137.850 4.280 ;
        RECT 1138.690 1.515 1141.070 4.280 ;
        RECT 1141.910 1.515 1144.750 4.280 ;
        RECT 1145.590 1.515 1148.430 4.280 ;
        RECT 1149.270 1.515 1152.110 4.280 ;
        RECT 1152.950 1.515 1155.790 4.280 ;
        RECT 1156.630 1.515 1159.010 4.280 ;
        RECT 1159.850 1.515 1162.690 4.280 ;
        RECT 1163.530 1.515 1166.370 4.280 ;
        RECT 1167.210 1.515 1170.050 4.280 ;
        RECT 1170.890 1.515 1173.730 4.280 ;
        RECT 1174.570 1.515 1176.950 4.280 ;
        RECT 1177.790 1.515 1180.630 4.280 ;
        RECT 1181.470 1.515 1184.310 4.280 ;
        RECT 1185.150 1.515 1187.990 4.280 ;
        RECT 1188.830 1.515 1191.210 4.280 ;
        RECT 1192.050 1.515 1194.890 4.280 ;
        RECT 1195.730 1.515 1198.570 4.280 ;
        RECT 1199.410 1.515 1202.250 4.280 ;
        RECT 1203.090 1.515 1205.930 4.280 ;
        RECT 1206.770 1.515 1209.150 4.280 ;
        RECT 1209.990 1.515 1212.830 4.280 ;
        RECT 1213.670 1.515 1216.510 4.280 ;
        RECT 1217.350 1.515 1220.190 4.280 ;
        RECT 1221.030 1.515 1223.870 4.280 ;
        RECT 1224.710 1.515 1227.090 4.280 ;
        RECT 1227.930 1.515 1230.770 4.280 ;
        RECT 1231.610 1.515 1234.450 4.280 ;
        RECT 1235.290 1.515 1238.130 4.280 ;
        RECT 1238.970 1.515 1241.810 4.280 ;
        RECT 1242.650 1.515 1245.030 4.280 ;
        RECT 1245.870 1.515 1248.710 4.280 ;
        RECT 1249.550 1.515 1252.390 4.280 ;
        RECT 1253.230 1.515 1256.070 4.280 ;
        RECT 1256.910 1.515 1259.750 4.280 ;
        RECT 1260.590 1.515 1262.970 4.280 ;
        RECT 1263.810 1.515 1266.650 4.280 ;
        RECT 1267.490 1.515 1270.330 4.280 ;
        RECT 1271.170 1.515 1274.010 4.280 ;
        RECT 1274.850 1.515 1277.690 4.280 ;
        RECT 1278.530 1.515 1280.910 4.280 ;
        RECT 1281.750 1.515 1284.590 4.280 ;
        RECT 1285.430 1.515 1288.270 4.280 ;
        RECT 1289.110 1.515 1291.950 4.280 ;
        RECT 1292.790 1.515 1295.630 4.280 ;
        RECT 1296.470 1.515 1298.850 4.280 ;
        RECT 1299.690 1.515 1302.530 4.280 ;
        RECT 1303.370 1.515 1306.210 4.280 ;
        RECT 1307.050 1.515 1309.890 4.280 ;
        RECT 1310.730 1.515 1313.570 4.280 ;
        RECT 1314.410 1.515 1316.790 4.280 ;
        RECT 1317.630 1.515 1320.470 4.280 ;
        RECT 1321.310 1.515 1324.150 4.280 ;
        RECT 1324.990 1.515 1327.830 4.280 ;
        RECT 1328.670 1.515 1331.050 4.280 ;
        RECT 1331.890 1.515 1334.730 4.280 ;
        RECT 1335.570 1.515 1338.410 4.280 ;
        RECT 1339.250 1.515 1342.090 4.280 ;
        RECT 1342.930 1.515 1345.770 4.280 ;
        RECT 1346.610 1.515 1348.990 4.280 ;
        RECT 1349.830 1.515 1352.670 4.280 ;
        RECT 1353.510 1.515 1356.350 4.280 ;
        RECT 1357.190 1.515 1360.030 4.280 ;
        RECT 1360.870 1.515 1363.710 4.280 ;
        RECT 1364.550 1.515 1366.930 4.280 ;
        RECT 1367.770 1.515 1370.610 4.280 ;
        RECT 1371.450 1.515 1374.290 4.280 ;
        RECT 1375.130 1.515 1377.970 4.280 ;
        RECT 1378.810 1.515 1381.650 4.280 ;
        RECT 1382.490 1.515 1384.870 4.280 ;
        RECT 1385.710 1.515 1388.550 4.280 ;
        RECT 1389.390 1.515 1392.230 4.280 ;
        RECT 1393.070 1.515 1395.910 4.280 ;
        RECT 1396.750 1.515 1399.590 4.280 ;
        RECT 1400.430 1.515 1402.810 4.280 ;
        RECT 1403.650 1.515 1406.490 4.280 ;
        RECT 1407.330 1.515 1410.170 4.280 ;
        RECT 1411.010 1.515 1413.850 4.280 ;
        RECT 1414.690 1.515 1417.530 4.280 ;
        RECT 1418.370 1.515 1420.750 4.280 ;
        RECT 1421.590 1.515 1424.430 4.280 ;
        RECT 1425.270 1.515 1428.110 4.280 ;
        RECT 1428.950 1.515 1431.790 4.280 ;
        RECT 1432.630 1.515 1435.470 4.280 ;
        RECT 1436.310 1.515 1438.690 4.280 ;
        RECT 1439.530 1.515 1442.370 4.280 ;
        RECT 1443.210 1.515 1446.050 4.280 ;
        RECT 1446.890 1.515 1449.730 4.280 ;
        RECT 1450.570 1.515 1453.410 4.280 ;
        RECT 1454.250 1.515 1456.630 4.280 ;
        RECT 1457.470 1.515 1460.310 4.280 ;
        RECT 1461.150 1.515 1463.990 4.280 ;
        RECT 1464.830 1.515 1467.670 4.280 ;
        RECT 1468.510 1.515 1471.350 4.280 ;
        RECT 1472.190 1.515 1474.570 4.280 ;
        RECT 1475.410 1.515 1478.250 4.280 ;
        RECT 1479.090 1.515 1481.930 4.280 ;
        RECT 1482.770 1.515 1485.610 4.280 ;
        RECT 1486.450 1.515 1488.830 4.280 ;
        RECT 1489.670 1.515 1492.510 4.280 ;
        RECT 1493.350 1.515 1496.190 4.280 ;
        RECT 1497.030 1.515 1499.870 4.280 ;
        RECT 1500.710 1.515 1503.550 4.280 ;
        RECT 1504.390 1.515 1506.770 4.280 ;
        RECT 1507.610 1.515 1510.450 4.280 ;
        RECT 1511.290 1.515 1514.130 4.280 ;
        RECT 1514.970 1.515 1517.810 4.280 ;
        RECT 1518.650 1.515 1521.490 4.280 ;
        RECT 1522.330 1.515 1524.710 4.280 ;
        RECT 1525.550 1.515 1528.390 4.280 ;
        RECT 1529.230 1.515 1532.070 4.280 ;
        RECT 1532.910 1.515 1535.750 4.280 ;
        RECT 1536.590 1.515 1539.430 4.280 ;
        RECT 1540.270 1.515 1542.650 4.280 ;
        RECT 1543.490 1.515 1546.330 4.280 ;
        RECT 1547.170 1.515 1550.010 4.280 ;
        RECT 1550.850 1.515 1553.690 4.280 ;
        RECT 1554.530 1.515 1557.370 4.280 ;
        RECT 1558.210 1.515 1560.590 4.280 ;
        RECT 1561.430 1.515 1564.270 4.280 ;
        RECT 1565.110 1.515 1567.950 4.280 ;
        RECT 1568.790 1.515 1571.630 4.280 ;
        RECT 1572.470 1.515 1575.310 4.280 ;
        RECT 1576.150 1.515 1578.530 4.280 ;
        RECT 1579.370 1.515 1582.210 4.280 ;
        RECT 1583.050 1.515 1585.890 4.280 ;
        RECT 1586.730 1.515 1589.570 4.280 ;
        RECT 1590.410 1.515 1593.250 4.280 ;
        RECT 1594.090 1.515 1596.470 4.280 ;
        RECT 1597.310 1.515 1600.150 4.280 ;
        RECT 1600.990 1.515 1603.830 4.280 ;
        RECT 1604.670 1.515 1607.510 4.280 ;
        RECT 1608.350 1.515 1611.190 4.280 ;
        RECT 1612.030 1.515 1614.410 4.280 ;
        RECT 1615.250 1.515 1618.090 4.280 ;
        RECT 1618.930 1.515 1621.770 4.280 ;
        RECT 1622.610 1.515 1625.450 4.280 ;
        RECT 1626.290 1.515 1628.670 4.280 ;
        RECT 1629.510 1.515 1632.350 4.280 ;
        RECT 1633.190 1.515 1636.030 4.280 ;
        RECT 1636.870 1.515 1639.710 4.280 ;
        RECT 1640.550 1.515 1643.390 4.280 ;
        RECT 1644.230 1.515 1646.610 4.280 ;
        RECT 1647.450 1.515 1650.290 4.280 ;
        RECT 1651.130 1.515 1653.970 4.280 ;
        RECT 1654.810 1.515 1657.650 4.280 ;
        RECT 1658.490 1.515 1661.330 4.280 ;
        RECT 1662.170 1.515 1664.550 4.280 ;
        RECT 1665.390 1.515 1668.230 4.280 ;
        RECT 1669.070 1.515 1671.910 4.280 ;
        RECT 1672.750 1.515 1675.590 4.280 ;
        RECT 1676.430 1.515 1679.270 4.280 ;
        RECT 1680.110 1.515 1682.490 4.280 ;
        RECT 1683.330 1.515 1686.170 4.280 ;
        RECT 1687.010 1.515 1689.850 4.280 ;
        RECT 1690.690 1.515 1693.530 4.280 ;
        RECT 1694.370 1.515 1697.210 4.280 ;
        RECT 1698.050 1.515 1700.430 4.280 ;
        RECT 1701.270 1.515 1704.110 4.280 ;
        RECT 1704.950 1.515 1707.790 4.280 ;
        RECT 1708.630 1.515 1711.470 4.280 ;
        RECT 1712.310 1.515 1715.150 4.280 ;
        RECT 1715.990 1.515 1718.370 4.280 ;
        RECT 1719.210 1.515 1722.050 4.280 ;
        RECT 1722.890 1.515 1725.730 4.280 ;
        RECT 1726.570 1.515 1729.410 4.280 ;
        RECT 1730.250 1.515 1733.090 4.280 ;
        RECT 1733.930 1.515 1736.310 4.280 ;
        RECT 1737.150 1.515 1739.990 4.280 ;
        RECT 1740.830 1.515 1743.670 4.280 ;
        RECT 1744.510 1.515 1747.350 4.280 ;
        RECT 1748.190 1.515 1751.030 4.280 ;
        RECT 1751.870 1.515 1754.250 4.280 ;
        RECT 1755.090 1.515 1757.930 4.280 ;
        RECT 1758.770 1.515 1761.610 4.280 ;
        RECT 1762.450 1.515 1765.290 4.280 ;
        RECT 1766.130 1.515 1767.600 4.280 ;
      LAYER met3 ;
        RECT 4.400 1775.120 1763.200 1775.305 ;
        RECT 1.445 1774.440 1763.200 1775.120 ;
        RECT 1.445 1773.120 1767.255 1774.440 ;
        RECT 4.400 1771.720 1767.255 1773.120 ;
        RECT 1.445 1770.400 1767.255 1771.720 ;
        RECT 1.445 1769.720 1763.200 1770.400 ;
        RECT 4.400 1769.000 1763.200 1769.720 ;
        RECT 4.400 1768.320 1767.255 1769.000 ;
        RECT 1.445 1766.320 1767.255 1768.320 ;
        RECT 4.400 1764.960 1767.255 1766.320 ;
        RECT 4.400 1764.920 1763.200 1764.960 ;
        RECT 1.445 1763.560 1763.200 1764.920 ;
        RECT 1.445 1762.920 1767.255 1763.560 ;
        RECT 4.400 1761.520 1767.255 1762.920 ;
        RECT 1.445 1759.520 1767.255 1761.520 ;
        RECT 1.445 1758.840 1763.200 1759.520 ;
        RECT 4.400 1758.120 1763.200 1758.840 ;
        RECT 4.400 1757.440 1767.255 1758.120 ;
        RECT 1.445 1755.440 1767.255 1757.440 ;
        RECT 4.400 1754.080 1767.255 1755.440 ;
        RECT 4.400 1754.040 1763.200 1754.080 ;
        RECT 1.445 1752.680 1763.200 1754.040 ;
        RECT 1.445 1752.040 1767.255 1752.680 ;
        RECT 4.400 1750.640 1767.255 1752.040 ;
        RECT 1.445 1748.640 1767.255 1750.640 ;
        RECT 4.400 1747.240 1763.200 1748.640 ;
        RECT 1.445 1745.240 1767.255 1747.240 ;
        RECT 4.400 1743.840 1767.255 1745.240 ;
        RECT 1.445 1743.200 1767.255 1743.840 ;
        RECT 1.445 1741.840 1763.200 1743.200 ;
        RECT 4.400 1741.800 1763.200 1741.840 ;
        RECT 4.400 1740.440 1767.255 1741.800 ;
        RECT 1.445 1737.760 1767.255 1740.440 ;
        RECT 4.400 1736.360 1763.200 1737.760 ;
        RECT 1.445 1734.360 1767.255 1736.360 ;
        RECT 4.400 1732.960 1767.255 1734.360 ;
        RECT 1.445 1732.320 1767.255 1732.960 ;
        RECT 1.445 1730.960 1763.200 1732.320 ;
        RECT 4.400 1730.920 1763.200 1730.960 ;
        RECT 4.400 1729.560 1767.255 1730.920 ;
        RECT 1.445 1727.560 1767.255 1729.560 ;
        RECT 4.400 1726.880 1767.255 1727.560 ;
        RECT 4.400 1726.160 1763.200 1726.880 ;
        RECT 1.445 1725.480 1763.200 1726.160 ;
        RECT 1.445 1724.160 1767.255 1725.480 ;
        RECT 4.400 1722.760 1767.255 1724.160 ;
        RECT 1.445 1721.440 1767.255 1722.760 ;
        RECT 1.445 1720.080 1763.200 1721.440 ;
        RECT 4.400 1720.040 1763.200 1720.080 ;
        RECT 4.400 1718.680 1767.255 1720.040 ;
        RECT 1.445 1716.680 1767.255 1718.680 ;
        RECT 4.400 1716.000 1767.255 1716.680 ;
        RECT 4.400 1715.280 1763.200 1716.000 ;
        RECT 1.445 1714.600 1763.200 1715.280 ;
        RECT 1.445 1713.280 1767.255 1714.600 ;
        RECT 4.400 1711.880 1767.255 1713.280 ;
        RECT 1.445 1710.560 1767.255 1711.880 ;
        RECT 1.445 1709.880 1763.200 1710.560 ;
        RECT 4.400 1709.160 1763.200 1709.880 ;
        RECT 4.400 1708.480 1767.255 1709.160 ;
        RECT 1.445 1706.480 1767.255 1708.480 ;
        RECT 4.400 1705.120 1767.255 1706.480 ;
        RECT 4.400 1705.080 1763.200 1705.120 ;
        RECT 1.445 1703.720 1763.200 1705.080 ;
        RECT 1.445 1703.080 1767.255 1703.720 ;
        RECT 4.400 1701.680 1767.255 1703.080 ;
        RECT 1.445 1699.680 1767.255 1701.680 ;
        RECT 1.445 1699.000 1763.200 1699.680 ;
        RECT 4.400 1698.280 1763.200 1699.000 ;
        RECT 4.400 1697.600 1767.255 1698.280 ;
        RECT 1.445 1695.600 1767.255 1697.600 ;
        RECT 4.400 1694.240 1767.255 1695.600 ;
        RECT 4.400 1694.200 1763.200 1694.240 ;
        RECT 1.445 1692.840 1763.200 1694.200 ;
        RECT 1.445 1692.200 1767.255 1692.840 ;
        RECT 4.400 1690.800 1767.255 1692.200 ;
        RECT 1.445 1688.800 1767.255 1690.800 ;
        RECT 4.400 1687.400 1763.200 1688.800 ;
        RECT 1.445 1685.400 1767.255 1687.400 ;
        RECT 4.400 1684.000 1767.255 1685.400 ;
        RECT 1.445 1683.360 1767.255 1684.000 ;
        RECT 1.445 1682.000 1763.200 1683.360 ;
        RECT 4.400 1681.960 1763.200 1682.000 ;
        RECT 4.400 1680.600 1767.255 1681.960 ;
        RECT 1.445 1677.920 1767.255 1680.600 ;
        RECT 4.400 1676.520 1763.200 1677.920 ;
        RECT 1.445 1674.520 1767.255 1676.520 ;
        RECT 4.400 1673.120 1767.255 1674.520 ;
        RECT 1.445 1672.480 1767.255 1673.120 ;
        RECT 1.445 1671.120 1763.200 1672.480 ;
        RECT 4.400 1671.080 1763.200 1671.120 ;
        RECT 4.400 1669.720 1767.255 1671.080 ;
        RECT 1.445 1667.720 1767.255 1669.720 ;
        RECT 4.400 1667.040 1767.255 1667.720 ;
        RECT 4.400 1666.320 1763.200 1667.040 ;
        RECT 1.445 1665.640 1763.200 1666.320 ;
        RECT 1.445 1664.320 1767.255 1665.640 ;
        RECT 4.400 1662.920 1767.255 1664.320 ;
        RECT 1.445 1661.600 1767.255 1662.920 ;
        RECT 1.445 1660.240 1763.200 1661.600 ;
        RECT 4.400 1660.200 1763.200 1660.240 ;
        RECT 4.400 1658.840 1767.255 1660.200 ;
        RECT 1.445 1656.840 1767.255 1658.840 ;
        RECT 4.400 1656.160 1767.255 1656.840 ;
        RECT 4.400 1655.440 1763.200 1656.160 ;
        RECT 1.445 1654.760 1763.200 1655.440 ;
        RECT 1.445 1653.440 1767.255 1654.760 ;
        RECT 4.400 1652.040 1767.255 1653.440 ;
        RECT 1.445 1650.720 1767.255 1652.040 ;
        RECT 1.445 1650.040 1763.200 1650.720 ;
        RECT 4.400 1649.320 1763.200 1650.040 ;
        RECT 4.400 1648.640 1767.255 1649.320 ;
        RECT 1.445 1646.640 1767.255 1648.640 ;
        RECT 4.400 1645.280 1767.255 1646.640 ;
        RECT 4.400 1645.240 1763.200 1645.280 ;
        RECT 1.445 1643.880 1763.200 1645.240 ;
        RECT 1.445 1643.240 1767.255 1643.880 ;
        RECT 4.400 1641.840 1767.255 1643.240 ;
        RECT 1.445 1639.840 1767.255 1641.840 ;
        RECT 1.445 1639.160 1763.200 1639.840 ;
        RECT 4.400 1638.440 1763.200 1639.160 ;
        RECT 4.400 1637.760 1767.255 1638.440 ;
        RECT 1.445 1635.760 1767.255 1637.760 ;
        RECT 4.400 1634.400 1767.255 1635.760 ;
        RECT 4.400 1634.360 1763.200 1634.400 ;
        RECT 1.445 1633.000 1763.200 1634.360 ;
        RECT 1.445 1632.360 1767.255 1633.000 ;
        RECT 4.400 1630.960 1767.255 1632.360 ;
        RECT 1.445 1628.960 1767.255 1630.960 ;
        RECT 4.400 1627.560 1763.200 1628.960 ;
        RECT 1.445 1625.560 1767.255 1627.560 ;
        RECT 4.400 1624.160 1767.255 1625.560 ;
        RECT 1.445 1623.520 1767.255 1624.160 ;
        RECT 1.445 1622.120 1763.200 1623.520 ;
        RECT 1.445 1621.480 1767.255 1622.120 ;
        RECT 4.400 1620.080 1767.255 1621.480 ;
        RECT 1.445 1618.080 1767.255 1620.080 ;
        RECT 4.400 1616.680 1763.200 1618.080 ;
        RECT 1.445 1614.680 1767.255 1616.680 ;
        RECT 4.400 1613.280 1767.255 1614.680 ;
        RECT 1.445 1612.640 1767.255 1613.280 ;
        RECT 1.445 1611.280 1763.200 1612.640 ;
        RECT 4.400 1611.240 1763.200 1611.280 ;
        RECT 4.400 1609.880 1767.255 1611.240 ;
        RECT 1.445 1607.880 1767.255 1609.880 ;
        RECT 4.400 1607.200 1767.255 1607.880 ;
        RECT 4.400 1606.480 1763.200 1607.200 ;
        RECT 1.445 1605.800 1763.200 1606.480 ;
        RECT 1.445 1604.480 1767.255 1605.800 ;
        RECT 4.400 1603.080 1767.255 1604.480 ;
        RECT 1.445 1601.760 1767.255 1603.080 ;
        RECT 1.445 1600.400 1763.200 1601.760 ;
        RECT 4.400 1600.360 1763.200 1600.400 ;
        RECT 4.400 1599.000 1767.255 1600.360 ;
        RECT 1.445 1597.000 1767.255 1599.000 ;
        RECT 4.400 1596.320 1767.255 1597.000 ;
        RECT 4.400 1595.600 1763.200 1596.320 ;
        RECT 1.445 1594.920 1763.200 1595.600 ;
        RECT 1.445 1593.600 1767.255 1594.920 ;
        RECT 4.400 1592.200 1767.255 1593.600 ;
        RECT 1.445 1590.880 1767.255 1592.200 ;
        RECT 1.445 1590.200 1763.200 1590.880 ;
        RECT 4.400 1589.480 1763.200 1590.200 ;
        RECT 4.400 1588.800 1767.255 1589.480 ;
        RECT 1.445 1586.800 1767.255 1588.800 ;
        RECT 4.400 1585.440 1767.255 1586.800 ;
        RECT 4.400 1585.400 1763.200 1585.440 ;
        RECT 1.445 1584.040 1763.200 1585.400 ;
        RECT 1.445 1583.400 1767.255 1584.040 ;
        RECT 4.400 1582.000 1767.255 1583.400 ;
        RECT 1.445 1580.680 1767.255 1582.000 ;
        RECT 1.445 1579.320 1763.200 1580.680 ;
        RECT 4.400 1579.280 1763.200 1579.320 ;
        RECT 4.400 1577.920 1767.255 1579.280 ;
        RECT 1.445 1575.920 1767.255 1577.920 ;
        RECT 4.400 1575.240 1767.255 1575.920 ;
        RECT 4.400 1574.520 1763.200 1575.240 ;
        RECT 1.445 1573.840 1763.200 1574.520 ;
        RECT 1.445 1572.520 1767.255 1573.840 ;
        RECT 4.400 1571.120 1767.255 1572.520 ;
        RECT 1.445 1569.800 1767.255 1571.120 ;
        RECT 1.445 1569.120 1763.200 1569.800 ;
        RECT 4.400 1568.400 1763.200 1569.120 ;
        RECT 4.400 1567.720 1767.255 1568.400 ;
        RECT 1.445 1565.720 1767.255 1567.720 ;
        RECT 4.400 1564.360 1767.255 1565.720 ;
        RECT 4.400 1564.320 1763.200 1564.360 ;
        RECT 1.445 1562.960 1763.200 1564.320 ;
        RECT 1.445 1561.640 1767.255 1562.960 ;
        RECT 4.400 1560.240 1767.255 1561.640 ;
        RECT 1.445 1558.920 1767.255 1560.240 ;
        RECT 1.445 1558.240 1763.200 1558.920 ;
        RECT 4.400 1557.520 1763.200 1558.240 ;
        RECT 4.400 1556.840 1767.255 1557.520 ;
        RECT 1.445 1554.840 1767.255 1556.840 ;
        RECT 4.400 1553.480 1767.255 1554.840 ;
        RECT 4.400 1553.440 1763.200 1553.480 ;
        RECT 1.445 1552.080 1763.200 1553.440 ;
        RECT 1.445 1551.440 1767.255 1552.080 ;
        RECT 4.400 1550.040 1767.255 1551.440 ;
        RECT 1.445 1548.040 1767.255 1550.040 ;
        RECT 4.400 1546.640 1763.200 1548.040 ;
        RECT 1.445 1544.640 1767.255 1546.640 ;
        RECT 4.400 1543.240 1767.255 1544.640 ;
        RECT 1.445 1542.600 1767.255 1543.240 ;
        RECT 1.445 1541.200 1763.200 1542.600 ;
        RECT 1.445 1540.560 1767.255 1541.200 ;
        RECT 4.400 1539.160 1767.255 1540.560 ;
        RECT 1.445 1537.160 1767.255 1539.160 ;
        RECT 4.400 1535.760 1763.200 1537.160 ;
        RECT 1.445 1533.760 1767.255 1535.760 ;
        RECT 4.400 1532.360 1767.255 1533.760 ;
        RECT 1.445 1531.720 1767.255 1532.360 ;
        RECT 1.445 1530.360 1763.200 1531.720 ;
        RECT 4.400 1530.320 1763.200 1530.360 ;
        RECT 4.400 1528.960 1767.255 1530.320 ;
        RECT 1.445 1526.960 1767.255 1528.960 ;
        RECT 4.400 1526.280 1767.255 1526.960 ;
        RECT 4.400 1525.560 1763.200 1526.280 ;
        RECT 1.445 1524.880 1763.200 1525.560 ;
        RECT 1.445 1522.880 1767.255 1524.880 ;
        RECT 4.400 1521.480 1767.255 1522.880 ;
        RECT 1.445 1520.840 1767.255 1521.480 ;
        RECT 1.445 1519.480 1763.200 1520.840 ;
        RECT 4.400 1519.440 1763.200 1519.480 ;
        RECT 4.400 1518.080 1767.255 1519.440 ;
        RECT 1.445 1516.080 1767.255 1518.080 ;
        RECT 4.400 1515.400 1767.255 1516.080 ;
        RECT 4.400 1514.680 1763.200 1515.400 ;
        RECT 1.445 1514.000 1763.200 1514.680 ;
        RECT 1.445 1512.680 1767.255 1514.000 ;
        RECT 4.400 1511.280 1767.255 1512.680 ;
        RECT 1.445 1509.960 1767.255 1511.280 ;
        RECT 1.445 1509.280 1763.200 1509.960 ;
        RECT 4.400 1508.560 1763.200 1509.280 ;
        RECT 4.400 1507.880 1767.255 1508.560 ;
        RECT 1.445 1505.880 1767.255 1507.880 ;
        RECT 4.400 1504.520 1767.255 1505.880 ;
        RECT 4.400 1504.480 1763.200 1504.520 ;
        RECT 1.445 1503.120 1763.200 1504.480 ;
        RECT 1.445 1501.800 1767.255 1503.120 ;
        RECT 4.400 1500.400 1767.255 1501.800 ;
        RECT 1.445 1499.080 1767.255 1500.400 ;
        RECT 1.445 1498.400 1763.200 1499.080 ;
        RECT 4.400 1497.680 1763.200 1498.400 ;
        RECT 4.400 1497.000 1767.255 1497.680 ;
        RECT 1.445 1495.000 1767.255 1497.000 ;
        RECT 4.400 1493.640 1767.255 1495.000 ;
        RECT 4.400 1493.600 1763.200 1493.640 ;
        RECT 1.445 1492.240 1763.200 1493.600 ;
        RECT 1.445 1491.600 1767.255 1492.240 ;
        RECT 4.400 1490.200 1767.255 1491.600 ;
        RECT 1.445 1488.200 1767.255 1490.200 ;
        RECT 4.400 1486.800 1763.200 1488.200 ;
        RECT 1.445 1484.800 1767.255 1486.800 ;
        RECT 4.400 1483.400 1767.255 1484.800 ;
        RECT 1.445 1482.760 1767.255 1483.400 ;
        RECT 1.445 1481.360 1763.200 1482.760 ;
        RECT 1.445 1480.720 1767.255 1481.360 ;
        RECT 4.400 1479.320 1767.255 1480.720 ;
        RECT 1.445 1477.320 1767.255 1479.320 ;
        RECT 4.400 1475.920 1763.200 1477.320 ;
        RECT 1.445 1473.920 1767.255 1475.920 ;
        RECT 4.400 1472.520 1767.255 1473.920 ;
        RECT 1.445 1471.880 1767.255 1472.520 ;
        RECT 1.445 1470.520 1763.200 1471.880 ;
        RECT 4.400 1470.480 1763.200 1470.520 ;
        RECT 4.400 1469.120 1767.255 1470.480 ;
        RECT 1.445 1467.120 1767.255 1469.120 ;
        RECT 4.400 1466.440 1767.255 1467.120 ;
        RECT 4.400 1465.720 1763.200 1466.440 ;
        RECT 1.445 1465.040 1763.200 1465.720 ;
        RECT 1.445 1463.040 1767.255 1465.040 ;
        RECT 4.400 1461.640 1767.255 1463.040 ;
        RECT 1.445 1461.000 1767.255 1461.640 ;
        RECT 1.445 1459.640 1763.200 1461.000 ;
        RECT 4.400 1459.600 1763.200 1459.640 ;
        RECT 4.400 1458.240 1767.255 1459.600 ;
        RECT 1.445 1456.240 1767.255 1458.240 ;
        RECT 4.400 1455.560 1767.255 1456.240 ;
        RECT 4.400 1454.840 1763.200 1455.560 ;
        RECT 1.445 1454.160 1763.200 1454.840 ;
        RECT 1.445 1452.840 1767.255 1454.160 ;
        RECT 4.400 1451.440 1767.255 1452.840 ;
        RECT 1.445 1450.120 1767.255 1451.440 ;
        RECT 1.445 1449.440 1763.200 1450.120 ;
        RECT 4.400 1448.720 1763.200 1449.440 ;
        RECT 4.400 1448.040 1767.255 1448.720 ;
        RECT 1.445 1446.040 1767.255 1448.040 ;
        RECT 4.400 1444.680 1767.255 1446.040 ;
        RECT 4.400 1444.640 1763.200 1444.680 ;
        RECT 1.445 1443.280 1763.200 1444.640 ;
        RECT 1.445 1441.960 1767.255 1443.280 ;
        RECT 4.400 1440.560 1767.255 1441.960 ;
        RECT 1.445 1439.240 1767.255 1440.560 ;
        RECT 1.445 1438.560 1763.200 1439.240 ;
        RECT 4.400 1437.840 1763.200 1438.560 ;
        RECT 4.400 1437.160 1767.255 1437.840 ;
        RECT 1.445 1435.160 1767.255 1437.160 ;
        RECT 4.400 1433.800 1767.255 1435.160 ;
        RECT 4.400 1433.760 1763.200 1433.800 ;
        RECT 1.445 1432.400 1763.200 1433.760 ;
        RECT 1.445 1431.760 1767.255 1432.400 ;
        RECT 4.400 1430.360 1767.255 1431.760 ;
        RECT 1.445 1428.360 1767.255 1430.360 ;
        RECT 4.400 1426.960 1763.200 1428.360 ;
        RECT 1.445 1424.960 1767.255 1426.960 ;
        RECT 4.400 1423.560 1767.255 1424.960 ;
        RECT 1.445 1422.920 1767.255 1423.560 ;
        RECT 1.445 1421.520 1763.200 1422.920 ;
        RECT 1.445 1420.880 1767.255 1421.520 ;
        RECT 4.400 1419.480 1767.255 1420.880 ;
        RECT 1.445 1417.480 1767.255 1419.480 ;
        RECT 4.400 1416.080 1763.200 1417.480 ;
        RECT 1.445 1414.080 1767.255 1416.080 ;
        RECT 4.400 1412.680 1767.255 1414.080 ;
        RECT 1.445 1412.040 1767.255 1412.680 ;
        RECT 1.445 1410.680 1763.200 1412.040 ;
        RECT 4.400 1410.640 1763.200 1410.680 ;
        RECT 4.400 1409.280 1767.255 1410.640 ;
        RECT 1.445 1407.280 1767.255 1409.280 ;
        RECT 4.400 1406.600 1767.255 1407.280 ;
        RECT 4.400 1405.880 1763.200 1406.600 ;
        RECT 1.445 1405.200 1763.200 1405.880 ;
        RECT 1.445 1403.200 1767.255 1405.200 ;
        RECT 4.400 1401.800 1767.255 1403.200 ;
        RECT 1.445 1401.160 1767.255 1401.800 ;
        RECT 1.445 1399.800 1763.200 1401.160 ;
        RECT 4.400 1399.760 1763.200 1399.800 ;
        RECT 4.400 1398.400 1767.255 1399.760 ;
        RECT 1.445 1396.400 1767.255 1398.400 ;
        RECT 4.400 1395.720 1767.255 1396.400 ;
        RECT 4.400 1395.000 1763.200 1395.720 ;
        RECT 1.445 1394.320 1763.200 1395.000 ;
        RECT 1.445 1393.000 1767.255 1394.320 ;
        RECT 4.400 1391.600 1767.255 1393.000 ;
        RECT 1.445 1390.280 1767.255 1391.600 ;
        RECT 1.445 1389.600 1763.200 1390.280 ;
        RECT 4.400 1388.880 1763.200 1389.600 ;
        RECT 4.400 1388.200 1767.255 1388.880 ;
        RECT 1.445 1386.200 1767.255 1388.200 ;
        RECT 4.400 1385.520 1767.255 1386.200 ;
        RECT 4.400 1384.800 1763.200 1385.520 ;
        RECT 1.445 1384.120 1763.200 1384.800 ;
        RECT 1.445 1382.120 1767.255 1384.120 ;
        RECT 4.400 1380.720 1767.255 1382.120 ;
        RECT 1.445 1380.080 1767.255 1380.720 ;
        RECT 1.445 1378.720 1763.200 1380.080 ;
        RECT 4.400 1378.680 1763.200 1378.720 ;
        RECT 4.400 1377.320 1767.255 1378.680 ;
        RECT 1.445 1375.320 1767.255 1377.320 ;
        RECT 4.400 1374.640 1767.255 1375.320 ;
        RECT 4.400 1373.920 1763.200 1374.640 ;
        RECT 1.445 1373.240 1763.200 1373.920 ;
        RECT 1.445 1371.920 1767.255 1373.240 ;
        RECT 4.400 1370.520 1767.255 1371.920 ;
        RECT 1.445 1369.200 1767.255 1370.520 ;
        RECT 1.445 1368.520 1763.200 1369.200 ;
        RECT 4.400 1367.800 1763.200 1368.520 ;
        RECT 4.400 1367.120 1767.255 1367.800 ;
        RECT 1.445 1364.440 1767.255 1367.120 ;
        RECT 4.400 1363.760 1767.255 1364.440 ;
        RECT 4.400 1363.040 1763.200 1363.760 ;
        RECT 1.445 1362.360 1763.200 1363.040 ;
        RECT 1.445 1361.040 1767.255 1362.360 ;
        RECT 4.400 1359.640 1767.255 1361.040 ;
        RECT 1.445 1358.320 1767.255 1359.640 ;
        RECT 1.445 1357.640 1763.200 1358.320 ;
        RECT 4.400 1356.920 1763.200 1357.640 ;
        RECT 4.400 1356.240 1767.255 1356.920 ;
        RECT 1.445 1354.240 1767.255 1356.240 ;
        RECT 4.400 1352.880 1767.255 1354.240 ;
        RECT 4.400 1352.840 1763.200 1352.880 ;
        RECT 1.445 1351.480 1763.200 1352.840 ;
        RECT 1.445 1350.840 1767.255 1351.480 ;
        RECT 4.400 1349.440 1767.255 1350.840 ;
        RECT 1.445 1347.440 1767.255 1349.440 ;
        RECT 4.400 1346.040 1763.200 1347.440 ;
        RECT 1.445 1343.360 1767.255 1346.040 ;
        RECT 4.400 1342.000 1767.255 1343.360 ;
        RECT 4.400 1341.960 1763.200 1342.000 ;
        RECT 1.445 1340.600 1763.200 1341.960 ;
        RECT 1.445 1339.960 1767.255 1340.600 ;
        RECT 4.400 1338.560 1767.255 1339.960 ;
        RECT 1.445 1336.560 1767.255 1338.560 ;
        RECT 4.400 1335.160 1763.200 1336.560 ;
        RECT 1.445 1333.160 1767.255 1335.160 ;
        RECT 4.400 1331.760 1767.255 1333.160 ;
        RECT 1.445 1331.120 1767.255 1331.760 ;
        RECT 1.445 1329.760 1763.200 1331.120 ;
        RECT 4.400 1329.720 1763.200 1329.760 ;
        RECT 4.400 1328.360 1767.255 1329.720 ;
        RECT 1.445 1326.360 1767.255 1328.360 ;
        RECT 4.400 1325.680 1767.255 1326.360 ;
        RECT 4.400 1324.960 1763.200 1325.680 ;
        RECT 1.445 1324.280 1763.200 1324.960 ;
        RECT 1.445 1322.280 1767.255 1324.280 ;
        RECT 4.400 1320.880 1767.255 1322.280 ;
        RECT 1.445 1320.240 1767.255 1320.880 ;
        RECT 1.445 1318.880 1763.200 1320.240 ;
        RECT 4.400 1318.840 1763.200 1318.880 ;
        RECT 4.400 1317.480 1767.255 1318.840 ;
        RECT 1.445 1315.480 1767.255 1317.480 ;
        RECT 4.400 1314.800 1767.255 1315.480 ;
        RECT 4.400 1314.080 1763.200 1314.800 ;
        RECT 1.445 1313.400 1763.200 1314.080 ;
        RECT 1.445 1312.080 1767.255 1313.400 ;
        RECT 4.400 1310.680 1767.255 1312.080 ;
        RECT 1.445 1309.360 1767.255 1310.680 ;
        RECT 1.445 1308.680 1763.200 1309.360 ;
        RECT 4.400 1307.960 1763.200 1308.680 ;
        RECT 4.400 1307.280 1767.255 1307.960 ;
        RECT 1.445 1304.600 1767.255 1307.280 ;
        RECT 4.400 1303.920 1767.255 1304.600 ;
        RECT 4.400 1303.200 1763.200 1303.920 ;
        RECT 1.445 1302.520 1763.200 1303.200 ;
        RECT 1.445 1301.200 1767.255 1302.520 ;
        RECT 4.400 1299.800 1767.255 1301.200 ;
        RECT 1.445 1298.480 1767.255 1299.800 ;
        RECT 1.445 1297.800 1763.200 1298.480 ;
        RECT 4.400 1297.080 1763.200 1297.800 ;
        RECT 4.400 1296.400 1767.255 1297.080 ;
        RECT 1.445 1294.400 1767.255 1296.400 ;
        RECT 4.400 1293.040 1767.255 1294.400 ;
        RECT 4.400 1293.000 1763.200 1293.040 ;
        RECT 1.445 1291.640 1763.200 1293.000 ;
        RECT 1.445 1291.000 1767.255 1291.640 ;
        RECT 4.400 1289.600 1767.255 1291.000 ;
        RECT 1.445 1287.600 1767.255 1289.600 ;
        RECT 4.400 1286.200 1763.200 1287.600 ;
        RECT 1.445 1283.520 1767.255 1286.200 ;
        RECT 4.400 1282.160 1767.255 1283.520 ;
        RECT 4.400 1282.120 1763.200 1282.160 ;
        RECT 1.445 1280.760 1763.200 1282.120 ;
        RECT 1.445 1280.120 1767.255 1280.760 ;
        RECT 4.400 1278.720 1767.255 1280.120 ;
        RECT 1.445 1276.720 1767.255 1278.720 ;
        RECT 4.400 1275.320 1763.200 1276.720 ;
        RECT 1.445 1273.320 1767.255 1275.320 ;
        RECT 4.400 1271.920 1767.255 1273.320 ;
        RECT 1.445 1271.280 1767.255 1271.920 ;
        RECT 1.445 1269.920 1763.200 1271.280 ;
        RECT 4.400 1269.880 1763.200 1269.920 ;
        RECT 4.400 1268.520 1767.255 1269.880 ;
        RECT 1.445 1265.840 1767.255 1268.520 ;
        RECT 4.400 1264.440 1763.200 1265.840 ;
        RECT 1.445 1262.440 1767.255 1264.440 ;
        RECT 4.400 1261.040 1767.255 1262.440 ;
        RECT 1.445 1260.400 1767.255 1261.040 ;
        RECT 1.445 1259.040 1763.200 1260.400 ;
        RECT 4.400 1259.000 1763.200 1259.040 ;
        RECT 4.400 1257.640 1767.255 1259.000 ;
        RECT 1.445 1255.640 1767.255 1257.640 ;
        RECT 4.400 1254.960 1767.255 1255.640 ;
        RECT 4.400 1254.240 1763.200 1254.960 ;
        RECT 1.445 1253.560 1763.200 1254.240 ;
        RECT 1.445 1252.240 1767.255 1253.560 ;
        RECT 4.400 1250.840 1767.255 1252.240 ;
        RECT 1.445 1249.520 1767.255 1250.840 ;
        RECT 1.445 1248.840 1763.200 1249.520 ;
        RECT 4.400 1248.120 1763.200 1248.840 ;
        RECT 4.400 1247.440 1767.255 1248.120 ;
        RECT 1.445 1244.760 1767.255 1247.440 ;
        RECT 4.400 1244.080 1767.255 1244.760 ;
        RECT 4.400 1243.360 1763.200 1244.080 ;
        RECT 1.445 1242.680 1763.200 1243.360 ;
        RECT 1.445 1241.360 1767.255 1242.680 ;
        RECT 4.400 1239.960 1767.255 1241.360 ;
        RECT 1.445 1238.640 1767.255 1239.960 ;
        RECT 1.445 1237.960 1763.200 1238.640 ;
        RECT 4.400 1237.240 1763.200 1237.960 ;
        RECT 4.400 1236.560 1767.255 1237.240 ;
        RECT 1.445 1234.560 1767.255 1236.560 ;
        RECT 4.400 1233.200 1767.255 1234.560 ;
        RECT 4.400 1233.160 1763.200 1233.200 ;
        RECT 1.445 1231.800 1763.200 1233.160 ;
        RECT 1.445 1231.160 1767.255 1231.800 ;
        RECT 4.400 1229.760 1767.255 1231.160 ;
        RECT 1.445 1227.760 1767.255 1229.760 ;
        RECT 4.400 1226.360 1763.200 1227.760 ;
        RECT 1.445 1223.680 1767.255 1226.360 ;
        RECT 4.400 1222.320 1767.255 1223.680 ;
        RECT 4.400 1222.280 1763.200 1222.320 ;
        RECT 1.445 1220.920 1763.200 1222.280 ;
        RECT 1.445 1220.280 1767.255 1220.920 ;
        RECT 4.400 1218.880 1767.255 1220.280 ;
        RECT 1.445 1216.880 1767.255 1218.880 ;
        RECT 4.400 1215.480 1763.200 1216.880 ;
        RECT 1.445 1213.480 1767.255 1215.480 ;
        RECT 4.400 1212.080 1767.255 1213.480 ;
        RECT 1.445 1211.440 1767.255 1212.080 ;
        RECT 1.445 1210.080 1763.200 1211.440 ;
        RECT 4.400 1210.040 1763.200 1210.080 ;
        RECT 4.400 1208.680 1767.255 1210.040 ;
        RECT 1.445 1206.000 1767.255 1208.680 ;
        RECT 4.400 1204.600 1763.200 1206.000 ;
        RECT 1.445 1202.600 1767.255 1204.600 ;
        RECT 4.400 1201.200 1767.255 1202.600 ;
        RECT 1.445 1200.560 1767.255 1201.200 ;
        RECT 1.445 1199.200 1763.200 1200.560 ;
        RECT 4.400 1199.160 1763.200 1199.200 ;
        RECT 4.400 1197.800 1767.255 1199.160 ;
        RECT 1.445 1195.800 1767.255 1197.800 ;
        RECT 4.400 1195.120 1767.255 1195.800 ;
        RECT 4.400 1194.400 1763.200 1195.120 ;
        RECT 1.445 1193.720 1763.200 1194.400 ;
        RECT 1.445 1192.400 1767.255 1193.720 ;
        RECT 4.400 1191.000 1767.255 1192.400 ;
        RECT 1.445 1189.680 1767.255 1191.000 ;
        RECT 1.445 1189.000 1763.200 1189.680 ;
        RECT 4.400 1188.280 1763.200 1189.000 ;
        RECT 4.400 1187.600 1767.255 1188.280 ;
        RECT 1.445 1184.920 1767.255 1187.600 ;
        RECT 4.400 1183.520 1763.200 1184.920 ;
        RECT 1.445 1181.520 1767.255 1183.520 ;
        RECT 4.400 1180.120 1767.255 1181.520 ;
        RECT 1.445 1179.480 1767.255 1180.120 ;
        RECT 1.445 1178.120 1763.200 1179.480 ;
        RECT 4.400 1178.080 1763.200 1178.120 ;
        RECT 4.400 1176.720 1767.255 1178.080 ;
        RECT 1.445 1174.720 1767.255 1176.720 ;
        RECT 4.400 1174.040 1767.255 1174.720 ;
        RECT 4.400 1173.320 1763.200 1174.040 ;
        RECT 1.445 1172.640 1763.200 1173.320 ;
        RECT 1.445 1171.320 1767.255 1172.640 ;
        RECT 4.400 1169.920 1767.255 1171.320 ;
        RECT 1.445 1168.600 1767.255 1169.920 ;
        RECT 1.445 1167.240 1763.200 1168.600 ;
        RECT 4.400 1167.200 1763.200 1167.240 ;
        RECT 4.400 1165.840 1767.255 1167.200 ;
        RECT 1.445 1163.840 1767.255 1165.840 ;
        RECT 4.400 1163.160 1767.255 1163.840 ;
        RECT 4.400 1162.440 1763.200 1163.160 ;
        RECT 1.445 1161.760 1763.200 1162.440 ;
        RECT 1.445 1160.440 1767.255 1161.760 ;
        RECT 4.400 1159.040 1767.255 1160.440 ;
        RECT 1.445 1157.720 1767.255 1159.040 ;
        RECT 1.445 1157.040 1763.200 1157.720 ;
        RECT 4.400 1156.320 1763.200 1157.040 ;
        RECT 4.400 1155.640 1767.255 1156.320 ;
        RECT 1.445 1153.640 1767.255 1155.640 ;
        RECT 4.400 1152.280 1767.255 1153.640 ;
        RECT 4.400 1152.240 1763.200 1152.280 ;
        RECT 1.445 1150.880 1763.200 1152.240 ;
        RECT 1.445 1150.240 1767.255 1150.880 ;
        RECT 4.400 1148.840 1767.255 1150.240 ;
        RECT 1.445 1146.840 1767.255 1148.840 ;
        RECT 1.445 1146.160 1763.200 1146.840 ;
        RECT 4.400 1145.440 1763.200 1146.160 ;
        RECT 4.400 1144.760 1767.255 1145.440 ;
        RECT 1.445 1142.760 1767.255 1144.760 ;
        RECT 4.400 1141.400 1767.255 1142.760 ;
        RECT 4.400 1141.360 1763.200 1141.400 ;
        RECT 1.445 1140.000 1763.200 1141.360 ;
        RECT 1.445 1139.360 1767.255 1140.000 ;
        RECT 4.400 1137.960 1767.255 1139.360 ;
        RECT 1.445 1135.960 1767.255 1137.960 ;
        RECT 4.400 1134.560 1763.200 1135.960 ;
        RECT 1.445 1132.560 1767.255 1134.560 ;
        RECT 4.400 1131.160 1767.255 1132.560 ;
        RECT 1.445 1130.520 1767.255 1131.160 ;
        RECT 1.445 1129.160 1763.200 1130.520 ;
        RECT 4.400 1129.120 1763.200 1129.160 ;
        RECT 4.400 1127.760 1767.255 1129.120 ;
        RECT 1.445 1125.080 1767.255 1127.760 ;
        RECT 4.400 1123.680 1763.200 1125.080 ;
        RECT 1.445 1121.680 1767.255 1123.680 ;
        RECT 4.400 1120.280 1767.255 1121.680 ;
        RECT 1.445 1119.640 1767.255 1120.280 ;
        RECT 1.445 1118.280 1763.200 1119.640 ;
        RECT 4.400 1118.240 1763.200 1118.280 ;
        RECT 4.400 1116.880 1767.255 1118.240 ;
        RECT 1.445 1114.880 1767.255 1116.880 ;
        RECT 4.400 1114.200 1767.255 1114.880 ;
        RECT 4.400 1113.480 1763.200 1114.200 ;
        RECT 1.445 1112.800 1763.200 1113.480 ;
        RECT 1.445 1111.480 1767.255 1112.800 ;
        RECT 4.400 1110.080 1767.255 1111.480 ;
        RECT 1.445 1108.760 1767.255 1110.080 ;
        RECT 1.445 1107.400 1763.200 1108.760 ;
        RECT 4.400 1107.360 1763.200 1107.400 ;
        RECT 4.400 1106.000 1767.255 1107.360 ;
        RECT 1.445 1104.000 1767.255 1106.000 ;
        RECT 4.400 1103.320 1767.255 1104.000 ;
        RECT 4.400 1102.600 1763.200 1103.320 ;
        RECT 1.445 1101.920 1763.200 1102.600 ;
        RECT 1.445 1100.600 1767.255 1101.920 ;
        RECT 4.400 1099.200 1767.255 1100.600 ;
        RECT 1.445 1097.880 1767.255 1099.200 ;
        RECT 1.445 1097.200 1763.200 1097.880 ;
        RECT 4.400 1096.480 1763.200 1097.200 ;
        RECT 4.400 1095.800 1767.255 1096.480 ;
        RECT 1.445 1093.800 1767.255 1095.800 ;
        RECT 4.400 1092.440 1767.255 1093.800 ;
        RECT 4.400 1092.400 1763.200 1092.440 ;
        RECT 1.445 1091.040 1763.200 1092.400 ;
        RECT 1.445 1090.400 1767.255 1091.040 ;
        RECT 4.400 1089.000 1767.255 1090.400 ;
        RECT 1.445 1087.000 1767.255 1089.000 ;
        RECT 1.445 1086.320 1763.200 1087.000 ;
        RECT 4.400 1085.600 1763.200 1086.320 ;
        RECT 4.400 1084.920 1767.255 1085.600 ;
        RECT 1.445 1082.920 1767.255 1084.920 ;
        RECT 4.400 1081.560 1767.255 1082.920 ;
        RECT 4.400 1081.520 1763.200 1081.560 ;
        RECT 1.445 1080.160 1763.200 1081.520 ;
        RECT 1.445 1079.520 1767.255 1080.160 ;
        RECT 4.400 1078.120 1767.255 1079.520 ;
        RECT 1.445 1076.120 1767.255 1078.120 ;
        RECT 4.400 1074.720 1763.200 1076.120 ;
        RECT 1.445 1072.720 1767.255 1074.720 ;
        RECT 4.400 1071.320 1767.255 1072.720 ;
        RECT 1.445 1070.680 1767.255 1071.320 ;
        RECT 1.445 1069.320 1763.200 1070.680 ;
        RECT 4.400 1069.280 1763.200 1069.320 ;
        RECT 4.400 1067.920 1767.255 1069.280 ;
        RECT 1.445 1065.240 1767.255 1067.920 ;
        RECT 4.400 1063.840 1763.200 1065.240 ;
        RECT 1.445 1061.840 1767.255 1063.840 ;
        RECT 4.400 1060.440 1767.255 1061.840 ;
        RECT 1.445 1059.800 1767.255 1060.440 ;
        RECT 1.445 1058.440 1763.200 1059.800 ;
        RECT 4.400 1058.400 1763.200 1058.440 ;
        RECT 4.400 1057.040 1767.255 1058.400 ;
        RECT 1.445 1055.040 1767.255 1057.040 ;
        RECT 4.400 1054.360 1767.255 1055.040 ;
        RECT 4.400 1053.640 1763.200 1054.360 ;
        RECT 1.445 1052.960 1763.200 1053.640 ;
        RECT 1.445 1051.640 1767.255 1052.960 ;
        RECT 4.400 1050.240 1767.255 1051.640 ;
        RECT 1.445 1048.920 1767.255 1050.240 ;
        RECT 1.445 1047.560 1763.200 1048.920 ;
        RECT 4.400 1047.520 1763.200 1047.560 ;
        RECT 4.400 1046.160 1767.255 1047.520 ;
        RECT 1.445 1044.160 1767.255 1046.160 ;
        RECT 4.400 1043.480 1767.255 1044.160 ;
        RECT 4.400 1042.760 1763.200 1043.480 ;
        RECT 1.445 1042.080 1763.200 1042.760 ;
        RECT 1.445 1040.760 1767.255 1042.080 ;
        RECT 4.400 1039.360 1767.255 1040.760 ;
        RECT 1.445 1038.040 1767.255 1039.360 ;
        RECT 1.445 1037.360 1763.200 1038.040 ;
        RECT 4.400 1036.640 1763.200 1037.360 ;
        RECT 4.400 1035.960 1767.255 1036.640 ;
        RECT 1.445 1033.960 1767.255 1035.960 ;
        RECT 4.400 1032.600 1767.255 1033.960 ;
        RECT 4.400 1032.560 1763.200 1032.600 ;
        RECT 1.445 1031.200 1763.200 1032.560 ;
        RECT 1.445 1030.560 1767.255 1031.200 ;
        RECT 4.400 1029.160 1767.255 1030.560 ;
        RECT 1.445 1027.160 1767.255 1029.160 ;
        RECT 1.445 1026.480 1763.200 1027.160 ;
        RECT 4.400 1025.760 1763.200 1026.480 ;
        RECT 4.400 1025.080 1767.255 1025.760 ;
        RECT 1.445 1023.080 1767.255 1025.080 ;
        RECT 4.400 1021.720 1767.255 1023.080 ;
        RECT 4.400 1021.680 1763.200 1021.720 ;
        RECT 1.445 1020.320 1763.200 1021.680 ;
        RECT 1.445 1019.680 1767.255 1020.320 ;
        RECT 4.400 1018.280 1767.255 1019.680 ;
        RECT 1.445 1016.280 1767.255 1018.280 ;
        RECT 4.400 1014.880 1763.200 1016.280 ;
        RECT 1.445 1012.880 1767.255 1014.880 ;
        RECT 4.400 1011.480 1767.255 1012.880 ;
        RECT 1.445 1010.840 1767.255 1011.480 ;
        RECT 1.445 1009.440 1763.200 1010.840 ;
        RECT 1.445 1008.800 1767.255 1009.440 ;
        RECT 4.400 1007.400 1767.255 1008.800 ;
        RECT 1.445 1005.400 1767.255 1007.400 ;
        RECT 4.400 1004.000 1763.200 1005.400 ;
        RECT 1.445 1002.000 1767.255 1004.000 ;
        RECT 4.400 1000.600 1767.255 1002.000 ;
        RECT 1.445 999.960 1767.255 1000.600 ;
        RECT 1.445 998.600 1763.200 999.960 ;
        RECT 4.400 998.560 1763.200 998.600 ;
        RECT 4.400 997.200 1767.255 998.560 ;
        RECT 1.445 995.200 1767.255 997.200 ;
        RECT 4.400 994.520 1767.255 995.200 ;
        RECT 4.400 993.800 1763.200 994.520 ;
        RECT 1.445 993.120 1763.200 993.800 ;
        RECT 1.445 991.800 1767.255 993.120 ;
        RECT 4.400 990.400 1767.255 991.800 ;
        RECT 1.445 989.760 1767.255 990.400 ;
        RECT 1.445 988.360 1763.200 989.760 ;
        RECT 1.445 987.720 1767.255 988.360 ;
        RECT 4.400 986.320 1767.255 987.720 ;
        RECT 1.445 984.320 1767.255 986.320 ;
        RECT 4.400 982.920 1763.200 984.320 ;
        RECT 1.445 980.920 1767.255 982.920 ;
        RECT 4.400 979.520 1767.255 980.920 ;
        RECT 1.445 978.880 1767.255 979.520 ;
        RECT 1.445 977.520 1763.200 978.880 ;
        RECT 4.400 977.480 1763.200 977.520 ;
        RECT 4.400 976.120 1767.255 977.480 ;
        RECT 1.445 974.120 1767.255 976.120 ;
        RECT 4.400 973.440 1767.255 974.120 ;
        RECT 4.400 972.720 1763.200 973.440 ;
        RECT 1.445 972.040 1763.200 972.720 ;
        RECT 1.445 970.720 1767.255 972.040 ;
        RECT 4.400 969.320 1767.255 970.720 ;
        RECT 1.445 968.000 1767.255 969.320 ;
        RECT 1.445 966.640 1763.200 968.000 ;
        RECT 4.400 966.600 1763.200 966.640 ;
        RECT 4.400 965.240 1767.255 966.600 ;
        RECT 1.445 963.240 1767.255 965.240 ;
        RECT 4.400 962.560 1767.255 963.240 ;
        RECT 4.400 961.840 1763.200 962.560 ;
        RECT 1.445 961.160 1763.200 961.840 ;
        RECT 1.445 959.840 1767.255 961.160 ;
        RECT 4.400 958.440 1767.255 959.840 ;
        RECT 1.445 957.120 1767.255 958.440 ;
        RECT 1.445 956.440 1763.200 957.120 ;
        RECT 4.400 955.720 1763.200 956.440 ;
        RECT 4.400 955.040 1767.255 955.720 ;
        RECT 1.445 953.040 1767.255 955.040 ;
        RECT 4.400 951.680 1767.255 953.040 ;
        RECT 4.400 951.640 1763.200 951.680 ;
        RECT 1.445 950.280 1763.200 951.640 ;
        RECT 1.445 948.960 1767.255 950.280 ;
        RECT 4.400 947.560 1767.255 948.960 ;
        RECT 1.445 946.240 1767.255 947.560 ;
        RECT 1.445 945.560 1763.200 946.240 ;
        RECT 4.400 944.840 1763.200 945.560 ;
        RECT 4.400 944.160 1767.255 944.840 ;
        RECT 1.445 942.160 1767.255 944.160 ;
        RECT 4.400 940.800 1767.255 942.160 ;
        RECT 4.400 940.760 1763.200 940.800 ;
        RECT 1.445 939.400 1763.200 940.760 ;
        RECT 1.445 938.760 1767.255 939.400 ;
        RECT 4.400 937.360 1767.255 938.760 ;
        RECT 1.445 935.360 1767.255 937.360 ;
        RECT 4.400 933.960 1763.200 935.360 ;
        RECT 1.445 931.960 1767.255 933.960 ;
        RECT 4.400 930.560 1767.255 931.960 ;
        RECT 1.445 929.920 1767.255 930.560 ;
        RECT 1.445 928.520 1763.200 929.920 ;
        RECT 1.445 927.880 1767.255 928.520 ;
        RECT 4.400 926.480 1767.255 927.880 ;
        RECT 1.445 924.480 1767.255 926.480 ;
        RECT 4.400 923.080 1763.200 924.480 ;
        RECT 1.445 921.080 1767.255 923.080 ;
        RECT 4.400 919.680 1767.255 921.080 ;
        RECT 1.445 919.040 1767.255 919.680 ;
        RECT 1.445 917.680 1763.200 919.040 ;
        RECT 4.400 917.640 1763.200 917.680 ;
        RECT 4.400 916.280 1767.255 917.640 ;
        RECT 1.445 914.280 1767.255 916.280 ;
        RECT 4.400 913.600 1767.255 914.280 ;
        RECT 4.400 912.880 1763.200 913.600 ;
        RECT 1.445 912.200 1763.200 912.880 ;
        RECT 1.445 910.200 1767.255 912.200 ;
        RECT 4.400 908.800 1767.255 910.200 ;
        RECT 1.445 908.160 1767.255 908.800 ;
        RECT 1.445 906.800 1763.200 908.160 ;
        RECT 4.400 906.760 1763.200 906.800 ;
        RECT 4.400 905.400 1767.255 906.760 ;
        RECT 1.445 903.400 1767.255 905.400 ;
        RECT 4.400 902.720 1767.255 903.400 ;
        RECT 4.400 902.000 1763.200 902.720 ;
        RECT 1.445 901.320 1763.200 902.000 ;
        RECT 1.445 900.000 1767.255 901.320 ;
        RECT 4.400 898.600 1767.255 900.000 ;
        RECT 1.445 897.280 1767.255 898.600 ;
        RECT 1.445 896.600 1763.200 897.280 ;
        RECT 4.400 895.880 1763.200 896.600 ;
        RECT 4.400 895.200 1767.255 895.880 ;
        RECT 1.445 893.200 1767.255 895.200 ;
        RECT 4.400 891.840 1767.255 893.200 ;
        RECT 4.400 891.800 1763.200 891.840 ;
        RECT 1.445 890.440 1763.200 891.800 ;
        RECT 1.445 889.120 1767.255 890.440 ;
        RECT 4.400 887.720 1767.255 889.120 ;
        RECT 1.445 886.400 1767.255 887.720 ;
        RECT 1.445 885.720 1763.200 886.400 ;
        RECT 4.400 885.000 1763.200 885.720 ;
        RECT 4.400 884.320 1767.255 885.000 ;
        RECT 1.445 882.320 1767.255 884.320 ;
        RECT 4.400 880.960 1767.255 882.320 ;
        RECT 4.400 880.920 1763.200 880.960 ;
        RECT 1.445 879.560 1763.200 880.920 ;
        RECT 1.445 878.920 1767.255 879.560 ;
        RECT 4.400 877.520 1767.255 878.920 ;
        RECT 1.445 875.520 1767.255 877.520 ;
        RECT 4.400 874.120 1763.200 875.520 ;
        RECT 1.445 872.120 1767.255 874.120 ;
        RECT 4.400 870.720 1767.255 872.120 ;
        RECT 1.445 870.080 1767.255 870.720 ;
        RECT 1.445 868.680 1763.200 870.080 ;
        RECT 1.445 868.040 1767.255 868.680 ;
        RECT 4.400 866.640 1767.255 868.040 ;
        RECT 1.445 864.640 1767.255 866.640 ;
        RECT 4.400 863.240 1763.200 864.640 ;
        RECT 1.445 861.240 1767.255 863.240 ;
        RECT 4.400 859.840 1767.255 861.240 ;
        RECT 1.445 859.200 1767.255 859.840 ;
        RECT 1.445 857.840 1763.200 859.200 ;
        RECT 4.400 857.800 1763.200 857.840 ;
        RECT 4.400 856.440 1767.255 857.800 ;
        RECT 1.445 854.440 1767.255 856.440 ;
        RECT 4.400 853.760 1767.255 854.440 ;
        RECT 4.400 853.040 1763.200 853.760 ;
        RECT 1.445 852.360 1763.200 853.040 ;
        RECT 1.445 850.360 1767.255 852.360 ;
        RECT 4.400 848.960 1767.255 850.360 ;
        RECT 1.445 848.320 1767.255 848.960 ;
        RECT 1.445 846.960 1763.200 848.320 ;
        RECT 4.400 846.920 1763.200 846.960 ;
        RECT 4.400 845.560 1767.255 846.920 ;
        RECT 1.445 843.560 1767.255 845.560 ;
        RECT 4.400 842.880 1767.255 843.560 ;
        RECT 4.400 842.160 1763.200 842.880 ;
        RECT 1.445 841.480 1763.200 842.160 ;
        RECT 1.445 840.160 1767.255 841.480 ;
        RECT 4.400 838.760 1767.255 840.160 ;
        RECT 1.445 837.440 1767.255 838.760 ;
        RECT 1.445 836.760 1763.200 837.440 ;
        RECT 4.400 836.040 1763.200 836.760 ;
        RECT 4.400 835.360 1767.255 836.040 ;
        RECT 1.445 833.360 1767.255 835.360 ;
        RECT 4.400 832.000 1767.255 833.360 ;
        RECT 4.400 831.960 1763.200 832.000 ;
        RECT 1.445 830.600 1763.200 831.960 ;
        RECT 1.445 829.280 1767.255 830.600 ;
        RECT 4.400 827.880 1767.255 829.280 ;
        RECT 1.445 826.560 1767.255 827.880 ;
        RECT 1.445 825.880 1763.200 826.560 ;
        RECT 4.400 825.160 1763.200 825.880 ;
        RECT 4.400 824.480 1767.255 825.160 ;
        RECT 1.445 822.480 1767.255 824.480 ;
        RECT 4.400 821.120 1767.255 822.480 ;
        RECT 4.400 821.080 1763.200 821.120 ;
        RECT 1.445 819.720 1763.200 821.080 ;
        RECT 1.445 819.080 1767.255 819.720 ;
        RECT 4.400 817.680 1767.255 819.080 ;
        RECT 1.445 815.680 1767.255 817.680 ;
        RECT 4.400 814.280 1763.200 815.680 ;
        RECT 1.445 811.600 1767.255 814.280 ;
        RECT 4.400 810.240 1767.255 811.600 ;
        RECT 4.400 810.200 1763.200 810.240 ;
        RECT 1.445 808.840 1763.200 810.200 ;
        RECT 1.445 808.200 1767.255 808.840 ;
        RECT 4.400 806.800 1767.255 808.200 ;
        RECT 1.445 804.800 1767.255 806.800 ;
        RECT 4.400 803.400 1763.200 804.800 ;
        RECT 1.445 801.400 1767.255 803.400 ;
        RECT 4.400 800.000 1767.255 801.400 ;
        RECT 1.445 799.360 1767.255 800.000 ;
        RECT 1.445 798.000 1763.200 799.360 ;
        RECT 4.400 797.960 1763.200 798.000 ;
        RECT 4.400 796.600 1767.255 797.960 ;
        RECT 1.445 794.600 1767.255 796.600 ;
        RECT 4.400 793.920 1767.255 794.600 ;
        RECT 4.400 793.200 1763.200 793.920 ;
        RECT 1.445 792.520 1763.200 793.200 ;
        RECT 1.445 790.520 1767.255 792.520 ;
        RECT 4.400 789.160 1767.255 790.520 ;
        RECT 4.400 789.120 1763.200 789.160 ;
        RECT 1.445 787.760 1763.200 789.120 ;
        RECT 1.445 787.120 1767.255 787.760 ;
        RECT 4.400 785.720 1767.255 787.120 ;
        RECT 1.445 783.720 1767.255 785.720 ;
        RECT 4.400 782.320 1763.200 783.720 ;
        RECT 1.445 780.320 1767.255 782.320 ;
        RECT 4.400 778.920 1767.255 780.320 ;
        RECT 1.445 778.280 1767.255 778.920 ;
        RECT 1.445 776.920 1763.200 778.280 ;
        RECT 4.400 776.880 1763.200 776.920 ;
        RECT 4.400 775.520 1767.255 776.880 ;
        RECT 1.445 773.520 1767.255 775.520 ;
        RECT 4.400 772.840 1767.255 773.520 ;
        RECT 4.400 772.120 1763.200 772.840 ;
        RECT 1.445 771.440 1763.200 772.120 ;
        RECT 1.445 769.440 1767.255 771.440 ;
        RECT 4.400 768.040 1767.255 769.440 ;
        RECT 1.445 767.400 1767.255 768.040 ;
        RECT 1.445 766.040 1763.200 767.400 ;
        RECT 4.400 766.000 1763.200 766.040 ;
        RECT 4.400 764.640 1767.255 766.000 ;
        RECT 1.445 762.640 1767.255 764.640 ;
        RECT 4.400 761.960 1767.255 762.640 ;
        RECT 4.400 761.240 1763.200 761.960 ;
        RECT 1.445 760.560 1763.200 761.240 ;
        RECT 1.445 759.240 1767.255 760.560 ;
        RECT 4.400 757.840 1767.255 759.240 ;
        RECT 1.445 756.520 1767.255 757.840 ;
        RECT 1.445 755.840 1763.200 756.520 ;
        RECT 4.400 755.120 1763.200 755.840 ;
        RECT 4.400 754.440 1767.255 755.120 ;
        RECT 1.445 751.760 1767.255 754.440 ;
        RECT 4.400 751.080 1767.255 751.760 ;
        RECT 4.400 750.360 1763.200 751.080 ;
        RECT 1.445 749.680 1763.200 750.360 ;
        RECT 1.445 748.360 1767.255 749.680 ;
        RECT 4.400 746.960 1767.255 748.360 ;
        RECT 1.445 745.640 1767.255 746.960 ;
        RECT 1.445 744.960 1763.200 745.640 ;
        RECT 4.400 744.240 1763.200 744.960 ;
        RECT 4.400 743.560 1767.255 744.240 ;
        RECT 1.445 741.560 1767.255 743.560 ;
        RECT 4.400 740.200 1767.255 741.560 ;
        RECT 4.400 740.160 1763.200 740.200 ;
        RECT 1.445 738.800 1763.200 740.160 ;
        RECT 1.445 738.160 1767.255 738.800 ;
        RECT 4.400 736.760 1767.255 738.160 ;
        RECT 1.445 734.760 1767.255 736.760 ;
        RECT 4.400 733.360 1763.200 734.760 ;
        RECT 1.445 730.680 1767.255 733.360 ;
        RECT 4.400 729.320 1767.255 730.680 ;
        RECT 4.400 729.280 1763.200 729.320 ;
        RECT 1.445 727.920 1763.200 729.280 ;
        RECT 1.445 727.280 1767.255 727.920 ;
        RECT 4.400 725.880 1767.255 727.280 ;
        RECT 1.445 723.880 1767.255 725.880 ;
        RECT 4.400 722.480 1763.200 723.880 ;
        RECT 1.445 720.480 1767.255 722.480 ;
        RECT 4.400 719.080 1767.255 720.480 ;
        RECT 1.445 718.440 1767.255 719.080 ;
        RECT 1.445 717.080 1763.200 718.440 ;
        RECT 4.400 717.040 1763.200 717.080 ;
        RECT 4.400 715.680 1767.255 717.040 ;
        RECT 1.445 713.680 1767.255 715.680 ;
        RECT 4.400 713.000 1767.255 713.680 ;
        RECT 4.400 712.280 1763.200 713.000 ;
        RECT 1.445 711.600 1763.200 712.280 ;
        RECT 1.445 709.600 1767.255 711.600 ;
        RECT 4.400 708.200 1767.255 709.600 ;
        RECT 1.445 707.560 1767.255 708.200 ;
        RECT 1.445 706.200 1763.200 707.560 ;
        RECT 4.400 706.160 1763.200 706.200 ;
        RECT 4.400 704.800 1767.255 706.160 ;
        RECT 1.445 702.800 1767.255 704.800 ;
        RECT 4.400 702.120 1767.255 702.800 ;
        RECT 4.400 701.400 1763.200 702.120 ;
        RECT 1.445 700.720 1763.200 701.400 ;
        RECT 1.445 699.400 1767.255 700.720 ;
        RECT 4.400 698.000 1767.255 699.400 ;
        RECT 1.445 696.680 1767.255 698.000 ;
        RECT 1.445 696.000 1763.200 696.680 ;
        RECT 4.400 695.280 1763.200 696.000 ;
        RECT 4.400 694.600 1767.255 695.280 ;
        RECT 1.445 691.920 1767.255 694.600 ;
        RECT 4.400 691.240 1767.255 691.920 ;
        RECT 4.400 690.520 1763.200 691.240 ;
        RECT 1.445 689.840 1763.200 690.520 ;
        RECT 1.445 688.520 1767.255 689.840 ;
        RECT 4.400 687.120 1767.255 688.520 ;
        RECT 1.445 685.800 1767.255 687.120 ;
        RECT 1.445 685.120 1763.200 685.800 ;
        RECT 4.400 684.400 1763.200 685.120 ;
        RECT 4.400 683.720 1767.255 684.400 ;
        RECT 1.445 681.720 1767.255 683.720 ;
        RECT 4.400 680.360 1767.255 681.720 ;
        RECT 4.400 680.320 1763.200 680.360 ;
        RECT 1.445 678.960 1763.200 680.320 ;
        RECT 1.445 678.320 1767.255 678.960 ;
        RECT 4.400 676.920 1767.255 678.320 ;
        RECT 1.445 674.920 1767.255 676.920 ;
        RECT 4.400 673.520 1763.200 674.920 ;
        RECT 1.445 670.840 1767.255 673.520 ;
        RECT 4.400 669.480 1767.255 670.840 ;
        RECT 4.400 669.440 1763.200 669.480 ;
        RECT 1.445 668.080 1763.200 669.440 ;
        RECT 1.445 667.440 1767.255 668.080 ;
        RECT 4.400 666.040 1767.255 667.440 ;
        RECT 1.445 664.040 1767.255 666.040 ;
        RECT 4.400 662.640 1763.200 664.040 ;
        RECT 1.445 660.640 1767.255 662.640 ;
        RECT 4.400 659.240 1767.255 660.640 ;
        RECT 1.445 658.600 1767.255 659.240 ;
        RECT 1.445 657.240 1763.200 658.600 ;
        RECT 4.400 657.200 1763.200 657.240 ;
        RECT 4.400 655.840 1767.255 657.200 ;
        RECT 1.445 653.160 1767.255 655.840 ;
        RECT 4.400 651.760 1763.200 653.160 ;
        RECT 1.445 649.760 1767.255 651.760 ;
        RECT 4.400 648.360 1767.255 649.760 ;
        RECT 1.445 647.720 1767.255 648.360 ;
        RECT 1.445 646.360 1763.200 647.720 ;
        RECT 4.400 646.320 1763.200 646.360 ;
        RECT 4.400 644.960 1767.255 646.320 ;
        RECT 1.445 642.960 1767.255 644.960 ;
        RECT 4.400 642.280 1767.255 642.960 ;
        RECT 4.400 641.560 1763.200 642.280 ;
        RECT 1.445 640.880 1763.200 641.560 ;
        RECT 1.445 639.560 1767.255 640.880 ;
        RECT 4.400 638.160 1767.255 639.560 ;
        RECT 1.445 636.840 1767.255 638.160 ;
        RECT 1.445 636.160 1763.200 636.840 ;
        RECT 4.400 635.440 1763.200 636.160 ;
        RECT 4.400 634.760 1767.255 635.440 ;
        RECT 1.445 632.080 1767.255 634.760 ;
        RECT 4.400 631.400 1767.255 632.080 ;
        RECT 4.400 630.680 1763.200 631.400 ;
        RECT 1.445 630.000 1763.200 630.680 ;
        RECT 1.445 628.680 1767.255 630.000 ;
        RECT 4.400 627.280 1767.255 628.680 ;
        RECT 1.445 625.960 1767.255 627.280 ;
        RECT 1.445 625.280 1763.200 625.960 ;
        RECT 4.400 624.560 1763.200 625.280 ;
        RECT 4.400 623.880 1767.255 624.560 ;
        RECT 1.445 621.880 1767.255 623.880 ;
        RECT 4.400 620.520 1767.255 621.880 ;
        RECT 4.400 620.480 1763.200 620.520 ;
        RECT 1.445 619.120 1763.200 620.480 ;
        RECT 1.445 618.480 1767.255 619.120 ;
        RECT 4.400 617.080 1767.255 618.480 ;
        RECT 1.445 615.080 1767.255 617.080 ;
        RECT 4.400 613.680 1763.200 615.080 ;
        RECT 1.445 611.000 1767.255 613.680 ;
        RECT 4.400 609.640 1767.255 611.000 ;
        RECT 4.400 609.600 1763.200 609.640 ;
        RECT 1.445 608.240 1763.200 609.600 ;
        RECT 1.445 607.600 1767.255 608.240 ;
        RECT 4.400 606.200 1767.255 607.600 ;
        RECT 1.445 604.200 1767.255 606.200 ;
        RECT 4.400 602.800 1763.200 604.200 ;
        RECT 1.445 600.800 1767.255 602.800 ;
        RECT 4.400 599.400 1767.255 600.800 ;
        RECT 1.445 598.760 1767.255 599.400 ;
        RECT 1.445 597.400 1763.200 598.760 ;
        RECT 4.400 597.360 1763.200 597.400 ;
        RECT 4.400 596.000 1767.255 597.360 ;
        RECT 1.445 594.000 1767.255 596.000 ;
        RECT 1.445 593.320 1763.200 594.000 ;
        RECT 4.400 592.600 1763.200 593.320 ;
        RECT 4.400 591.920 1767.255 592.600 ;
        RECT 1.445 589.920 1767.255 591.920 ;
        RECT 4.400 588.560 1767.255 589.920 ;
        RECT 4.400 588.520 1763.200 588.560 ;
        RECT 1.445 587.160 1763.200 588.520 ;
        RECT 1.445 586.520 1767.255 587.160 ;
        RECT 4.400 585.120 1767.255 586.520 ;
        RECT 1.445 583.120 1767.255 585.120 ;
        RECT 4.400 581.720 1763.200 583.120 ;
        RECT 1.445 579.720 1767.255 581.720 ;
        RECT 4.400 578.320 1767.255 579.720 ;
        RECT 1.445 577.680 1767.255 578.320 ;
        RECT 1.445 576.320 1763.200 577.680 ;
        RECT 4.400 576.280 1763.200 576.320 ;
        RECT 4.400 574.920 1767.255 576.280 ;
        RECT 1.445 572.240 1767.255 574.920 ;
        RECT 4.400 570.840 1763.200 572.240 ;
        RECT 1.445 568.840 1767.255 570.840 ;
        RECT 4.400 567.440 1767.255 568.840 ;
        RECT 1.445 566.800 1767.255 567.440 ;
        RECT 1.445 565.440 1763.200 566.800 ;
        RECT 4.400 565.400 1763.200 565.440 ;
        RECT 4.400 564.040 1767.255 565.400 ;
        RECT 1.445 562.040 1767.255 564.040 ;
        RECT 4.400 561.360 1767.255 562.040 ;
        RECT 4.400 560.640 1763.200 561.360 ;
        RECT 1.445 559.960 1763.200 560.640 ;
        RECT 1.445 558.640 1767.255 559.960 ;
        RECT 4.400 557.240 1767.255 558.640 ;
        RECT 1.445 555.920 1767.255 557.240 ;
        RECT 1.445 554.560 1763.200 555.920 ;
        RECT 4.400 554.520 1763.200 554.560 ;
        RECT 4.400 553.160 1767.255 554.520 ;
        RECT 1.445 551.160 1767.255 553.160 ;
        RECT 4.400 550.480 1767.255 551.160 ;
        RECT 4.400 549.760 1763.200 550.480 ;
        RECT 1.445 549.080 1763.200 549.760 ;
        RECT 1.445 547.760 1767.255 549.080 ;
        RECT 4.400 546.360 1767.255 547.760 ;
        RECT 1.445 545.040 1767.255 546.360 ;
        RECT 1.445 544.360 1763.200 545.040 ;
        RECT 4.400 543.640 1763.200 544.360 ;
        RECT 4.400 542.960 1767.255 543.640 ;
        RECT 1.445 540.960 1767.255 542.960 ;
        RECT 4.400 539.600 1767.255 540.960 ;
        RECT 4.400 539.560 1763.200 539.600 ;
        RECT 1.445 538.200 1763.200 539.560 ;
        RECT 1.445 537.560 1767.255 538.200 ;
        RECT 4.400 536.160 1767.255 537.560 ;
        RECT 1.445 534.160 1767.255 536.160 ;
        RECT 1.445 533.480 1763.200 534.160 ;
        RECT 4.400 532.760 1763.200 533.480 ;
        RECT 4.400 532.080 1767.255 532.760 ;
        RECT 1.445 530.080 1767.255 532.080 ;
        RECT 4.400 528.720 1767.255 530.080 ;
        RECT 4.400 528.680 1763.200 528.720 ;
        RECT 1.445 527.320 1763.200 528.680 ;
        RECT 1.445 526.680 1767.255 527.320 ;
        RECT 4.400 525.280 1767.255 526.680 ;
        RECT 1.445 523.280 1767.255 525.280 ;
        RECT 4.400 521.880 1763.200 523.280 ;
        RECT 1.445 519.880 1767.255 521.880 ;
        RECT 4.400 518.480 1767.255 519.880 ;
        RECT 1.445 517.840 1767.255 518.480 ;
        RECT 1.445 516.480 1763.200 517.840 ;
        RECT 4.400 516.440 1763.200 516.480 ;
        RECT 4.400 515.080 1767.255 516.440 ;
        RECT 1.445 512.400 1767.255 515.080 ;
        RECT 4.400 511.000 1763.200 512.400 ;
        RECT 1.445 509.000 1767.255 511.000 ;
        RECT 4.400 507.600 1767.255 509.000 ;
        RECT 1.445 506.960 1767.255 507.600 ;
        RECT 1.445 505.600 1763.200 506.960 ;
        RECT 4.400 505.560 1763.200 505.600 ;
        RECT 4.400 504.200 1767.255 505.560 ;
        RECT 1.445 502.200 1767.255 504.200 ;
        RECT 4.400 501.520 1767.255 502.200 ;
        RECT 4.400 500.800 1763.200 501.520 ;
        RECT 1.445 500.120 1763.200 500.800 ;
        RECT 1.445 498.800 1767.255 500.120 ;
        RECT 4.400 497.400 1767.255 498.800 ;
        RECT 1.445 496.080 1767.255 497.400 ;
        RECT 1.445 494.720 1763.200 496.080 ;
        RECT 4.400 494.680 1763.200 494.720 ;
        RECT 4.400 493.320 1767.255 494.680 ;
        RECT 1.445 491.320 1767.255 493.320 ;
        RECT 4.400 490.640 1767.255 491.320 ;
        RECT 4.400 489.920 1763.200 490.640 ;
        RECT 1.445 489.240 1763.200 489.920 ;
        RECT 1.445 487.920 1767.255 489.240 ;
        RECT 4.400 486.520 1767.255 487.920 ;
        RECT 1.445 485.200 1767.255 486.520 ;
        RECT 1.445 484.520 1763.200 485.200 ;
        RECT 4.400 483.800 1763.200 484.520 ;
        RECT 4.400 483.120 1767.255 483.800 ;
        RECT 1.445 481.120 1767.255 483.120 ;
        RECT 4.400 479.760 1767.255 481.120 ;
        RECT 4.400 479.720 1763.200 479.760 ;
        RECT 1.445 478.360 1763.200 479.720 ;
        RECT 1.445 477.720 1767.255 478.360 ;
        RECT 4.400 476.320 1767.255 477.720 ;
        RECT 1.445 474.320 1767.255 476.320 ;
        RECT 1.445 473.640 1763.200 474.320 ;
        RECT 4.400 472.920 1763.200 473.640 ;
        RECT 4.400 472.240 1767.255 472.920 ;
        RECT 1.445 470.240 1767.255 472.240 ;
        RECT 4.400 468.880 1767.255 470.240 ;
        RECT 4.400 468.840 1763.200 468.880 ;
        RECT 1.445 467.480 1763.200 468.840 ;
        RECT 1.445 466.840 1767.255 467.480 ;
        RECT 4.400 465.440 1767.255 466.840 ;
        RECT 1.445 463.440 1767.255 465.440 ;
        RECT 4.400 462.040 1763.200 463.440 ;
        RECT 1.445 460.040 1767.255 462.040 ;
        RECT 4.400 458.640 1767.255 460.040 ;
        RECT 1.445 458.000 1767.255 458.640 ;
        RECT 1.445 456.600 1763.200 458.000 ;
        RECT 1.445 455.960 1767.255 456.600 ;
        RECT 4.400 454.560 1767.255 455.960 ;
        RECT 1.445 452.560 1767.255 454.560 ;
        RECT 4.400 451.160 1763.200 452.560 ;
        RECT 1.445 449.160 1767.255 451.160 ;
        RECT 4.400 447.760 1767.255 449.160 ;
        RECT 1.445 447.120 1767.255 447.760 ;
        RECT 1.445 445.760 1763.200 447.120 ;
        RECT 4.400 445.720 1763.200 445.760 ;
        RECT 4.400 444.360 1767.255 445.720 ;
        RECT 1.445 442.360 1767.255 444.360 ;
        RECT 4.400 441.680 1767.255 442.360 ;
        RECT 4.400 440.960 1763.200 441.680 ;
        RECT 1.445 440.280 1763.200 440.960 ;
        RECT 1.445 438.960 1767.255 440.280 ;
        RECT 4.400 437.560 1767.255 438.960 ;
        RECT 1.445 436.240 1767.255 437.560 ;
        RECT 1.445 434.880 1763.200 436.240 ;
        RECT 4.400 434.840 1763.200 434.880 ;
        RECT 4.400 433.480 1767.255 434.840 ;
        RECT 1.445 431.480 1767.255 433.480 ;
        RECT 4.400 430.800 1767.255 431.480 ;
        RECT 4.400 430.080 1763.200 430.800 ;
        RECT 1.445 429.400 1763.200 430.080 ;
        RECT 1.445 428.080 1767.255 429.400 ;
        RECT 4.400 426.680 1767.255 428.080 ;
        RECT 1.445 425.360 1767.255 426.680 ;
        RECT 1.445 424.680 1763.200 425.360 ;
        RECT 4.400 423.960 1763.200 424.680 ;
        RECT 4.400 423.280 1767.255 423.960 ;
        RECT 1.445 421.280 1767.255 423.280 ;
        RECT 4.400 419.920 1767.255 421.280 ;
        RECT 4.400 419.880 1763.200 419.920 ;
        RECT 1.445 418.520 1763.200 419.880 ;
        RECT 1.445 417.880 1767.255 418.520 ;
        RECT 4.400 416.480 1767.255 417.880 ;
        RECT 1.445 414.480 1767.255 416.480 ;
        RECT 1.445 413.800 1763.200 414.480 ;
        RECT 4.400 413.080 1763.200 413.800 ;
        RECT 4.400 412.400 1767.255 413.080 ;
        RECT 1.445 410.400 1767.255 412.400 ;
        RECT 4.400 409.040 1767.255 410.400 ;
        RECT 4.400 409.000 1763.200 409.040 ;
        RECT 1.445 407.640 1763.200 409.000 ;
        RECT 1.445 407.000 1767.255 407.640 ;
        RECT 4.400 405.600 1767.255 407.000 ;
        RECT 1.445 403.600 1767.255 405.600 ;
        RECT 4.400 402.200 1763.200 403.600 ;
        RECT 1.445 400.200 1767.255 402.200 ;
        RECT 4.400 398.800 1767.255 400.200 ;
        RECT 1.445 398.160 1767.255 398.800 ;
        RECT 1.445 396.760 1763.200 398.160 ;
        RECT 1.445 396.120 1767.255 396.760 ;
        RECT 4.400 394.720 1767.255 396.120 ;
        RECT 1.445 393.400 1767.255 394.720 ;
        RECT 1.445 392.720 1763.200 393.400 ;
        RECT 4.400 392.000 1763.200 392.720 ;
        RECT 4.400 391.320 1767.255 392.000 ;
        RECT 1.445 389.320 1767.255 391.320 ;
        RECT 4.400 387.960 1767.255 389.320 ;
        RECT 4.400 387.920 1763.200 387.960 ;
        RECT 1.445 386.560 1763.200 387.920 ;
        RECT 1.445 385.920 1767.255 386.560 ;
        RECT 4.400 384.520 1767.255 385.920 ;
        RECT 1.445 382.520 1767.255 384.520 ;
        RECT 4.400 381.120 1763.200 382.520 ;
        RECT 1.445 379.120 1767.255 381.120 ;
        RECT 4.400 377.720 1767.255 379.120 ;
        RECT 1.445 377.080 1767.255 377.720 ;
        RECT 1.445 375.680 1763.200 377.080 ;
        RECT 1.445 375.040 1767.255 375.680 ;
        RECT 4.400 373.640 1767.255 375.040 ;
        RECT 1.445 371.640 1767.255 373.640 ;
        RECT 4.400 370.240 1763.200 371.640 ;
        RECT 1.445 368.240 1767.255 370.240 ;
        RECT 4.400 366.840 1767.255 368.240 ;
        RECT 1.445 366.200 1767.255 366.840 ;
        RECT 1.445 364.840 1763.200 366.200 ;
        RECT 4.400 364.800 1763.200 364.840 ;
        RECT 4.400 363.440 1767.255 364.800 ;
        RECT 1.445 361.440 1767.255 363.440 ;
        RECT 4.400 360.760 1767.255 361.440 ;
        RECT 4.400 360.040 1763.200 360.760 ;
        RECT 1.445 359.360 1763.200 360.040 ;
        RECT 1.445 358.040 1767.255 359.360 ;
        RECT 4.400 356.640 1767.255 358.040 ;
        RECT 1.445 355.320 1767.255 356.640 ;
        RECT 1.445 353.960 1763.200 355.320 ;
        RECT 4.400 353.920 1763.200 353.960 ;
        RECT 4.400 352.560 1767.255 353.920 ;
        RECT 1.445 350.560 1767.255 352.560 ;
        RECT 4.400 349.880 1767.255 350.560 ;
        RECT 4.400 349.160 1763.200 349.880 ;
        RECT 1.445 348.480 1763.200 349.160 ;
        RECT 1.445 347.160 1767.255 348.480 ;
        RECT 4.400 345.760 1767.255 347.160 ;
        RECT 1.445 344.440 1767.255 345.760 ;
        RECT 1.445 343.760 1763.200 344.440 ;
        RECT 4.400 343.040 1763.200 343.760 ;
        RECT 4.400 342.360 1767.255 343.040 ;
        RECT 1.445 340.360 1767.255 342.360 ;
        RECT 4.400 339.000 1767.255 340.360 ;
        RECT 4.400 338.960 1763.200 339.000 ;
        RECT 1.445 337.600 1763.200 338.960 ;
        RECT 1.445 336.280 1767.255 337.600 ;
        RECT 4.400 334.880 1767.255 336.280 ;
        RECT 1.445 333.560 1767.255 334.880 ;
        RECT 1.445 332.880 1763.200 333.560 ;
        RECT 4.400 332.160 1763.200 332.880 ;
        RECT 4.400 331.480 1767.255 332.160 ;
        RECT 1.445 329.480 1767.255 331.480 ;
        RECT 4.400 328.120 1767.255 329.480 ;
        RECT 4.400 328.080 1763.200 328.120 ;
        RECT 1.445 326.720 1763.200 328.080 ;
        RECT 1.445 326.080 1767.255 326.720 ;
        RECT 4.400 324.680 1767.255 326.080 ;
        RECT 1.445 322.680 1767.255 324.680 ;
        RECT 4.400 321.280 1763.200 322.680 ;
        RECT 1.445 319.280 1767.255 321.280 ;
        RECT 4.400 317.880 1767.255 319.280 ;
        RECT 1.445 317.240 1767.255 317.880 ;
        RECT 1.445 315.840 1763.200 317.240 ;
        RECT 1.445 315.200 1767.255 315.840 ;
        RECT 4.400 313.800 1767.255 315.200 ;
        RECT 1.445 311.800 1767.255 313.800 ;
        RECT 4.400 310.400 1763.200 311.800 ;
        RECT 1.445 308.400 1767.255 310.400 ;
        RECT 4.400 307.000 1767.255 308.400 ;
        RECT 1.445 306.360 1767.255 307.000 ;
        RECT 1.445 305.000 1763.200 306.360 ;
        RECT 4.400 304.960 1763.200 305.000 ;
        RECT 4.400 303.600 1767.255 304.960 ;
        RECT 1.445 301.600 1767.255 303.600 ;
        RECT 4.400 300.920 1767.255 301.600 ;
        RECT 4.400 300.200 1763.200 300.920 ;
        RECT 1.445 299.520 1763.200 300.200 ;
        RECT 1.445 297.520 1767.255 299.520 ;
        RECT 4.400 296.120 1767.255 297.520 ;
        RECT 1.445 295.480 1767.255 296.120 ;
        RECT 1.445 294.120 1763.200 295.480 ;
        RECT 4.400 294.080 1763.200 294.120 ;
        RECT 4.400 292.720 1767.255 294.080 ;
        RECT 1.445 290.720 1767.255 292.720 ;
        RECT 4.400 290.040 1767.255 290.720 ;
        RECT 4.400 289.320 1763.200 290.040 ;
        RECT 1.445 288.640 1763.200 289.320 ;
        RECT 1.445 287.320 1767.255 288.640 ;
        RECT 4.400 285.920 1767.255 287.320 ;
        RECT 1.445 284.600 1767.255 285.920 ;
        RECT 1.445 283.920 1763.200 284.600 ;
        RECT 4.400 283.200 1763.200 283.920 ;
        RECT 4.400 282.520 1767.255 283.200 ;
        RECT 1.445 280.520 1767.255 282.520 ;
        RECT 4.400 279.160 1767.255 280.520 ;
        RECT 4.400 279.120 1763.200 279.160 ;
        RECT 1.445 277.760 1763.200 279.120 ;
        RECT 1.445 276.440 1767.255 277.760 ;
        RECT 4.400 275.040 1767.255 276.440 ;
        RECT 1.445 273.720 1767.255 275.040 ;
        RECT 1.445 273.040 1763.200 273.720 ;
        RECT 4.400 272.320 1763.200 273.040 ;
        RECT 4.400 271.640 1767.255 272.320 ;
        RECT 1.445 269.640 1767.255 271.640 ;
        RECT 4.400 268.280 1767.255 269.640 ;
        RECT 4.400 268.240 1763.200 268.280 ;
        RECT 1.445 266.880 1763.200 268.240 ;
        RECT 1.445 266.240 1767.255 266.880 ;
        RECT 4.400 264.840 1767.255 266.240 ;
        RECT 1.445 262.840 1767.255 264.840 ;
        RECT 4.400 261.440 1763.200 262.840 ;
        RECT 1.445 259.440 1767.255 261.440 ;
        RECT 4.400 258.040 1767.255 259.440 ;
        RECT 1.445 257.400 1767.255 258.040 ;
        RECT 1.445 256.000 1763.200 257.400 ;
        RECT 1.445 255.360 1767.255 256.000 ;
        RECT 4.400 253.960 1767.255 255.360 ;
        RECT 1.445 251.960 1767.255 253.960 ;
        RECT 4.400 250.560 1763.200 251.960 ;
        RECT 1.445 248.560 1767.255 250.560 ;
        RECT 4.400 247.160 1767.255 248.560 ;
        RECT 1.445 246.520 1767.255 247.160 ;
        RECT 1.445 245.160 1763.200 246.520 ;
        RECT 4.400 245.120 1763.200 245.160 ;
        RECT 4.400 243.760 1767.255 245.120 ;
        RECT 1.445 241.760 1767.255 243.760 ;
        RECT 4.400 241.080 1767.255 241.760 ;
        RECT 4.400 240.360 1763.200 241.080 ;
        RECT 1.445 239.680 1763.200 240.360 ;
        RECT 1.445 237.680 1767.255 239.680 ;
        RECT 4.400 236.280 1767.255 237.680 ;
        RECT 1.445 235.640 1767.255 236.280 ;
        RECT 1.445 234.280 1763.200 235.640 ;
        RECT 4.400 234.240 1763.200 234.280 ;
        RECT 4.400 232.880 1767.255 234.240 ;
        RECT 1.445 230.880 1767.255 232.880 ;
        RECT 4.400 230.200 1767.255 230.880 ;
        RECT 4.400 229.480 1763.200 230.200 ;
        RECT 1.445 228.800 1763.200 229.480 ;
        RECT 1.445 227.480 1767.255 228.800 ;
        RECT 4.400 226.080 1767.255 227.480 ;
        RECT 1.445 224.760 1767.255 226.080 ;
        RECT 1.445 224.080 1763.200 224.760 ;
        RECT 4.400 223.360 1763.200 224.080 ;
        RECT 4.400 222.680 1767.255 223.360 ;
        RECT 1.445 220.680 1767.255 222.680 ;
        RECT 4.400 219.320 1767.255 220.680 ;
        RECT 4.400 219.280 1763.200 219.320 ;
        RECT 1.445 217.920 1763.200 219.280 ;
        RECT 1.445 216.600 1767.255 217.920 ;
        RECT 4.400 215.200 1767.255 216.600 ;
        RECT 1.445 213.880 1767.255 215.200 ;
        RECT 1.445 213.200 1763.200 213.880 ;
        RECT 4.400 212.480 1763.200 213.200 ;
        RECT 4.400 211.800 1767.255 212.480 ;
        RECT 1.445 209.800 1767.255 211.800 ;
        RECT 4.400 208.440 1767.255 209.800 ;
        RECT 4.400 208.400 1763.200 208.440 ;
        RECT 1.445 207.040 1763.200 208.400 ;
        RECT 1.445 206.400 1767.255 207.040 ;
        RECT 4.400 205.000 1767.255 206.400 ;
        RECT 1.445 203.000 1767.255 205.000 ;
        RECT 4.400 201.600 1763.200 203.000 ;
        RECT 1.445 198.920 1767.255 201.600 ;
        RECT 4.400 198.240 1767.255 198.920 ;
        RECT 4.400 197.520 1763.200 198.240 ;
        RECT 1.445 196.840 1763.200 197.520 ;
        RECT 1.445 195.520 1767.255 196.840 ;
        RECT 4.400 194.120 1767.255 195.520 ;
        RECT 1.445 192.800 1767.255 194.120 ;
        RECT 1.445 192.120 1763.200 192.800 ;
        RECT 4.400 191.400 1763.200 192.120 ;
        RECT 4.400 190.720 1767.255 191.400 ;
        RECT 1.445 188.720 1767.255 190.720 ;
        RECT 4.400 187.360 1767.255 188.720 ;
        RECT 4.400 187.320 1763.200 187.360 ;
        RECT 1.445 185.960 1763.200 187.320 ;
        RECT 1.445 185.320 1767.255 185.960 ;
        RECT 4.400 183.920 1767.255 185.320 ;
        RECT 1.445 181.920 1767.255 183.920 ;
        RECT 4.400 180.520 1763.200 181.920 ;
        RECT 1.445 177.840 1767.255 180.520 ;
        RECT 4.400 176.480 1767.255 177.840 ;
        RECT 4.400 176.440 1763.200 176.480 ;
        RECT 1.445 175.080 1763.200 176.440 ;
        RECT 1.445 174.440 1767.255 175.080 ;
        RECT 4.400 173.040 1767.255 174.440 ;
        RECT 1.445 171.040 1767.255 173.040 ;
        RECT 4.400 169.640 1763.200 171.040 ;
        RECT 1.445 167.640 1767.255 169.640 ;
        RECT 4.400 166.240 1767.255 167.640 ;
        RECT 1.445 165.600 1767.255 166.240 ;
        RECT 1.445 164.240 1763.200 165.600 ;
        RECT 4.400 164.200 1763.200 164.240 ;
        RECT 4.400 162.840 1767.255 164.200 ;
        RECT 1.445 160.840 1767.255 162.840 ;
        RECT 4.400 160.160 1767.255 160.840 ;
        RECT 4.400 159.440 1763.200 160.160 ;
        RECT 1.445 158.760 1763.200 159.440 ;
        RECT 1.445 156.760 1767.255 158.760 ;
        RECT 4.400 155.360 1767.255 156.760 ;
        RECT 1.445 154.720 1767.255 155.360 ;
        RECT 1.445 153.360 1763.200 154.720 ;
        RECT 4.400 153.320 1763.200 153.360 ;
        RECT 4.400 151.960 1767.255 153.320 ;
        RECT 1.445 149.960 1767.255 151.960 ;
        RECT 4.400 149.280 1767.255 149.960 ;
        RECT 4.400 148.560 1763.200 149.280 ;
        RECT 1.445 147.880 1763.200 148.560 ;
        RECT 1.445 146.560 1767.255 147.880 ;
        RECT 4.400 145.160 1767.255 146.560 ;
        RECT 1.445 143.840 1767.255 145.160 ;
        RECT 1.445 143.160 1763.200 143.840 ;
        RECT 4.400 142.440 1763.200 143.160 ;
        RECT 4.400 141.760 1767.255 142.440 ;
        RECT 1.445 139.080 1767.255 141.760 ;
        RECT 4.400 138.400 1767.255 139.080 ;
        RECT 4.400 137.680 1763.200 138.400 ;
        RECT 1.445 137.000 1763.200 137.680 ;
        RECT 1.445 135.680 1767.255 137.000 ;
        RECT 4.400 134.280 1767.255 135.680 ;
        RECT 1.445 132.960 1767.255 134.280 ;
        RECT 1.445 132.280 1763.200 132.960 ;
        RECT 4.400 131.560 1763.200 132.280 ;
        RECT 4.400 130.880 1767.255 131.560 ;
        RECT 1.445 128.880 1767.255 130.880 ;
        RECT 4.400 127.520 1767.255 128.880 ;
        RECT 4.400 127.480 1763.200 127.520 ;
        RECT 1.445 126.120 1763.200 127.480 ;
        RECT 1.445 125.480 1767.255 126.120 ;
        RECT 4.400 124.080 1767.255 125.480 ;
        RECT 1.445 122.080 1767.255 124.080 ;
        RECT 4.400 120.680 1763.200 122.080 ;
        RECT 1.445 118.000 1767.255 120.680 ;
        RECT 4.400 116.640 1767.255 118.000 ;
        RECT 4.400 116.600 1763.200 116.640 ;
        RECT 1.445 115.240 1763.200 116.600 ;
        RECT 1.445 114.600 1767.255 115.240 ;
        RECT 4.400 113.200 1767.255 114.600 ;
        RECT 1.445 111.200 1767.255 113.200 ;
        RECT 4.400 109.800 1763.200 111.200 ;
        RECT 1.445 107.800 1767.255 109.800 ;
        RECT 4.400 106.400 1767.255 107.800 ;
        RECT 1.445 105.760 1767.255 106.400 ;
        RECT 1.445 104.400 1763.200 105.760 ;
        RECT 4.400 104.360 1763.200 104.400 ;
        RECT 4.400 103.000 1767.255 104.360 ;
        RECT 1.445 100.320 1767.255 103.000 ;
        RECT 4.400 98.920 1763.200 100.320 ;
        RECT 1.445 96.920 1767.255 98.920 ;
        RECT 4.400 95.520 1767.255 96.920 ;
        RECT 1.445 94.880 1767.255 95.520 ;
        RECT 1.445 93.520 1763.200 94.880 ;
        RECT 4.400 93.480 1763.200 93.520 ;
        RECT 4.400 92.120 1767.255 93.480 ;
        RECT 1.445 90.120 1767.255 92.120 ;
        RECT 4.400 89.440 1767.255 90.120 ;
        RECT 4.400 88.720 1763.200 89.440 ;
        RECT 1.445 88.040 1763.200 88.720 ;
        RECT 1.445 86.720 1767.255 88.040 ;
        RECT 4.400 85.320 1767.255 86.720 ;
        RECT 1.445 84.000 1767.255 85.320 ;
        RECT 1.445 83.320 1763.200 84.000 ;
        RECT 4.400 82.600 1763.200 83.320 ;
        RECT 4.400 81.920 1767.255 82.600 ;
        RECT 1.445 79.240 1767.255 81.920 ;
        RECT 4.400 78.560 1767.255 79.240 ;
        RECT 4.400 77.840 1763.200 78.560 ;
        RECT 1.445 77.160 1763.200 77.840 ;
        RECT 1.445 75.840 1767.255 77.160 ;
        RECT 4.400 74.440 1767.255 75.840 ;
        RECT 1.445 73.120 1767.255 74.440 ;
        RECT 1.445 72.440 1763.200 73.120 ;
        RECT 4.400 71.720 1763.200 72.440 ;
        RECT 4.400 71.040 1767.255 71.720 ;
        RECT 1.445 69.040 1767.255 71.040 ;
        RECT 4.400 67.680 1767.255 69.040 ;
        RECT 4.400 67.640 1763.200 67.680 ;
        RECT 1.445 66.280 1763.200 67.640 ;
        RECT 1.445 65.640 1767.255 66.280 ;
        RECT 4.400 64.240 1767.255 65.640 ;
        RECT 1.445 62.240 1767.255 64.240 ;
        RECT 4.400 60.840 1763.200 62.240 ;
        RECT 1.445 58.160 1767.255 60.840 ;
        RECT 4.400 56.800 1767.255 58.160 ;
        RECT 4.400 56.760 1763.200 56.800 ;
        RECT 1.445 55.400 1763.200 56.760 ;
        RECT 1.445 54.760 1767.255 55.400 ;
        RECT 4.400 53.360 1767.255 54.760 ;
        RECT 1.445 51.360 1767.255 53.360 ;
        RECT 4.400 49.960 1763.200 51.360 ;
        RECT 1.445 47.960 1767.255 49.960 ;
        RECT 4.400 46.560 1767.255 47.960 ;
        RECT 1.445 45.920 1767.255 46.560 ;
        RECT 1.445 44.560 1763.200 45.920 ;
        RECT 4.400 44.520 1763.200 44.560 ;
        RECT 4.400 43.160 1767.255 44.520 ;
        RECT 1.445 40.480 1767.255 43.160 ;
        RECT 4.400 39.080 1763.200 40.480 ;
        RECT 1.445 37.080 1767.255 39.080 ;
        RECT 4.400 35.680 1767.255 37.080 ;
        RECT 1.445 35.040 1767.255 35.680 ;
        RECT 1.445 33.680 1763.200 35.040 ;
        RECT 4.400 33.640 1763.200 33.680 ;
        RECT 4.400 32.280 1767.255 33.640 ;
        RECT 1.445 30.280 1767.255 32.280 ;
        RECT 4.400 29.600 1767.255 30.280 ;
        RECT 4.400 28.880 1763.200 29.600 ;
        RECT 1.445 28.200 1763.200 28.880 ;
        RECT 1.445 26.880 1767.255 28.200 ;
        RECT 4.400 25.480 1767.255 26.880 ;
        RECT 1.445 24.160 1767.255 25.480 ;
        RECT 1.445 23.480 1763.200 24.160 ;
        RECT 4.400 22.760 1763.200 23.480 ;
        RECT 4.400 22.080 1767.255 22.760 ;
        RECT 1.445 19.400 1767.255 22.080 ;
        RECT 4.400 18.720 1767.255 19.400 ;
        RECT 4.400 18.000 1763.200 18.720 ;
        RECT 1.445 17.320 1763.200 18.000 ;
        RECT 1.445 16.000 1767.255 17.320 ;
        RECT 4.400 14.600 1767.255 16.000 ;
        RECT 1.445 13.280 1767.255 14.600 ;
        RECT 1.445 12.600 1763.200 13.280 ;
        RECT 4.400 11.880 1763.200 12.600 ;
        RECT 4.400 11.200 1767.255 11.880 ;
        RECT 1.445 9.200 1767.255 11.200 ;
        RECT 4.400 7.840 1767.255 9.200 ;
        RECT 4.400 7.800 1763.200 7.840 ;
        RECT 1.445 6.440 1763.200 7.800 ;
        RECT 1.445 5.800 1767.255 6.440 ;
        RECT 4.400 4.400 1767.255 5.800 ;
        RECT 1.445 3.080 1767.255 4.400 ;
        RECT 1.445 2.400 1763.200 3.080 ;
        RECT 4.400 1.680 1763.200 2.400 ;
        RECT 4.400 1.535 1767.255 1.680 ;
      LAYER met4 ;
        RECT 3.975 1765.920 1767.025 1767.825 ;
        RECT 3.975 10.240 20.640 1765.920 ;
        RECT 23.040 10.240 97.440 1765.920 ;
        RECT 99.840 10.240 174.240 1765.920 ;
        RECT 176.640 10.240 251.040 1765.920 ;
        RECT 253.440 10.240 327.840 1765.920 ;
        RECT 330.240 10.240 404.640 1765.920 ;
        RECT 407.040 10.240 481.440 1765.920 ;
        RECT 483.840 10.240 558.240 1765.920 ;
        RECT 560.640 10.240 635.040 1765.920 ;
        RECT 637.440 10.240 711.840 1765.920 ;
        RECT 714.240 10.240 788.640 1765.920 ;
        RECT 791.040 10.240 865.440 1765.920 ;
        RECT 867.840 10.240 942.240 1765.920 ;
        RECT 944.640 10.240 1019.040 1765.920 ;
        RECT 1021.440 10.240 1095.840 1765.920 ;
        RECT 1098.240 10.240 1172.640 1765.920 ;
        RECT 1175.040 10.240 1249.440 1765.920 ;
        RECT 1251.840 10.240 1326.240 1765.920 ;
        RECT 1328.640 10.240 1403.040 1765.920 ;
        RECT 1405.440 10.240 1479.840 1765.920 ;
        RECT 1482.240 10.240 1556.640 1765.920 ;
        RECT 1559.040 10.240 1633.440 1765.920 ;
        RECT 1635.840 10.240 1710.240 1765.920 ;
        RECT 1712.640 10.240 1767.025 1765.920 ;
        RECT 3.975 9.695 1767.025 10.240 ;
  END
END Marmot
END LIBRARY

