VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Marmot
  CLASS BLOCK ;
  FOREIGN Marmot ;
  ORIGIN 0.000 0.000 ;
  SIZE 1756.625 BY 1767.345 ;
  PIN data_arrays_0_0_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1700.040 4.000 1700.640 ;
    END
  END data_arrays_0_0_ext_ram_addr1[0]
  PIN data_arrays_0_0_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1708.200 4.000 1708.800 ;
    END
  END data_arrays_0_0_ext_ram_addr1[1]
  PIN data_arrays_0_0_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.680 4.000 1716.280 ;
    END
  END data_arrays_0_0_ext_ram_addr1[2]
  PIN data_arrays_0_0_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.840 4.000 1724.440 ;
    END
  END data_arrays_0_0_ext_ram_addr1[3]
  PIN data_arrays_0_0_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1731.320 4.000 1731.920 ;
    END
  END data_arrays_0_0_ext_ram_addr1[4]
  PIN data_arrays_0_0_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1739.480 4.000 1740.080 ;
    END
  END data_arrays_0_0_ext_ram_addr1[5]
  PIN data_arrays_0_0_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1746.960 4.000 1747.560 ;
    END
  END data_arrays_0_0_ext_ram_addr1[6]
  PIN data_arrays_0_0_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1755.120 4.000 1755.720 ;
    END
  END data_arrays_0_0_ext_ram_addr1[7]
  PIN data_arrays_0_0_ext_ram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1762.600 4.000 1763.200 ;
    END
  END data_arrays_0_0_ext_ram_addr1[8]
  PIN data_arrays_0_0_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1004.400 4.000 1005.000 ;
    END
  END data_arrays_0_0_ext_ram_addr[0]
  PIN data_arrays_0_0_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END data_arrays_0_0_ext_ram_addr[1]
  PIN data_arrays_0_0_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END data_arrays_0_0_ext_ram_addr[2]
  PIN data_arrays_0_0_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1027.520 4.000 1028.120 ;
    END
  END data_arrays_0_0_ext_ram_addr[3]
  PIN data_arrays_0_0_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1035.680 4.000 1036.280 ;
    END
  END data_arrays_0_0_ext_ram_addr[4]
  PIN data_arrays_0_0_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.160 4.000 1043.760 ;
    END
  END data_arrays_0_0_ext_ram_addr[5]
  PIN data_arrays_0_0_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1051.320 4.000 1051.920 ;
    END
  END data_arrays_0_0_ext_ram_addr[6]
  PIN data_arrays_0_0_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1058.800 4.000 1059.400 ;
    END
  END data_arrays_0_0_ext_ram_addr[7]
  PIN data_arrays_0_0_ext_ram_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.960 4.000 1067.560 ;
    END
  END data_arrays_0_0_ext_ram_addr[8]
  PIN data_arrays_0_0_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END data_arrays_0_0_ext_ram_clk
  PIN data_arrays_0_0_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1637.480 4.000 1638.080 ;
    END
  END data_arrays_0_0_ext_ram_csb1[0]
  PIN data_arrays_0_0_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1645.640 4.000 1646.240 ;
    END
  END data_arrays_0_0_ext_ram_csb1[1]
  PIN data_arrays_0_0_ext_ram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1653.120 4.000 1653.720 ;
    END
  END data_arrays_0_0_ext_ram_csb1[2]
  PIN data_arrays_0_0_ext_ram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1661.280 4.000 1661.880 ;
    END
  END data_arrays_0_0_ext_ram_csb1[3]
  PIN data_arrays_0_0_ext_ram_csb1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1668.760 4.000 1669.360 ;
    END
  END data_arrays_0_0_ext_ram_csb1[4]
  PIN data_arrays_0_0_ext_ram_csb1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1676.920 4.000 1677.520 ;
    END
  END data_arrays_0_0_ext_ram_csb1[5]
  PIN data_arrays_0_0_ext_ram_csb1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1684.400 4.000 1685.000 ;
    END
  END data_arrays_0_0_ext_ram_csb1[6]
  PIN data_arrays_0_0_ext_ram_csb1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1692.560 4.000 1693.160 ;
    END
  END data_arrays_0_0_ext_ram_csb1[7]
  PIN data_arrays_0_0_ext_ram_csb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1598.720 4.000 1599.320 ;
    END
  END data_arrays_0_0_ext_ram_csb[0]
  PIN data_arrays_0_0_ext_ram_csb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1606.200 4.000 1606.800 ;
    END
  END data_arrays_0_0_ext_ram_csb[1]
  PIN data_arrays_0_0_ext_ram_csb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1614.360 4.000 1614.960 ;
    END
  END data_arrays_0_0_ext_ram_csb[2]
  PIN data_arrays_0_0_ext_ram_csb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1621.840 4.000 1622.440 ;
    END
  END data_arrays_0_0_ext_ram_csb[3]
  PIN data_arrays_0_0_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[0]
  PIN data_arrays_0_0_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[10]
  PIN data_arrays_0_0_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[11]
  PIN data_arrays_0_0_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[12]
  PIN data_arrays_0_0_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[13]
  PIN data_arrays_0_0_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[14]
  PIN data_arrays_0_0_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[15]
  PIN data_arrays_0_0_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[16]
  PIN data_arrays_0_0_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[17]
  PIN data_arrays_0_0_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[18]
  PIN data_arrays_0_0_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[19]
  PIN data_arrays_0_0_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[1]
  PIN data_arrays_0_0_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[20]
  PIN data_arrays_0_0_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[21]
  PIN data_arrays_0_0_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[22]
  PIN data_arrays_0_0_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[23]
  PIN data_arrays_0_0_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[24]
  PIN data_arrays_0_0_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[25]
  PIN data_arrays_0_0_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[26]
  PIN data_arrays_0_0_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[27]
  PIN data_arrays_0_0_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[28]
  PIN data_arrays_0_0_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[29]
  PIN data_arrays_0_0_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[2]
  PIN data_arrays_0_0_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[30]
  PIN data_arrays_0_0_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[31]
  PIN data_arrays_0_0_ext_ram_rdata0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[32]
  PIN data_arrays_0_0_ext_ram_rdata0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[33]
  PIN data_arrays_0_0_ext_ram_rdata0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[34]
  PIN data_arrays_0_0_ext_ram_rdata0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[35]
  PIN data_arrays_0_0_ext_ram_rdata0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[36]
  PIN data_arrays_0_0_ext_ram_rdata0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[37]
  PIN data_arrays_0_0_ext_ram_rdata0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[38]
  PIN data_arrays_0_0_ext_ram_rdata0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[39]
  PIN data_arrays_0_0_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[3]
  PIN data_arrays_0_0_ext_ram_rdata0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[40]
  PIN data_arrays_0_0_ext_ram_rdata0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[41]
  PIN data_arrays_0_0_ext_ram_rdata0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[42]
  PIN data_arrays_0_0_ext_ram_rdata0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[43]
  PIN data_arrays_0_0_ext_ram_rdata0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.520 4.000 348.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[44]
  PIN data_arrays_0_0_ext_ram_rdata0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[45]
  PIN data_arrays_0_0_ext_ram_rdata0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[46]
  PIN data_arrays_0_0_ext_ram_rdata0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[47]
  PIN data_arrays_0_0_ext_ram_rdata0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[48]
  PIN data_arrays_0_0_ext_ram_rdata0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[49]
  PIN data_arrays_0_0_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[4]
  PIN data_arrays_0_0_ext_ram_rdata0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[50]
  PIN data_arrays_0_0_ext_ram_rdata0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[51]
  PIN data_arrays_0_0_ext_ram_rdata0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[52]
  PIN data_arrays_0_0_ext_ram_rdata0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[53]
  PIN data_arrays_0_0_ext_ram_rdata0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[54]
  PIN data_arrays_0_0_ext_ram_rdata0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[55]
  PIN data_arrays_0_0_ext_ram_rdata0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[56]
  PIN data_arrays_0_0_ext_ram_rdata0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[57]
  PIN data_arrays_0_0_ext_ram_rdata0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[58]
  PIN data_arrays_0_0_ext_ram_rdata0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 464.480 4.000 465.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[59]
  PIN data_arrays_0_0_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[5]
  PIN data_arrays_0_0_ext_ram_rdata0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[60]
  PIN data_arrays_0_0_ext_ram_rdata0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[61]
  PIN data_arrays_0_0_ext_ram_rdata0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[62]
  PIN data_arrays_0_0_ext_ram_rdata0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.760 4.000 496.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[63]
  PIN data_arrays_0_0_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[6]
  PIN data_arrays_0_0_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[7]
  PIN data_arrays_0_0_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[8]
  PIN data_arrays_0_0_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[9]
  PIN data_arrays_0_0_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 4.000 504.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[0]
  PIN data_arrays_0_0_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[10]
  PIN data_arrays_0_0_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[11]
  PIN data_arrays_0_0_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[12]
  PIN data_arrays_0_0_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[13]
  PIN data_arrays_0_0_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[14]
  PIN data_arrays_0_0_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.880 4.000 621.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[15]
  PIN data_arrays_0_0_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[16]
  PIN data_arrays_0_0_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[17]
  PIN data_arrays_0_0_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[18]
  PIN data_arrays_0_0_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[19]
  PIN data_arrays_0_0_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[1]
  PIN data_arrays_0_0_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[20]
  PIN data_arrays_0_0_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[21]
  PIN data_arrays_0_0_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[22]
  PIN data_arrays_0_0_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[23]
  PIN data_arrays_0_0_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[24]
  PIN data_arrays_0_0_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[25]
  PIN data_arrays_0_0_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[26]
  PIN data_arrays_0_0_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.720 4.000 715.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[27]
  PIN data_arrays_0_0_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[28]
  PIN data_arrays_0_0_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[29]
  PIN data_arrays_0_0_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[2]
  PIN data_arrays_0_0_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[30]
  PIN data_arrays_0_0_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.000 4.000 746.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[31]
  PIN data_arrays_0_0_ext_ram_rdata1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.160 4.000 754.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[32]
  PIN data_arrays_0_0_ext_ram_rdata1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[33]
  PIN data_arrays_0_0_ext_ram_rdata1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[34]
  PIN data_arrays_0_0_ext_ram_rdata1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.280 4.000 777.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[35]
  PIN data_arrays_0_0_ext_ram_rdata1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[36]
  PIN data_arrays_0_0_ext_ram_rdata1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[37]
  PIN data_arrays_0_0_ext_ram_rdata1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[38]
  PIN data_arrays_0_0_ext_ram_rdata1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 808.560 4.000 809.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[39]
  PIN data_arrays_0_0_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[3]
  PIN data_arrays_0_0_ext_ram_rdata1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.720 4.000 817.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[40]
  PIN data_arrays_0_0_ext_ram_rdata1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.200 4.000 824.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[41]
  PIN data_arrays_0_0_ext_ram_rdata1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[42]
  PIN data_arrays_0_0_ext_ram_rdata1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[43]
  PIN data_arrays_0_0_ext_ram_rdata1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.000 4.000 848.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[44]
  PIN data_arrays_0_0_ext_ram_rdata1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[45]
  PIN data_arrays_0_0_ext_ram_rdata1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[46]
  PIN data_arrays_0_0_ext_ram_rdata1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.120 4.000 871.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[47]
  PIN data_arrays_0_0_ext_ram_rdata1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.280 4.000 879.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[48]
  PIN data_arrays_0_0_ext_ram_rdata1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.760 4.000 887.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[49]
  PIN data_arrays_0_0_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[4]
  PIN data_arrays_0_0_ext_ram_rdata1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.920 4.000 895.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[50]
  PIN data_arrays_0_0_ext_ram_rdata1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 902.400 4.000 903.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[51]
  PIN data_arrays_0_0_ext_ram_rdata1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 910.560 4.000 911.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[52]
  PIN data_arrays_0_0_ext_ram_rdata1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[53]
  PIN data_arrays_0_0_ext_ram_rdata1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.200 4.000 926.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[54]
  PIN data_arrays_0_0_ext_ram_rdata1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.680 4.000 934.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[55]
  PIN data_arrays_0_0_ext_ram_rdata1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[56]
  PIN data_arrays_0_0_ext_ram_rdata1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 949.320 4.000 949.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[57]
  PIN data_arrays_0_0_ext_ram_rdata1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 957.480 4.000 958.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[58]
  PIN data_arrays_0_0_ext_ram_rdata1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.960 4.000 965.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[59]
  PIN data_arrays_0_0_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[5]
  PIN data_arrays_0_0_ext_ram_rdata1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.120 4.000 973.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[60]
  PIN data_arrays_0_0_ext_ram_rdata1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[61]
  PIN data_arrays_0_0_ext_ram_rdata1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 988.760 4.000 989.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[62]
  PIN data_arrays_0_0_ext_ram_rdata1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[63]
  PIN data_arrays_0_0_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[6]
  PIN data_arrays_0_0_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[7]
  PIN data_arrays_0_0_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[8]
  PIN data_arrays_0_0_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[9]
  PIN data_arrays_0_0_ext_ram_rdata2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.430 1763.345 1186.710 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[0]
  PIN data_arrays_0_0_ext_ram_rdata2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 1763.345 1231.330 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[10]
  PIN data_arrays_0_0_ext_ram_rdata2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.650 1763.345 1235.930 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[11]
  PIN data_arrays_0_0_ext_ram_rdata2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 1763.345 1240.070 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[12]
  PIN data_arrays_0_0_ext_ram_rdata2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.390 1763.345 1244.670 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[13]
  PIN data_arrays_0_0_ext_ram_rdata2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990 1763.345 1249.270 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[14]
  PIN data_arrays_0_0_ext_ram_rdata2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 1763.345 1253.410 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[15]
  PIN data_arrays_0_0_ext_ram_rdata2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.730 1763.345 1258.010 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[16]
  PIN data_arrays_0_0_ext_ram_rdata2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 1763.345 1262.610 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[17]
  PIN data_arrays_0_0_ext_ram_rdata2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 1763.345 1267.210 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[18]
  PIN data_arrays_0_0_ext_ram_rdata2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.070 1763.345 1271.350 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[19]
  PIN data_arrays_0_0_ext_ram_rdata2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.570 1763.345 1190.850 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[1]
  PIN data_arrays_0_0_ext_ram_rdata2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.670 1763.345 1275.950 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[20]
  PIN data_arrays_0_0_ext_ram_rdata2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 1763.345 1280.550 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[21]
  PIN data_arrays_0_0_ext_ram_rdata2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.410 1763.345 1284.690 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[22]
  PIN data_arrays_0_0_ext_ram_rdata2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 1763.345 1289.290 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[23]
  PIN data_arrays_0_0_ext_ram_rdata2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.610 1763.345 1293.890 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[24]
  PIN data_arrays_0_0_ext_ram_rdata2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 1763.345 1298.490 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[25]
  PIN data_arrays_0_0_ext_ram_rdata2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.350 1763.345 1302.630 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[26]
  PIN data_arrays_0_0_ext_ram_rdata2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.950 1763.345 1307.230 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[27]
  PIN data_arrays_0_0_ext_ram_rdata2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.550 1763.345 1311.830 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[28]
  PIN data_arrays_0_0_ext_ram_rdata2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.690 1763.345 1315.970 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[29]
  PIN data_arrays_0_0_ext_ram_rdata2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 1763.345 1195.450 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[2]
  PIN data_arrays_0_0_ext_ram_rdata2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 1763.345 1320.570 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[30]
  PIN data_arrays_0_0_ext_ram_rdata2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.890 1763.345 1325.170 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[31]
  PIN data_arrays_0_0_ext_ram_rdata2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.490 1763.345 1329.770 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[32]
  PIN data_arrays_0_0_ext_ram_rdata2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 1763.345 1333.910 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[33]
  PIN data_arrays_0_0_ext_ram_rdata2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.230 1763.345 1338.510 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[34]
  PIN data_arrays_0_0_ext_ram_rdata2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 1763.345 1343.110 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[35]
  PIN data_arrays_0_0_ext_ram_rdata2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.970 1763.345 1347.250 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[36]
  PIN data_arrays_0_0_ext_ram_rdata2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.570 1763.345 1351.850 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[37]
  PIN data_arrays_0_0_ext_ram_rdata2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.170 1763.345 1356.450 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[38]
  PIN data_arrays_0_0_ext_ram_rdata2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 1763.345 1361.050 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[39]
  PIN data_arrays_0_0_ext_ram_rdata2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.770 1763.345 1200.050 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[3]
  PIN data_arrays_0_0_ext_ram_rdata2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.910 1763.345 1365.190 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[40]
  PIN data_arrays_0_0_ext_ram_rdata2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.510 1763.345 1369.790 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[41]
  PIN data_arrays_0_0_ext_ram_rdata2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.110 1763.345 1374.390 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[42]
  PIN data_arrays_0_0_ext_ram_rdata2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 1763.345 1378.990 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[43]
  PIN data_arrays_0_0_ext_ram_rdata2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.850 1763.345 1383.130 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[44]
  PIN data_arrays_0_0_ext_ram_rdata2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.450 1763.345 1387.730 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[45]
  PIN data_arrays_0_0_ext_ram_rdata2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.050 1763.345 1392.330 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[46]
  PIN data_arrays_0_0_ext_ram_rdata2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.190 1763.345 1396.470 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[47]
  PIN data_arrays_0_0_ext_ram_rdata2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 1763.345 1401.070 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[48]
  PIN data_arrays_0_0_ext_ram_rdata2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.390 1763.345 1405.670 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[49]
  PIN data_arrays_0_0_ext_ram_rdata2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 1763.345 1204.650 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[4]
  PIN data_arrays_0_0_ext_ram_rdata2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.990 1763.345 1410.270 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[50]
  PIN data_arrays_0_0_ext_ram_rdata2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.130 1763.345 1414.410 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[51]
  PIN data_arrays_0_0_ext_ram_rdata2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 1763.345 1419.010 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[52]
  PIN data_arrays_0_0_ext_ram_rdata2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 1763.345 1423.610 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[53]
  PIN data_arrays_0_0_ext_ram_rdata2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.470 1763.345 1427.750 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[54]
  PIN data_arrays_0_0_ext_ram_rdata2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.070 1763.345 1432.350 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[55]
  PIN data_arrays_0_0_ext_ram_rdata2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.670 1763.345 1436.950 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[56]
  PIN data_arrays_0_0_ext_ram_rdata2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.270 1763.345 1441.550 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[57]
  PIN data_arrays_0_0_ext_ram_rdata2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.410 1763.345 1445.690 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[58]
  PIN data_arrays_0_0_ext_ram_rdata2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.010 1763.345 1450.290 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[59]
  PIN data_arrays_0_0_ext_ram_rdata2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 1763.345 1208.790 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[5]
  PIN data_arrays_0_0_ext_ram_rdata2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.610 1763.345 1454.890 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[60]
  PIN data_arrays_0_0_ext_ram_rdata2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 1763.345 1459.030 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[61]
  PIN data_arrays_0_0_ext_ram_rdata2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.350 1763.345 1463.630 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[62]
  PIN data_arrays_0_0_ext_ram_rdata2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.950 1763.345 1468.230 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[63]
  PIN data_arrays_0_0_ext_ram_rdata2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.110 1763.345 1213.390 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[6]
  PIN data_arrays_0_0_ext_ram_rdata2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.710 1763.345 1217.990 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[7]
  PIN data_arrays_0_0_ext_ram_rdata2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.850 1763.345 1222.130 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[8]
  PIN data_arrays_0_0_ext_ram_rdata2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.450 1763.345 1226.730 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[9]
  PIN data_arrays_0_0_ext_ram_rdata3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.550 1763.345 1472.830 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[0]
  PIN data_arrays_0_0_ext_ram_rdata3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.170 1763.345 1517.450 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[10]
  PIN data_arrays_0_0_ext_ram_rdata3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.310 1763.345 1521.590 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[11]
  PIN data_arrays_0_0_ext_ram_rdata3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.910 1763.345 1526.190 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[12]
  PIN data_arrays_0_0_ext_ram_rdata3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.510 1763.345 1530.790 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[13]
  PIN data_arrays_0_0_ext_ram_rdata3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.110 1763.345 1535.390 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[14]
  PIN data_arrays_0_0_ext_ram_rdata3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 1763.345 1539.530 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[15]
  PIN data_arrays_0_0_ext_ram_rdata3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.850 1763.345 1544.130 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[16]
  PIN data_arrays_0_0_ext_ram_rdata3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.450 1763.345 1548.730 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[17]
  PIN data_arrays_0_0_ext_ram_rdata3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.590 1763.345 1552.870 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[18]
  PIN data_arrays_0_0_ext_ram_rdata3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 1763.345 1557.470 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[19]
  PIN data_arrays_0_0_ext_ram_rdata3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.690 1763.345 1476.970 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[1]
  PIN data_arrays_0_0_ext_ram_rdata3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 1763.345 1562.070 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[20]
  PIN data_arrays_0_0_ext_ram_rdata3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.390 1763.345 1566.670 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[21]
  PIN data_arrays_0_0_ext_ram_rdata3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.530 1763.345 1570.810 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[22]
  PIN data_arrays_0_0_ext_ram_rdata3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.130 1763.345 1575.410 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[23]
  PIN data_arrays_0_0_ext_ram_rdata3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.730 1763.345 1580.010 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[24]
  PIN data_arrays_0_0_ext_ram_rdata3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 1763.345 1584.610 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[25]
  PIN data_arrays_0_0_ext_ram_rdata3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.470 1763.345 1588.750 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[26]
  PIN data_arrays_0_0_ext_ram_rdata3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.070 1763.345 1593.350 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[27]
  PIN data_arrays_0_0_ext_ram_rdata3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.670 1763.345 1597.950 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[28]
  PIN data_arrays_0_0_ext_ram_rdata3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.810 1763.345 1602.090 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[29]
  PIN data_arrays_0_0_ext_ram_rdata3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 1763.345 1481.570 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[2]
  PIN data_arrays_0_0_ext_ram_rdata3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.410 1763.345 1606.690 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[30]
  PIN data_arrays_0_0_ext_ram_rdata3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.010 1763.345 1611.290 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[31]
  PIN data_arrays_0_0_ext_ram_rdata3[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.610 1763.345 1615.890 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[32]
  PIN data_arrays_0_0_ext_ram_rdata3[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.750 1763.345 1620.030 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[33]
  PIN data_arrays_0_0_ext_ram_rdata3[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.350 1763.345 1624.630 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[34]
  PIN data_arrays_0_0_ext_ram_rdata3[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.950 1763.345 1629.230 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[35]
  PIN data_arrays_0_0_ext_ram_rdata3[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.090 1763.345 1633.370 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[36]
  PIN data_arrays_0_0_ext_ram_rdata3[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1637.690 1763.345 1637.970 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[37]
  PIN data_arrays_0_0_ext_ram_rdata3[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 1763.345 1642.570 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[38]
  PIN data_arrays_0_0_ext_ram_rdata3[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.890 1763.345 1647.170 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[39]
  PIN data_arrays_0_0_ext_ram_rdata3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.890 1763.345 1486.170 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[3]
  PIN data_arrays_0_0_ext_ram_rdata3[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.030 1763.345 1651.310 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[40]
  PIN data_arrays_0_0_ext_ram_rdata3[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.630 1763.345 1655.910 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[41]
  PIN data_arrays_0_0_ext_ram_rdata3[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.230 1763.345 1660.510 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[42]
  PIN data_arrays_0_0_ext_ram_rdata3[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.370 1763.345 1664.650 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[43]
  PIN data_arrays_0_0_ext_ram_rdata3[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.970 1763.345 1669.250 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[44]
  PIN data_arrays_0_0_ext_ram_rdata3[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1673.570 1763.345 1673.850 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[45]
  PIN data_arrays_0_0_ext_ram_rdata3[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.170 1763.345 1678.450 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[46]
  PIN data_arrays_0_0_ext_ram_rdata3[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.310 1763.345 1682.590 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[47]
  PIN data_arrays_0_0_ext_ram_rdata3[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.910 1763.345 1687.190 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[48]
  PIN data_arrays_0_0_ext_ram_rdata3[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.510 1763.345 1691.790 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[49]
  PIN data_arrays_0_0_ext_ram_rdata3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.030 1763.345 1490.310 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[4]
  PIN data_arrays_0_0_ext_ram_rdata3[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1695.650 1763.345 1695.930 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[50]
  PIN data_arrays_0_0_ext_ram_rdata3[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 1763.345 1700.530 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[51]
  PIN data_arrays_0_0_ext_ram_rdata3[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.850 1763.345 1705.130 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[52]
  PIN data_arrays_0_0_ext_ram_rdata3[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.450 1763.345 1709.730 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[53]
  PIN data_arrays_0_0_ext_ram_rdata3[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.590 1763.345 1713.870 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[54]
  PIN data_arrays_0_0_ext_ram_rdata3[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 1763.345 1718.470 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[55]
  PIN data_arrays_0_0_ext_ram_rdata3[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.790 1763.345 1723.070 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[56]
  PIN data_arrays_0_0_ext_ram_rdata3[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.930 1763.345 1727.210 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[57]
  PIN data_arrays_0_0_ext_ram_rdata3[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.530 1763.345 1731.810 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[58]
  PIN data_arrays_0_0_ext_ram_rdata3[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.130 1763.345 1736.410 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[59]
  PIN data_arrays_0_0_ext_ram_rdata3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.630 1763.345 1494.910 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[5]
  PIN data_arrays_0_0_ext_ram_rdata3[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.730 1763.345 1741.010 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[60]
  PIN data_arrays_0_0_ext_ram_rdata3[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.870 1763.345 1745.150 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[61]
  PIN data_arrays_0_0_ext_ram_rdata3[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.470 1763.345 1749.750 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[62]
  PIN data_arrays_0_0_ext_ram_rdata3[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.070 1763.345 1754.350 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[63]
  PIN data_arrays_0_0_ext_ram_rdata3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.230 1763.345 1499.510 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[6]
  PIN data_arrays_0_0_ext_ram_rdata3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 1763.345 1504.110 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[7]
  PIN data_arrays_0_0_ext_ram_rdata3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.970 1763.345 1508.250 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[8]
  PIN data_arrays_0_0_ext_ram_rdata3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.570 1763.345 1512.850 1767.345 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[9]
  PIN data_arrays_0_0_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1082.600 4.000 1083.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[0]
  PIN data_arrays_0_0_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1160.800 4.000 1161.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[10]
  PIN data_arrays_0_0_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1168.280 4.000 1168.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata[11]
  PIN data_arrays_0_0_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata[12]
  PIN data_arrays_0_0_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.920 4.000 1184.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[13]
  PIN data_arrays_0_0_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1192.080 4.000 1192.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[14]
  PIN data_arrays_0_0_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1199.560 4.000 1200.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[15]
  PIN data_arrays_0_0_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.720 4.000 1208.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[16]
  PIN data_arrays_0_0_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1215.200 4.000 1215.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[17]
  PIN data_arrays_0_0_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1223.360 4.000 1223.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata[18]
  PIN data_arrays_0_0_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata[19]
  PIN data_arrays_0_0_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1090.080 4.000 1090.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[1]
  PIN data_arrays_0_0_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.000 4.000 1239.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[20]
  PIN data_arrays_0_0_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1246.480 4.000 1247.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[21]
  PIN data_arrays_0_0_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[22]
  PIN data_arrays_0_0_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1262.120 4.000 1262.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata[23]
  PIN data_arrays_0_0_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.280 4.000 1270.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata[24]
  PIN data_arrays_0_0_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1277.760 4.000 1278.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata[25]
  PIN data_arrays_0_0_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.920 4.000 1286.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[26]
  PIN data_arrays_0_0_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[27]
  PIN data_arrays_0_0_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1301.560 4.000 1302.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[28]
  PIN data_arrays_0_0_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.040 4.000 1309.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata[29]
  PIN data_arrays_0_0_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata[2]
  PIN data_arrays_0_0_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1317.200 4.000 1317.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[30]
  PIN data_arrays_0_0_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1324.680 4.000 1325.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata[31]
  PIN data_arrays_0_0_ext_ram_wdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata[32]
  PIN data_arrays_0_0_ext_ram_wdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1340.320 4.000 1340.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[33]
  PIN data_arrays_0_0_ext_ram_wdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1348.480 4.000 1349.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[34]
  PIN data_arrays_0_0_ext_ram_wdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1355.960 4.000 1356.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata[35]
  PIN data_arrays_0_0_ext_ram_wdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1364.120 4.000 1364.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata[36]
  PIN data_arrays_0_0_ext_ram_wdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1371.600 4.000 1372.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[37]
  PIN data_arrays_0_0_ext_ram_wdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1379.760 4.000 1380.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata[38]
  PIN data_arrays_0_0_ext_ram_wdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1387.240 4.000 1387.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata[39]
  PIN data_arrays_0_0_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.720 4.000 1106.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[3]
  PIN data_arrays_0_0_ext_ram_wdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1395.400 4.000 1396.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[40]
  PIN data_arrays_0_0_ext_ram_wdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1402.880 4.000 1403.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[41]
  PIN data_arrays_0_0_ext_ram_wdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata[42]
  PIN data_arrays_0_0_ext_ram_wdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1418.520 4.000 1419.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[43]
  PIN data_arrays_0_0_ext_ram_wdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1426.680 4.000 1427.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata[44]
  PIN data_arrays_0_0_ext_ram_wdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.160 4.000 1434.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[45]
  PIN data_arrays_0_0_ext_ram_wdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1442.320 4.000 1442.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[46]
  PIN data_arrays_0_0_ext_ram_wdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1449.800 4.000 1450.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[47]
  PIN data_arrays_0_0_ext_ram_wdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1457.960 4.000 1458.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata[48]
  PIN data_arrays_0_0_ext_ram_wdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata[49]
  PIN data_arrays_0_0_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1113.880 4.000 1114.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[4]
  PIN data_arrays_0_0_ext_ram_wdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1473.600 4.000 1474.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[50]
  PIN data_arrays_0_0_ext_ram_wdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1481.080 4.000 1481.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[51]
  PIN data_arrays_0_0_ext_ram_wdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata[52]
  PIN data_arrays_0_0_ext_ram_wdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1496.720 4.000 1497.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[53]
  PIN data_arrays_0_0_ext_ram_wdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1504.880 4.000 1505.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[54]
  PIN data_arrays_0_0_ext_ram_wdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1512.360 4.000 1512.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata[55]
  PIN data_arrays_0_0_ext_ram_wdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1520.520 4.000 1521.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[56]
  PIN data_arrays_0_0_ext_ram_wdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1528.000 4.000 1528.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[57]
  PIN data_arrays_0_0_ext_ram_wdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.160 4.000 1536.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[58]
  PIN data_arrays_0_0_ext_ram_wdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[59]
  PIN data_arrays_0_0_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1121.360 4.000 1121.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata[5]
  PIN data_arrays_0_0_ext_ram_wdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1551.800 4.000 1552.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[60]
  PIN data_arrays_0_0_ext_ram_wdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1559.280 4.000 1559.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata[61]
  PIN data_arrays_0_0_ext_ram_wdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1567.440 4.000 1568.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata[62]
  PIN data_arrays_0_0_ext_ram_wdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.920 4.000 1575.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[63]
  PIN data_arrays_0_0_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1129.520 4.000 1130.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[6]
  PIN data_arrays_0_0_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.000 4.000 1137.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[7]
  PIN data_arrays_0_0_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.160 4.000 1145.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[8]
  PIN data_arrays_0_0_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[9]
  PIN data_arrays_0_0_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1630.000 4.000 1630.600 ;
    END
  END data_arrays_0_0_ext_ram_web
  PIN data_arrays_0_0_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1583.080 4.000 1583.680 ;
    END
  END data_arrays_0_0_ext_ram_wmask[0]
  PIN data_arrays_0_0_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1590.560 4.000 1591.160 ;
    END
  END data_arrays_0_0_ext_ram_wmask[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 1763.345 677.030 1767.345 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 1763.345 810.890 1767.345 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1763.345 824.690 1767.345 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 1763.345 838.030 1767.345 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 1763.345 851.370 1767.345 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 1763.345 864.710 1767.345 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 1763.345 878.050 1767.345 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 1763.345 891.390 1767.345 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.450 1763.345 904.730 1767.345 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 1763.345 918.530 1767.345 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 1763.345 931.870 1767.345 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 1763.345 690.370 1767.345 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 1763.345 945.210 1767.345 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.270 1763.345 958.550 1767.345 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 1763.345 971.890 1767.345 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 1763.345 985.230 1767.345 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 1763.345 999.030 1767.345 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.090 1763.345 1012.370 1767.345 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.430 1763.345 1025.710 1767.345 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.770 1763.345 1039.050 1767.345 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 1763.345 1052.390 1767.345 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 1763.345 1065.730 1767.345 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 1763.345 703.710 1767.345 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 1763.345 1079.070 1767.345 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 1763.345 1092.870 1767.345 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.930 1763.345 1106.210 1767.345 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.270 1763.345 1119.550 1767.345 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.610 1763.345 1132.890 1767.345 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 1763.345 1146.230 1767.345 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 1763.345 1159.570 1767.345 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 1763.345 1173.370 1767.345 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 1763.345 717.050 1767.345 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 1763.345 730.390 1767.345 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 1763.345 744.190 1767.345 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 1763.345 757.530 1767.345 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 1763.345 770.870 1767.345 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 1763.345 784.210 1767.345 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 1763.345 797.550 1767.345 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 1763.345 681.630 1767.345 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 1763.345 815.490 1767.345 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 1763.345 828.830 1767.345 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 1763.345 842.170 1767.345 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 1763.345 855.970 1767.345 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 1763.345 869.310 1767.345 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 1763.345 882.650 1767.345 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 1763.345 895.990 1767.345 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 1763.345 909.330 1767.345 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 1763.345 922.670 1767.345 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 1763.345 936.010 1767.345 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 1763.345 694.970 1767.345 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 1763.345 949.810 1767.345 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 1763.345 963.150 1767.345 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 1763.345 976.490 1767.345 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 1763.345 989.830 1767.345 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 1763.345 1003.170 1767.345 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 1763.345 1016.510 1767.345 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.030 1763.345 1030.310 1767.345 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 1763.345 1043.650 1767.345 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 1763.345 1056.990 1767.345 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 1763.345 1070.330 1767.345 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 1763.345 708.310 1767.345 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.390 1763.345 1083.670 1767.345 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.730 1763.345 1097.010 1767.345 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 1763.345 1110.350 1767.345 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 1763.345 1124.150 1767.345 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 1763.345 1137.490 1767.345 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.550 1763.345 1150.830 1767.345 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 1763.345 1164.170 1767.345 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 1763.345 1177.510 1767.345 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1763.345 721.650 1767.345 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 1763.345 734.990 1767.345 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 1763.345 748.330 1767.345 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 1763.345 761.670 1767.345 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 1763.345 775.470 1767.345 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 1763.345 788.810 1767.345 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 1763.345 802.150 1767.345 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 1763.345 685.770 1767.345 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 1763.345 820.090 1767.345 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 1763.345 833.430 1767.345 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 1763.345 846.770 1767.345 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 1763.345 860.110 1767.345 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 1763.345 873.450 1767.345 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 1763.345 887.250 1767.345 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 1763.345 900.590 1767.345 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 1763.345 913.930 1767.345 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 1763.345 927.270 1767.345 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 1763.345 940.610 1767.345 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 1763.345 699.110 1767.345 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 1763.345 953.950 1767.345 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.010 1763.345 967.290 1767.345 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 1763.345 981.090 1767.345 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 1763.345 994.430 1767.345 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 1763.345 1007.770 1767.345 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 1763.345 1021.110 1767.345 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 1763.345 1034.450 1767.345 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 1763.345 1047.790 1767.345 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 1763.345 1061.590 1767.345 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.650 1763.345 1074.930 1767.345 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 1763.345 712.910 1767.345 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.990 1763.345 1088.270 1767.345 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 1763.345 1101.610 1767.345 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.670 1763.345 1114.950 1767.345 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 1763.345 1128.290 1767.345 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 1763.345 1141.630 1767.345 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.150 1763.345 1155.430 1767.345 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.490 1763.345 1168.770 1767.345 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 1763.345 1182.110 1767.345 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 1763.345 726.250 1767.345 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 1763.345 739.590 1767.345 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 1763.345 752.930 1767.345 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 1763.345 766.270 1767.345 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1763.345 779.610 1767.345 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 1763.345 793.410 1767.345 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 1763.345 806.750 1767.345 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 0.000 1747.450 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.850 0.000 1751.130 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.530 0.000 1754.810 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.170 0.000 1448.450 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 0.000 1459.030 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1469.330 0.000 1469.610 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.910 0.000 1480.190 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.530 0.000 1501.810 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.110 0.000 1512.390 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.690 0.000 1522.970 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.270 0.000 1533.550 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.310 0.000 1544.590 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.890 0.000 1555.170 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.470 0.000 1565.750 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.050 0.000 1576.330 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.090 0.000 1587.370 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.670 0.000 1597.950 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.250 0.000 1608.530 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.830 0.000 1619.110 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.870 0.000 1630.150 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.450 0.000 1640.730 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.030 0.000 1651.310 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 0.000 1661.890 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.650 0.000 1672.930 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.230 0.000 1683.510 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.390 0.000 1704.670 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.430 0.000 1715.710 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 0.000 1726.290 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.590 0.000 1736.870 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 0.000 753.390 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 0.000 774.550 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 0.000 806.750 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.250 0.000 849.530 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.010 0.000 967.290 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.590 0.000 977.870 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 0.000 988.450 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 0.000 999.490 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.370 0.000 1020.650 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 0.000 1031.230 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.530 0.000 1041.810 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.570 0.000 1052.850 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.150 0.000 1063.430 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 0.000 1074.010 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 0.000 1084.590 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 0.000 1095.630 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.930 0.000 1106.210 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 0.000 1116.790 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.710 0.000 1148.990 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 0.000 1170.150 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 0.000 1191.770 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 0.000 1202.350 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.650 0.000 1212.930 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.270 0.000 1234.550 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.850 0.000 1245.130 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.430 0.000 1255.710 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.050 0.000 1277.330 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.630 0.000 1287.910 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 0.000 1298.490 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.790 0.000 1309.070 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.830 0.000 1320.110 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 0.000 1330.690 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 0.000 1341.270 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.570 0.000 1351.850 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.610 0.000 1362.890 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.190 0.000 1373.470 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.770 0.000 1384.050 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.390 0.000 1405.670 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.970 0.000 1416.250 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 0.000 1426.830 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.130 0.000 1437.410 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.390 0.000 1451.670 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.430 0.000 1462.710 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.010 0.000 1473.290 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.590 0.000 1483.870 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 0.000 1494.450 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1505.210 0.000 1505.490 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.790 0.000 1516.070 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 0.000 1526.650 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.950 0.000 1537.230 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.530 0.000 1547.810 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 0.000 1558.850 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.150 0.000 1569.430 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.730 0.000 1580.010 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.310 0.000 1590.590 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.350 0.000 1601.630 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.930 0.000 1612.210 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.510 0.000 1622.790 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.090 0.000 1633.370 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.130 0.000 1644.410 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.710 0.000 1654.990 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.290 0.000 1665.570 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.870 0.000 1676.150 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.910 0.000 1687.190 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.490 0.000 1697.770 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.070 0.000 1708.350 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.650 0.000 1718.930 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.690 0.000 1729.970 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.270 0.000 1740.550 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 0.000 639.310 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 0.000 703.710 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 0.000 735.450 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 0.000 746.490 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.570 0.000 799.850 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 0.000 821.010 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 0.000 842.630 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 0.000 874.370 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 0.000 885.410 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.290 0.000 906.570 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 0.000 928.190 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 0.000 938.770 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 0.000 949.350 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.690 0.000 970.970 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 0.000 981.550 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.630 0.000 1034.910 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.210 0.000 1045.490 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.830 0.000 1067.110 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.410 0.000 1077.690 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.990 0.000 1088.270 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.770 0.000 1131.050 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 0.000 1141.630 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.390 0.000 1152.670 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.970 0.000 1163.250 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.550 0.000 1173.830 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.130 0.000 1184.410 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.750 0.000 1206.030 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.330 0.000 1216.610 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.950 0.000 1238.230 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.530 0.000 1248.810 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 0.000 1259.390 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 0.000 1269.970 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 0.000 1280.550 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.890 0.000 1302.170 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.470 0.000 1312.750 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 0.000 1323.330 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.090 0.000 1334.370 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.670 0.000 1344.950 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.250 0.000 1355.530 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.830 0.000 1366.110 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.870 0.000 1377.150 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.450 0.000 1387.730 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.030 0.000 1398.310 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.610 0.000 1408.890 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.650 0.000 1419.930 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1430.230 0.000 1430.510 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.810 0.000 1441.090 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.070 0.000 1455.350 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.650 0.000 1465.930 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.690 0.000 1476.970 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.270 0.000 1487.550 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.850 0.000 1498.130 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.430 0.000 1508.710 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.010 0.000 1519.290 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.050 0.000 1530.330 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.630 0.000 1540.910 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.210 0.000 1551.490 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 0.000 1562.070 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.830 0.000 1573.110 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.410 0.000 1583.690 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.990 0.000 1594.270 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.570 0.000 1604.850 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.610 0.000 1615.890 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.190 0.000 1626.470 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.770 0.000 1637.050 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.350 0.000 1647.630 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 0.000 1658.670 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.970 0.000 1669.250 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.550 0.000 1679.830 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.130 0.000 1690.410 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1701.170 0.000 1701.450 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.750 0.000 1712.030 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.330 0.000 1722.610 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.910 0.000 1733.190 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.950 0.000 1744.230 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 0.000 781.910 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 0.000 803.070 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 0.000 835.270 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.190 0.000 867.470 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 0.000 878.050 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.970 0.000 910.250 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 0.000 920.830 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 0.000 931.410 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 0.000 953.030 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 0.000 963.610 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.910 0.000 974.190 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.530 0.000 995.810 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.110 0.000 1006.390 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 0.000 1038.590 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 0.000 1049.170 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 0.000 1070.330 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.090 0.000 1081.370 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 0.000 1091.950 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.830 0.000 1113.110 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.610 0.000 1155.890 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.650 0.000 1166.930 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 0.000 1177.510 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 0.000 1188.090 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 0.000 1198.670 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.430 0.000 1209.710 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.010 0.000 1220.290 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.590 0.000 1230.870 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.210 0.000 1252.490 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.790 0.000 1263.070 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.370 0.000 1273.650 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.950 0.000 1284.230 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.570 0.000 1305.850 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 0.000 1316.430 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.310 0.000 1337.590 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.510 0.000 1369.790 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 0.000 1380.370 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.710 0.000 1401.990 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.290 0.000 1412.570 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.910 0.000 1434.190 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.490 0.000 1444.770 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END la_oenb[9]
  PIN tag_array_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 1763.345 498.090 1767.345 ;
    END
  END tag_array_ext_ram_addr1[0]
  PIN tag_array_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 1763.345 502.690 1767.345 ;
    END
  END tag_array_ext_ram_addr1[1]
  PIN tag_array_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 1763.345 507.290 1767.345 ;
    END
  END tag_array_ext_ram_addr1[2]
  PIN tag_array_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 1763.345 511.430 1767.345 ;
    END
  END tag_array_ext_ram_addr1[3]
  PIN tag_array_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 1763.345 516.030 1767.345 ;
    END
  END tag_array_ext_ram_addr1[4]
  PIN tag_array_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 1763.345 520.630 1767.345 ;
    END
  END tag_array_ext_ram_addr1[5]
  PIN tag_array_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 1763.345 524.770 1767.345 ;
    END
  END tag_array_ext_ram_addr1[6]
  PIN tag_array_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 1763.345 529.370 1767.345 ;
    END
  END tag_array_ext_ram_addr1[7]
  PIN tag_array_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 1763.345 144.810 1767.345 ;
    END
  END tag_array_ext_ram_addr[0]
  PIN tag_array_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 1763.345 149.410 1767.345 ;
    END
  END tag_array_ext_ram_addr[1]
  PIN tag_array_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 1763.345 154.010 1767.345 ;
    END
  END tag_array_ext_ram_addr[2]
  PIN tag_array_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 1763.345 158.610 1767.345 ;
    END
  END tag_array_ext_ram_addr[3]
  PIN tag_array_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 1763.345 162.750 1767.345 ;
    END
  END tag_array_ext_ram_addr[4]
  PIN tag_array_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 1763.345 167.350 1767.345 ;
    END
  END tag_array_ext_ram_addr[5]
  PIN tag_array_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 1763.345 171.950 1767.345 ;
    END
  END tag_array_ext_ram_addr[6]
  PIN tag_array_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 1763.345 176.090 1767.345 ;
    END
  END tag_array_ext_ram_addr[7]
  PIN tag_array_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1763.345 180.690 1767.345 ;
    END
  END tag_array_ext_ram_clk
  PIN tag_array_ext_ram_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1763.345 480.150 1767.345 ;
    END
  END tag_array_ext_ram_csb
  PIN tag_array_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 1763.345 489.350 1767.345 ;
    END
  END tag_array_ext_ram_csb1[0]
  PIN tag_array_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 1763.345 493.490 1767.345 ;
    END
  END tag_array_ext_ram_csb1[1]
  PIN tag_array_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 1763.345 2.210 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[0]
  PIN tag_array_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 1763.345 46.830 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[10]
  PIN tag_array_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 1763.345 50.970 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[11]
  PIN tag_array_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 1763.345 55.570 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[12]
  PIN tag_array_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 1763.345 60.170 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[13]
  PIN tag_array_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1763.345 64.770 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[14]
  PIN tag_array_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 1763.345 68.910 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[15]
  PIN tag_array_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 1763.345 73.510 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[16]
  PIN tag_array_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 1763.345 78.110 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[17]
  PIN tag_array_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 1763.345 82.250 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[18]
  PIN tag_array_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 1763.345 86.850 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[19]
  PIN tag_array_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 1763.345 6.350 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[1]
  PIN tag_array_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 1763.345 91.450 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[20]
  PIN tag_array_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 1763.345 96.050 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[21]
  PIN tag_array_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1763.345 100.190 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[22]
  PIN tag_array_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 1763.345 104.790 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[23]
  PIN tag_array_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 1763.345 109.390 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[24]
  PIN tag_array_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 1763.345 113.530 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[25]
  PIN tag_array_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 1763.345 118.130 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[26]
  PIN tag_array_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1763.345 122.730 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[27]
  PIN tag_array_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 1763.345 127.330 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[28]
  PIN tag_array_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 1763.345 131.470 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[29]
  PIN tag_array_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 1763.345 10.950 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[2]
  PIN tag_array_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 1763.345 136.070 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[30]
  PIN tag_array_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 1763.345 140.670 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[31]
  PIN tag_array_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 1763.345 15.550 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[3]
  PIN tag_array_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1763.345 19.690 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[4]
  PIN tag_array_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 1763.345 24.290 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[5]
  PIN tag_array_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 1763.345 28.890 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[6]
  PIN tag_array_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 1763.345 33.490 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[7]
  PIN tag_array_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 1763.345 37.630 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[8]
  PIN tag_array_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 1763.345 42.230 1767.345 ;
    END
  END tag_array_ext_ram_rdata0[9]
  PIN tag_array_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 1763.345 533.970 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[0]
  PIN tag_array_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 1763.345 578.590 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[10]
  PIN tag_array_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 1763.345 583.190 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[11]
  PIN tag_array_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 1763.345 587.790 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[12]
  PIN tag_array_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 1763.345 591.930 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[13]
  PIN tag_array_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 1763.345 596.530 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[14]
  PIN tag_array_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 1763.345 601.130 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[15]
  PIN tag_array_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 1763.345 605.270 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[16]
  PIN tag_array_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 1763.345 609.870 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[17]
  PIN tag_array_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 1763.345 614.470 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[18]
  PIN tag_array_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 1763.345 619.070 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[19]
  PIN tag_array_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 1763.345 538.570 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[1]
  PIN tag_array_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 1763.345 623.210 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[20]
  PIN tag_array_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 1763.345 627.810 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[21]
  PIN tag_array_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 1763.345 632.410 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[22]
  PIN tag_array_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 1763.345 636.550 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[23]
  PIN tag_array_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 1763.345 641.150 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[24]
  PIN tag_array_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 1763.345 645.750 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[25]
  PIN tag_array_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 1763.345 650.350 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[26]
  PIN tag_array_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 1763.345 654.490 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[27]
  PIN tag_array_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 1763.345 659.090 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[28]
  PIN tag_array_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 1763.345 663.690 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[29]
  PIN tag_array_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 1763.345 542.710 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[2]
  PIN tag_array_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 1763.345 667.830 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[30]
  PIN tag_array_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 1763.345 672.430 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[31]
  PIN tag_array_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 1763.345 547.310 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[3]
  PIN tag_array_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 1763.345 551.910 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[4]
  PIN tag_array_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 1763.345 556.050 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[5]
  PIN tag_array_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1763.345 560.650 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[6]
  PIN tag_array_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 1763.345 565.250 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[7]
  PIN tag_array_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 1763.345 569.850 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[8]
  PIN tag_array_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 1763.345 573.990 1767.345 ;
    END
  END tag_array_ext_ram_rdata1[9]
  PIN tag_array_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 1763.345 185.290 1767.345 ;
    END
  END tag_array_ext_ram_wdata[0]
  PIN tag_array_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 1763.345 229.910 1767.345 ;
    END
  END tag_array_ext_ram_wdata[10]
  PIN tag_array_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 1763.345 234.510 1767.345 ;
    END
  END tag_array_ext_ram_wdata[11]
  PIN tag_array_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 1763.345 239.110 1767.345 ;
    END
  END tag_array_ext_ram_wdata[12]
  PIN tag_array_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 1763.345 243.250 1767.345 ;
    END
  END tag_array_ext_ram_wdata[13]
  PIN tag_array_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 1763.345 247.850 1767.345 ;
    END
  END tag_array_ext_ram_wdata[14]
  PIN tag_array_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 1763.345 252.450 1767.345 ;
    END
  END tag_array_ext_ram_wdata[15]
  PIN tag_array_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 1763.345 256.590 1767.345 ;
    END
  END tag_array_ext_ram_wdata[16]
  PIN tag_array_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 1763.345 261.190 1767.345 ;
    END
  END tag_array_ext_ram_wdata[17]
  PIN tag_array_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 1763.345 265.790 1767.345 ;
    END
  END tag_array_ext_ram_wdata[18]
  PIN tag_array_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 1763.345 270.390 1767.345 ;
    END
  END tag_array_ext_ram_wdata[19]
  PIN tag_array_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 1763.345 189.890 1767.345 ;
    END
  END tag_array_ext_ram_wdata[1]
  PIN tag_array_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 1763.345 274.530 1767.345 ;
    END
  END tag_array_ext_ram_wdata[20]
  PIN tag_array_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 1763.345 279.130 1767.345 ;
    END
  END tag_array_ext_ram_wdata[21]
  PIN tag_array_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1763.345 283.730 1767.345 ;
    END
  END tag_array_ext_ram_wdata[22]
  PIN tag_array_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 1763.345 287.870 1767.345 ;
    END
  END tag_array_ext_ram_wdata[23]
  PIN tag_array_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 1763.345 292.470 1767.345 ;
    END
  END tag_array_ext_ram_wdata[24]
  PIN tag_array_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 1763.345 297.070 1767.345 ;
    END
  END tag_array_ext_ram_wdata[25]
  PIN tag_array_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 1763.345 301.670 1767.345 ;
    END
  END tag_array_ext_ram_wdata[26]
  PIN tag_array_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 1763.345 305.810 1767.345 ;
    END
  END tag_array_ext_ram_wdata[27]
  PIN tag_array_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 1763.345 310.410 1767.345 ;
    END
  END tag_array_ext_ram_wdata[28]
  PIN tag_array_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 1763.345 315.010 1767.345 ;
    END
  END tag_array_ext_ram_wdata[29]
  PIN tag_array_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 1763.345 194.030 1767.345 ;
    END
  END tag_array_ext_ram_wdata[2]
  PIN tag_array_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 1763.345 319.150 1767.345 ;
    END
  END tag_array_ext_ram_wdata[30]
  PIN tag_array_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 1763.345 323.750 1767.345 ;
    END
  END tag_array_ext_ram_wdata[31]
  PIN tag_array_ext_ram_wdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 1763.345 328.350 1767.345 ;
    END
  END tag_array_ext_ram_wdata[32]
  PIN tag_array_ext_ram_wdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 1763.345 332.950 1767.345 ;
    END
  END tag_array_ext_ram_wdata[33]
  PIN tag_array_ext_ram_wdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 1763.345 337.090 1767.345 ;
    END
  END tag_array_ext_ram_wdata[34]
  PIN tag_array_ext_ram_wdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 1763.345 341.690 1767.345 ;
    END
  END tag_array_ext_ram_wdata[35]
  PIN tag_array_ext_ram_wdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 1763.345 346.290 1767.345 ;
    END
  END tag_array_ext_ram_wdata[36]
  PIN tag_array_ext_ram_wdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 1763.345 350.430 1767.345 ;
    END
  END tag_array_ext_ram_wdata[37]
  PIN tag_array_ext_ram_wdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 1763.345 355.030 1767.345 ;
    END
  END tag_array_ext_ram_wdata[38]
  PIN tag_array_ext_ram_wdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 1763.345 359.630 1767.345 ;
    END
  END tag_array_ext_ram_wdata[39]
  PIN tag_array_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 1763.345 198.630 1767.345 ;
    END
  END tag_array_ext_ram_wdata[3]
  PIN tag_array_ext_ram_wdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1763.345 364.230 1767.345 ;
    END
  END tag_array_ext_ram_wdata[40]
  PIN tag_array_ext_ram_wdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 1763.345 368.370 1767.345 ;
    END
  END tag_array_ext_ram_wdata[41]
  PIN tag_array_ext_ram_wdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 1763.345 372.970 1767.345 ;
    END
  END tag_array_ext_ram_wdata[42]
  PIN tag_array_ext_ram_wdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 1763.345 377.570 1767.345 ;
    END
  END tag_array_ext_ram_wdata[43]
  PIN tag_array_ext_ram_wdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 1763.345 381.710 1767.345 ;
    END
  END tag_array_ext_ram_wdata[44]
  PIN tag_array_ext_ram_wdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 1763.345 386.310 1767.345 ;
    END
  END tag_array_ext_ram_wdata[45]
  PIN tag_array_ext_ram_wdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 1763.345 390.910 1767.345 ;
    END
  END tag_array_ext_ram_wdata[46]
  PIN tag_array_ext_ram_wdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 1763.345 395.510 1767.345 ;
    END
  END tag_array_ext_ram_wdata[47]
  PIN tag_array_ext_ram_wdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1763.345 399.650 1767.345 ;
    END
  END tag_array_ext_ram_wdata[48]
  PIN tag_array_ext_ram_wdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 1763.345 404.250 1767.345 ;
    END
  END tag_array_ext_ram_wdata[49]
  PIN tag_array_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 1763.345 203.230 1767.345 ;
    END
  END tag_array_ext_ram_wdata[4]
  PIN tag_array_ext_ram_wdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 1763.345 408.850 1767.345 ;
    END
  END tag_array_ext_ram_wdata[50]
  PIN tag_array_ext_ram_wdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 1763.345 413.450 1767.345 ;
    END
  END tag_array_ext_ram_wdata[51]
  PIN tag_array_ext_ram_wdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 1763.345 417.590 1767.345 ;
    END
  END tag_array_ext_ram_wdata[52]
  PIN tag_array_ext_ram_wdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 1763.345 422.190 1767.345 ;
    END
  END tag_array_ext_ram_wdata[53]
  PIN tag_array_ext_ram_wdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 1763.345 426.790 1767.345 ;
    END
  END tag_array_ext_ram_wdata[54]
  PIN tag_array_ext_ram_wdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 1763.345 430.930 1767.345 ;
    END
  END tag_array_ext_ram_wdata[55]
  PIN tag_array_ext_ram_wdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 1763.345 435.530 1767.345 ;
    END
  END tag_array_ext_ram_wdata[56]
  PIN tag_array_ext_ram_wdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 1763.345 440.130 1767.345 ;
    END
  END tag_array_ext_ram_wdata[57]
  PIN tag_array_ext_ram_wdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 1763.345 444.730 1767.345 ;
    END
  END tag_array_ext_ram_wdata[58]
  PIN tag_array_ext_ram_wdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 1763.345 448.870 1767.345 ;
    END
  END tag_array_ext_ram_wdata[59]
  PIN tag_array_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 1763.345 207.830 1767.345 ;
    END
  END tag_array_ext_ram_wdata[5]
  PIN tag_array_ext_ram_wdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 1763.345 453.470 1767.345 ;
    END
  END tag_array_ext_ram_wdata[60]
  PIN tag_array_ext_ram_wdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 1763.345 458.070 1767.345 ;
    END
  END tag_array_ext_ram_wdata[61]
  PIN tag_array_ext_ram_wdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 1763.345 462.210 1767.345 ;
    END
  END tag_array_ext_ram_wdata[62]
  PIN tag_array_ext_ram_wdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 1763.345 466.810 1767.345 ;
    END
  END tag_array_ext_ram_wdata[63]
  PIN tag_array_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 1763.345 211.970 1767.345 ;
    END
  END tag_array_ext_ram_wdata[6]
  PIN tag_array_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 1763.345 216.570 1767.345 ;
    END
  END tag_array_ext_ram_wdata[7]
  PIN tag_array_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 1763.345 221.170 1767.345 ;
    END
  END tag_array_ext_ram_wdata[8]
  PIN tag_array_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 1763.345 225.310 1767.345 ;
    END
  END tag_array_ext_ram_wdata[9]
  PIN tag_array_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 1763.345 484.750 1767.345 ;
    END
  END tag_array_ext_ram_web
  PIN tag_array_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 1763.345 471.410 1767.345 ;
    END
  END tag_array_ext_ram_wmask[0]
  PIN tag_array_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 1763.345 476.010 1767.345 ;
    END
  END tag_array_ext_ram_wmask[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1754.640 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1754.640 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1750.760 1754.485 ;
      LAYER met1 ;
        RECT 1.450 6.160 1754.830 1767.280 ;
      LAYER met2 ;
        RECT 1.480 1763.065 1.650 1767.310 ;
        RECT 2.490 1763.065 5.790 1767.310 ;
        RECT 6.630 1763.065 10.390 1767.310 ;
        RECT 11.230 1763.065 14.990 1767.310 ;
        RECT 15.830 1763.065 19.130 1767.310 ;
        RECT 19.970 1763.065 23.730 1767.310 ;
        RECT 24.570 1763.065 28.330 1767.310 ;
        RECT 29.170 1763.065 32.930 1767.310 ;
        RECT 33.770 1763.065 37.070 1767.310 ;
        RECT 37.910 1763.065 41.670 1767.310 ;
        RECT 42.510 1763.065 46.270 1767.310 ;
        RECT 47.110 1763.065 50.410 1767.310 ;
        RECT 51.250 1763.065 55.010 1767.310 ;
        RECT 55.850 1763.065 59.610 1767.310 ;
        RECT 60.450 1763.065 64.210 1767.310 ;
        RECT 65.050 1763.065 68.350 1767.310 ;
        RECT 69.190 1763.065 72.950 1767.310 ;
        RECT 73.790 1763.065 77.550 1767.310 ;
        RECT 78.390 1763.065 81.690 1767.310 ;
        RECT 82.530 1763.065 86.290 1767.310 ;
        RECT 87.130 1763.065 90.890 1767.310 ;
        RECT 91.730 1763.065 95.490 1767.310 ;
        RECT 96.330 1763.065 99.630 1767.310 ;
        RECT 100.470 1763.065 104.230 1767.310 ;
        RECT 105.070 1763.065 108.830 1767.310 ;
        RECT 109.670 1763.065 112.970 1767.310 ;
        RECT 113.810 1763.065 117.570 1767.310 ;
        RECT 118.410 1763.065 122.170 1767.310 ;
        RECT 123.010 1763.065 126.770 1767.310 ;
        RECT 127.610 1763.065 130.910 1767.310 ;
        RECT 131.750 1763.065 135.510 1767.310 ;
        RECT 136.350 1763.065 140.110 1767.310 ;
        RECT 140.950 1763.065 144.250 1767.310 ;
        RECT 145.090 1763.065 148.850 1767.310 ;
        RECT 149.690 1763.065 153.450 1767.310 ;
        RECT 154.290 1763.065 158.050 1767.310 ;
        RECT 158.890 1763.065 162.190 1767.310 ;
        RECT 163.030 1763.065 166.790 1767.310 ;
        RECT 167.630 1763.065 171.390 1767.310 ;
        RECT 172.230 1763.065 175.530 1767.310 ;
        RECT 176.370 1763.065 180.130 1767.310 ;
        RECT 180.970 1763.065 184.730 1767.310 ;
        RECT 185.570 1763.065 189.330 1767.310 ;
        RECT 190.170 1763.065 193.470 1767.310 ;
        RECT 194.310 1763.065 198.070 1767.310 ;
        RECT 198.910 1763.065 202.670 1767.310 ;
        RECT 203.510 1763.065 207.270 1767.310 ;
        RECT 208.110 1763.065 211.410 1767.310 ;
        RECT 212.250 1763.065 216.010 1767.310 ;
        RECT 216.850 1763.065 220.610 1767.310 ;
        RECT 221.450 1763.065 224.750 1767.310 ;
        RECT 225.590 1763.065 229.350 1767.310 ;
        RECT 230.190 1763.065 233.950 1767.310 ;
        RECT 234.790 1763.065 238.550 1767.310 ;
        RECT 239.390 1763.065 242.690 1767.310 ;
        RECT 243.530 1763.065 247.290 1767.310 ;
        RECT 248.130 1763.065 251.890 1767.310 ;
        RECT 252.730 1763.065 256.030 1767.310 ;
        RECT 256.870 1763.065 260.630 1767.310 ;
        RECT 261.470 1763.065 265.230 1767.310 ;
        RECT 266.070 1763.065 269.830 1767.310 ;
        RECT 270.670 1763.065 273.970 1767.310 ;
        RECT 274.810 1763.065 278.570 1767.310 ;
        RECT 279.410 1763.065 283.170 1767.310 ;
        RECT 284.010 1763.065 287.310 1767.310 ;
        RECT 288.150 1763.065 291.910 1767.310 ;
        RECT 292.750 1763.065 296.510 1767.310 ;
        RECT 297.350 1763.065 301.110 1767.310 ;
        RECT 301.950 1763.065 305.250 1767.310 ;
        RECT 306.090 1763.065 309.850 1767.310 ;
        RECT 310.690 1763.065 314.450 1767.310 ;
        RECT 315.290 1763.065 318.590 1767.310 ;
        RECT 319.430 1763.065 323.190 1767.310 ;
        RECT 324.030 1763.065 327.790 1767.310 ;
        RECT 328.630 1763.065 332.390 1767.310 ;
        RECT 333.230 1763.065 336.530 1767.310 ;
        RECT 337.370 1763.065 341.130 1767.310 ;
        RECT 341.970 1763.065 345.730 1767.310 ;
        RECT 346.570 1763.065 349.870 1767.310 ;
        RECT 350.710 1763.065 354.470 1767.310 ;
        RECT 355.310 1763.065 359.070 1767.310 ;
        RECT 359.910 1763.065 363.670 1767.310 ;
        RECT 364.510 1763.065 367.810 1767.310 ;
        RECT 368.650 1763.065 372.410 1767.310 ;
        RECT 373.250 1763.065 377.010 1767.310 ;
        RECT 377.850 1763.065 381.150 1767.310 ;
        RECT 381.990 1763.065 385.750 1767.310 ;
        RECT 386.590 1763.065 390.350 1767.310 ;
        RECT 391.190 1763.065 394.950 1767.310 ;
        RECT 395.790 1763.065 399.090 1767.310 ;
        RECT 399.930 1763.065 403.690 1767.310 ;
        RECT 404.530 1763.065 408.290 1767.310 ;
        RECT 409.130 1763.065 412.890 1767.310 ;
        RECT 413.730 1763.065 417.030 1767.310 ;
        RECT 417.870 1763.065 421.630 1767.310 ;
        RECT 422.470 1763.065 426.230 1767.310 ;
        RECT 427.070 1763.065 430.370 1767.310 ;
        RECT 431.210 1763.065 434.970 1767.310 ;
        RECT 435.810 1763.065 439.570 1767.310 ;
        RECT 440.410 1763.065 444.170 1767.310 ;
        RECT 445.010 1763.065 448.310 1767.310 ;
        RECT 449.150 1763.065 452.910 1767.310 ;
        RECT 453.750 1763.065 457.510 1767.310 ;
        RECT 458.350 1763.065 461.650 1767.310 ;
        RECT 462.490 1763.065 466.250 1767.310 ;
        RECT 467.090 1763.065 470.850 1767.310 ;
        RECT 471.690 1763.065 475.450 1767.310 ;
        RECT 476.290 1763.065 479.590 1767.310 ;
        RECT 480.430 1763.065 484.190 1767.310 ;
        RECT 485.030 1763.065 488.790 1767.310 ;
        RECT 489.630 1763.065 492.930 1767.310 ;
        RECT 493.770 1763.065 497.530 1767.310 ;
        RECT 498.370 1763.065 502.130 1767.310 ;
        RECT 502.970 1763.065 506.730 1767.310 ;
        RECT 507.570 1763.065 510.870 1767.310 ;
        RECT 511.710 1763.065 515.470 1767.310 ;
        RECT 516.310 1763.065 520.070 1767.310 ;
        RECT 520.910 1763.065 524.210 1767.310 ;
        RECT 525.050 1763.065 528.810 1767.310 ;
        RECT 529.650 1763.065 533.410 1767.310 ;
        RECT 534.250 1763.065 538.010 1767.310 ;
        RECT 538.850 1763.065 542.150 1767.310 ;
        RECT 542.990 1763.065 546.750 1767.310 ;
        RECT 547.590 1763.065 551.350 1767.310 ;
        RECT 552.190 1763.065 555.490 1767.310 ;
        RECT 556.330 1763.065 560.090 1767.310 ;
        RECT 560.930 1763.065 564.690 1767.310 ;
        RECT 565.530 1763.065 569.290 1767.310 ;
        RECT 570.130 1763.065 573.430 1767.310 ;
        RECT 574.270 1763.065 578.030 1767.310 ;
        RECT 578.870 1763.065 582.630 1767.310 ;
        RECT 583.470 1763.065 587.230 1767.310 ;
        RECT 588.070 1763.065 591.370 1767.310 ;
        RECT 592.210 1763.065 595.970 1767.310 ;
        RECT 596.810 1763.065 600.570 1767.310 ;
        RECT 601.410 1763.065 604.710 1767.310 ;
        RECT 605.550 1763.065 609.310 1767.310 ;
        RECT 610.150 1763.065 613.910 1767.310 ;
        RECT 614.750 1763.065 618.510 1767.310 ;
        RECT 619.350 1763.065 622.650 1767.310 ;
        RECT 623.490 1763.065 627.250 1767.310 ;
        RECT 628.090 1763.065 631.850 1767.310 ;
        RECT 632.690 1763.065 635.990 1767.310 ;
        RECT 636.830 1763.065 640.590 1767.310 ;
        RECT 641.430 1763.065 645.190 1767.310 ;
        RECT 646.030 1763.065 649.790 1767.310 ;
        RECT 650.630 1763.065 653.930 1767.310 ;
        RECT 654.770 1763.065 658.530 1767.310 ;
        RECT 659.370 1763.065 663.130 1767.310 ;
        RECT 663.970 1763.065 667.270 1767.310 ;
        RECT 668.110 1763.065 671.870 1767.310 ;
        RECT 672.710 1763.065 676.470 1767.310 ;
        RECT 677.310 1763.065 681.070 1767.310 ;
        RECT 681.910 1763.065 685.210 1767.310 ;
        RECT 686.050 1763.065 689.810 1767.310 ;
        RECT 690.650 1763.065 694.410 1767.310 ;
        RECT 695.250 1763.065 698.550 1767.310 ;
        RECT 699.390 1763.065 703.150 1767.310 ;
        RECT 703.990 1763.065 707.750 1767.310 ;
        RECT 708.590 1763.065 712.350 1767.310 ;
        RECT 713.190 1763.065 716.490 1767.310 ;
        RECT 717.330 1763.065 721.090 1767.310 ;
        RECT 721.930 1763.065 725.690 1767.310 ;
        RECT 726.530 1763.065 729.830 1767.310 ;
        RECT 730.670 1763.065 734.430 1767.310 ;
        RECT 735.270 1763.065 739.030 1767.310 ;
        RECT 739.870 1763.065 743.630 1767.310 ;
        RECT 744.470 1763.065 747.770 1767.310 ;
        RECT 748.610 1763.065 752.370 1767.310 ;
        RECT 753.210 1763.065 756.970 1767.310 ;
        RECT 757.810 1763.065 761.110 1767.310 ;
        RECT 761.950 1763.065 765.710 1767.310 ;
        RECT 766.550 1763.065 770.310 1767.310 ;
        RECT 771.150 1763.065 774.910 1767.310 ;
        RECT 775.750 1763.065 779.050 1767.310 ;
        RECT 779.890 1763.065 783.650 1767.310 ;
        RECT 784.490 1763.065 788.250 1767.310 ;
        RECT 789.090 1763.065 792.850 1767.310 ;
        RECT 793.690 1763.065 796.990 1767.310 ;
        RECT 797.830 1763.065 801.590 1767.310 ;
        RECT 802.430 1763.065 806.190 1767.310 ;
        RECT 807.030 1763.065 810.330 1767.310 ;
        RECT 811.170 1763.065 814.930 1767.310 ;
        RECT 815.770 1763.065 819.530 1767.310 ;
        RECT 820.370 1763.065 824.130 1767.310 ;
        RECT 824.970 1763.065 828.270 1767.310 ;
        RECT 829.110 1763.065 832.870 1767.310 ;
        RECT 833.710 1763.065 837.470 1767.310 ;
        RECT 838.310 1763.065 841.610 1767.310 ;
        RECT 842.450 1763.065 846.210 1767.310 ;
        RECT 847.050 1763.065 850.810 1767.310 ;
        RECT 851.650 1763.065 855.410 1767.310 ;
        RECT 856.250 1763.065 859.550 1767.310 ;
        RECT 860.390 1763.065 864.150 1767.310 ;
        RECT 864.990 1763.065 868.750 1767.310 ;
        RECT 869.590 1763.065 872.890 1767.310 ;
        RECT 873.730 1763.065 877.490 1767.310 ;
        RECT 878.330 1763.065 882.090 1767.310 ;
        RECT 882.930 1763.065 886.690 1767.310 ;
        RECT 887.530 1763.065 890.830 1767.310 ;
        RECT 891.670 1763.065 895.430 1767.310 ;
        RECT 896.270 1763.065 900.030 1767.310 ;
        RECT 900.870 1763.065 904.170 1767.310 ;
        RECT 905.010 1763.065 908.770 1767.310 ;
        RECT 909.610 1763.065 913.370 1767.310 ;
        RECT 914.210 1763.065 917.970 1767.310 ;
        RECT 918.810 1763.065 922.110 1767.310 ;
        RECT 922.950 1763.065 926.710 1767.310 ;
        RECT 927.550 1763.065 931.310 1767.310 ;
        RECT 932.150 1763.065 935.450 1767.310 ;
        RECT 936.290 1763.065 940.050 1767.310 ;
        RECT 940.890 1763.065 944.650 1767.310 ;
        RECT 945.490 1763.065 949.250 1767.310 ;
        RECT 950.090 1763.065 953.390 1767.310 ;
        RECT 954.230 1763.065 957.990 1767.310 ;
        RECT 958.830 1763.065 962.590 1767.310 ;
        RECT 963.430 1763.065 966.730 1767.310 ;
        RECT 967.570 1763.065 971.330 1767.310 ;
        RECT 972.170 1763.065 975.930 1767.310 ;
        RECT 976.770 1763.065 980.530 1767.310 ;
        RECT 981.370 1763.065 984.670 1767.310 ;
        RECT 985.510 1763.065 989.270 1767.310 ;
        RECT 990.110 1763.065 993.870 1767.310 ;
        RECT 994.710 1763.065 998.470 1767.310 ;
        RECT 999.310 1763.065 1002.610 1767.310 ;
        RECT 1003.450 1763.065 1007.210 1767.310 ;
        RECT 1008.050 1763.065 1011.810 1767.310 ;
        RECT 1012.650 1763.065 1015.950 1767.310 ;
        RECT 1016.790 1763.065 1020.550 1767.310 ;
        RECT 1021.390 1763.065 1025.150 1767.310 ;
        RECT 1025.990 1763.065 1029.750 1767.310 ;
        RECT 1030.590 1763.065 1033.890 1767.310 ;
        RECT 1034.730 1763.065 1038.490 1767.310 ;
        RECT 1039.330 1763.065 1043.090 1767.310 ;
        RECT 1043.930 1763.065 1047.230 1767.310 ;
        RECT 1048.070 1763.065 1051.830 1767.310 ;
        RECT 1052.670 1763.065 1056.430 1767.310 ;
        RECT 1057.270 1763.065 1061.030 1767.310 ;
        RECT 1061.870 1763.065 1065.170 1767.310 ;
        RECT 1066.010 1763.065 1069.770 1767.310 ;
        RECT 1070.610 1763.065 1074.370 1767.310 ;
        RECT 1075.210 1763.065 1078.510 1767.310 ;
        RECT 1079.350 1763.065 1083.110 1767.310 ;
        RECT 1083.950 1763.065 1087.710 1767.310 ;
        RECT 1088.550 1763.065 1092.310 1767.310 ;
        RECT 1093.150 1763.065 1096.450 1767.310 ;
        RECT 1097.290 1763.065 1101.050 1767.310 ;
        RECT 1101.890 1763.065 1105.650 1767.310 ;
        RECT 1106.490 1763.065 1109.790 1767.310 ;
        RECT 1110.630 1763.065 1114.390 1767.310 ;
        RECT 1115.230 1763.065 1118.990 1767.310 ;
        RECT 1119.830 1763.065 1123.590 1767.310 ;
        RECT 1124.430 1763.065 1127.730 1767.310 ;
        RECT 1128.570 1763.065 1132.330 1767.310 ;
        RECT 1133.170 1763.065 1136.930 1767.310 ;
        RECT 1137.770 1763.065 1141.070 1767.310 ;
        RECT 1141.910 1763.065 1145.670 1767.310 ;
        RECT 1146.510 1763.065 1150.270 1767.310 ;
        RECT 1151.110 1763.065 1154.870 1767.310 ;
        RECT 1155.710 1763.065 1159.010 1767.310 ;
        RECT 1159.850 1763.065 1163.610 1767.310 ;
        RECT 1164.450 1763.065 1168.210 1767.310 ;
        RECT 1169.050 1763.065 1172.810 1767.310 ;
        RECT 1173.650 1763.065 1176.950 1767.310 ;
        RECT 1177.790 1763.065 1181.550 1767.310 ;
        RECT 1182.390 1763.065 1186.150 1767.310 ;
        RECT 1186.990 1763.065 1190.290 1767.310 ;
        RECT 1191.130 1763.065 1194.890 1767.310 ;
        RECT 1195.730 1763.065 1199.490 1767.310 ;
        RECT 1200.330 1763.065 1204.090 1767.310 ;
        RECT 1204.930 1763.065 1208.230 1767.310 ;
        RECT 1209.070 1763.065 1212.830 1767.310 ;
        RECT 1213.670 1763.065 1217.430 1767.310 ;
        RECT 1218.270 1763.065 1221.570 1767.310 ;
        RECT 1222.410 1763.065 1226.170 1767.310 ;
        RECT 1227.010 1763.065 1230.770 1767.310 ;
        RECT 1231.610 1763.065 1235.370 1767.310 ;
        RECT 1236.210 1763.065 1239.510 1767.310 ;
        RECT 1240.350 1763.065 1244.110 1767.310 ;
        RECT 1244.950 1763.065 1248.710 1767.310 ;
        RECT 1249.550 1763.065 1252.850 1767.310 ;
        RECT 1253.690 1763.065 1257.450 1767.310 ;
        RECT 1258.290 1763.065 1262.050 1767.310 ;
        RECT 1262.890 1763.065 1266.650 1767.310 ;
        RECT 1267.490 1763.065 1270.790 1767.310 ;
        RECT 1271.630 1763.065 1275.390 1767.310 ;
        RECT 1276.230 1763.065 1279.990 1767.310 ;
        RECT 1280.830 1763.065 1284.130 1767.310 ;
        RECT 1284.970 1763.065 1288.730 1767.310 ;
        RECT 1289.570 1763.065 1293.330 1767.310 ;
        RECT 1294.170 1763.065 1297.930 1767.310 ;
        RECT 1298.770 1763.065 1302.070 1767.310 ;
        RECT 1302.910 1763.065 1306.670 1767.310 ;
        RECT 1307.510 1763.065 1311.270 1767.310 ;
        RECT 1312.110 1763.065 1315.410 1767.310 ;
        RECT 1316.250 1763.065 1320.010 1767.310 ;
        RECT 1320.850 1763.065 1324.610 1767.310 ;
        RECT 1325.450 1763.065 1329.210 1767.310 ;
        RECT 1330.050 1763.065 1333.350 1767.310 ;
        RECT 1334.190 1763.065 1337.950 1767.310 ;
        RECT 1338.790 1763.065 1342.550 1767.310 ;
        RECT 1343.390 1763.065 1346.690 1767.310 ;
        RECT 1347.530 1763.065 1351.290 1767.310 ;
        RECT 1352.130 1763.065 1355.890 1767.310 ;
        RECT 1356.730 1763.065 1360.490 1767.310 ;
        RECT 1361.330 1763.065 1364.630 1767.310 ;
        RECT 1365.470 1763.065 1369.230 1767.310 ;
        RECT 1370.070 1763.065 1373.830 1767.310 ;
        RECT 1374.670 1763.065 1378.430 1767.310 ;
        RECT 1379.270 1763.065 1382.570 1767.310 ;
        RECT 1383.410 1763.065 1387.170 1767.310 ;
        RECT 1388.010 1763.065 1391.770 1767.310 ;
        RECT 1392.610 1763.065 1395.910 1767.310 ;
        RECT 1396.750 1763.065 1400.510 1767.310 ;
        RECT 1401.350 1763.065 1405.110 1767.310 ;
        RECT 1405.950 1763.065 1409.710 1767.310 ;
        RECT 1410.550 1763.065 1413.850 1767.310 ;
        RECT 1414.690 1763.065 1418.450 1767.310 ;
        RECT 1419.290 1763.065 1423.050 1767.310 ;
        RECT 1423.890 1763.065 1427.190 1767.310 ;
        RECT 1428.030 1763.065 1431.790 1767.310 ;
        RECT 1432.630 1763.065 1436.390 1767.310 ;
        RECT 1437.230 1763.065 1440.990 1767.310 ;
        RECT 1441.830 1763.065 1445.130 1767.310 ;
        RECT 1445.970 1763.065 1449.730 1767.310 ;
        RECT 1450.570 1763.065 1454.330 1767.310 ;
        RECT 1455.170 1763.065 1458.470 1767.310 ;
        RECT 1459.310 1763.065 1463.070 1767.310 ;
        RECT 1463.910 1763.065 1467.670 1767.310 ;
        RECT 1468.510 1763.065 1472.270 1767.310 ;
        RECT 1473.110 1763.065 1476.410 1767.310 ;
        RECT 1477.250 1763.065 1481.010 1767.310 ;
        RECT 1481.850 1763.065 1485.610 1767.310 ;
        RECT 1486.450 1763.065 1489.750 1767.310 ;
        RECT 1490.590 1763.065 1494.350 1767.310 ;
        RECT 1495.190 1763.065 1498.950 1767.310 ;
        RECT 1499.790 1763.065 1503.550 1767.310 ;
        RECT 1504.390 1763.065 1507.690 1767.310 ;
        RECT 1508.530 1763.065 1512.290 1767.310 ;
        RECT 1513.130 1763.065 1516.890 1767.310 ;
        RECT 1517.730 1763.065 1521.030 1767.310 ;
        RECT 1521.870 1763.065 1525.630 1767.310 ;
        RECT 1526.470 1763.065 1530.230 1767.310 ;
        RECT 1531.070 1763.065 1534.830 1767.310 ;
        RECT 1535.670 1763.065 1538.970 1767.310 ;
        RECT 1539.810 1763.065 1543.570 1767.310 ;
        RECT 1544.410 1763.065 1548.170 1767.310 ;
        RECT 1549.010 1763.065 1552.310 1767.310 ;
        RECT 1553.150 1763.065 1556.910 1767.310 ;
        RECT 1557.750 1763.065 1561.510 1767.310 ;
        RECT 1562.350 1763.065 1566.110 1767.310 ;
        RECT 1566.950 1763.065 1570.250 1767.310 ;
        RECT 1571.090 1763.065 1574.850 1767.310 ;
        RECT 1575.690 1763.065 1579.450 1767.310 ;
        RECT 1580.290 1763.065 1584.050 1767.310 ;
        RECT 1584.890 1763.065 1588.190 1767.310 ;
        RECT 1589.030 1763.065 1592.790 1767.310 ;
        RECT 1593.630 1763.065 1597.390 1767.310 ;
        RECT 1598.230 1763.065 1601.530 1767.310 ;
        RECT 1602.370 1763.065 1606.130 1767.310 ;
        RECT 1606.970 1763.065 1610.730 1767.310 ;
        RECT 1611.570 1763.065 1615.330 1767.310 ;
        RECT 1616.170 1763.065 1619.470 1767.310 ;
        RECT 1620.310 1763.065 1624.070 1767.310 ;
        RECT 1624.910 1763.065 1628.670 1767.310 ;
        RECT 1629.510 1763.065 1632.810 1767.310 ;
        RECT 1633.650 1763.065 1637.410 1767.310 ;
        RECT 1638.250 1763.065 1642.010 1767.310 ;
        RECT 1642.850 1763.065 1646.610 1767.310 ;
        RECT 1647.450 1763.065 1650.750 1767.310 ;
        RECT 1651.590 1763.065 1655.350 1767.310 ;
        RECT 1656.190 1763.065 1659.950 1767.310 ;
        RECT 1660.790 1763.065 1664.090 1767.310 ;
        RECT 1664.930 1763.065 1668.690 1767.310 ;
        RECT 1669.530 1763.065 1673.290 1767.310 ;
        RECT 1674.130 1763.065 1677.890 1767.310 ;
        RECT 1678.730 1763.065 1682.030 1767.310 ;
        RECT 1682.870 1763.065 1686.630 1767.310 ;
        RECT 1687.470 1763.065 1691.230 1767.310 ;
        RECT 1692.070 1763.065 1695.370 1767.310 ;
        RECT 1696.210 1763.065 1699.970 1767.310 ;
        RECT 1700.810 1763.065 1704.570 1767.310 ;
        RECT 1705.410 1763.065 1709.170 1767.310 ;
        RECT 1710.010 1763.065 1713.310 1767.310 ;
        RECT 1714.150 1763.065 1717.910 1767.310 ;
        RECT 1718.750 1763.065 1722.510 1767.310 ;
        RECT 1723.350 1763.065 1726.650 1767.310 ;
        RECT 1727.490 1763.065 1731.250 1767.310 ;
        RECT 1732.090 1763.065 1735.850 1767.310 ;
        RECT 1736.690 1763.065 1740.450 1767.310 ;
        RECT 1741.290 1763.065 1744.590 1767.310 ;
        RECT 1745.430 1763.065 1749.190 1767.310 ;
        RECT 1750.030 1763.065 1753.790 1767.310 ;
        RECT 1754.630 1763.065 1754.800 1767.310 ;
        RECT 1.480 4.280 1754.800 1763.065 ;
        RECT 2.030 3.670 4.410 4.280 ;
        RECT 5.250 3.670 8.090 4.280 ;
        RECT 8.930 3.670 11.770 4.280 ;
        RECT 12.610 3.670 14.990 4.280 ;
        RECT 15.830 3.670 18.670 4.280 ;
        RECT 19.510 3.670 22.350 4.280 ;
        RECT 23.190 3.670 26.030 4.280 ;
        RECT 26.870 3.670 29.250 4.280 ;
        RECT 30.090 3.670 32.930 4.280 ;
        RECT 33.770 3.670 36.610 4.280 ;
        RECT 37.450 3.670 40.290 4.280 ;
        RECT 41.130 3.670 43.510 4.280 ;
        RECT 44.350 3.670 47.190 4.280 ;
        RECT 48.030 3.670 50.870 4.280 ;
        RECT 51.710 3.670 54.550 4.280 ;
        RECT 55.390 3.670 57.770 4.280 ;
        RECT 58.610 3.670 61.450 4.280 ;
        RECT 62.290 3.670 65.130 4.280 ;
        RECT 65.970 3.670 68.810 4.280 ;
        RECT 69.650 3.670 72.030 4.280 ;
        RECT 72.870 3.670 75.710 4.280 ;
        RECT 76.550 3.670 79.390 4.280 ;
        RECT 80.230 3.670 83.070 4.280 ;
        RECT 83.910 3.670 86.290 4.280 ;
        RECT 87.130 3.670 89.970 4.280 ;
        RECT 90.810 3.670 93.650 4.280 ;
        RECT 94.490 3.670 97.330 4.280 ;
        RECT 98.170 3.670 100.550 4.280 ;
        RECT 101.390 3.670 104.230 4.280 ;
        RECT 105.070 3.670 107.910 4.280 ;
        RECT 108.750 3.670 111.590 4.280 ;
        RECT 112.430 3.670 114.810 4.280 ;
        RECT 115.650 3.670 118.490 4.280 ;
        RECT 119.330 3.670 122.170 4.280 ;
        RECT 123.010 3.670 125.850 4.280 ;
        RECT 126.690 3.670 129.070 4.280 ;
        RECT 129.910 3.670 132.750 4.280 ;
        RECT 133.590 3.670 136.430 4.280 ;
        RECT 137.270 3.670 140.110 4.280 ;
        RECT 140.950 3.670 143.330 4.280 ;
        RECT 144.170 3.670 147.010 4.280 ;
        RECT 147.850 3.670 150.690 4.280 ;
        RECT 151.530 3.670 154.370 4.280 ;
        RECT 155.210 3.670 157.590 4.280 ;
        RECT 158.430 3.670 161.270 4.280 ;
        RECT 162.110 3.670 164.950 4.280 ;
        RECT 165.790 3.670 168.630 4.280 ;
        RECT 169.470 3.670 171.850 4.280 ;
        RECT 172.690 3.670 175.530 4.280 ;
        RECT 176.370 3.670 179.210 4.280 ;
        RECT 180.050 3.670 182.890 4.280 ;
        RECT 183.730 3.670 186.110 4.280 ;
        RECT 186.950 3.670 189.790 4.280 ;
        RECT 190.630 3.670 193.470 4.280 ;
        RECT 194.310 3.670 197.150 4.280 ;
        RECT 197.990 3.670 200.370 4.280 ;
        RECT 201.210 3.670 204.050 4.280 ;
        RECT 204.890 3.670 207.730 4.280 ;
        RECT 208.570 3.670 211.410 4.280 ;
        RECT 212.250 3.670 214.630 4.280 ;
        RECT 215.470 3.670 218.310 4.280 ;
        RECT 219.150 3.670 221.990 4.280 ;
        RECT 222.830 3.670 225.670 4.280 ;
        RECT 226.510 3.670 228.890 4.280 ;
        RECT 229.730 3.670 232.570 4.280 ;
        RECT 233.410 3.670 236.250 4.280 ;
        RECT 237.090 3.670 239.930 4.280 ;
        RECT 240.770 3.670 243.150 4.280 ;
        RECT 243.990 3.670 246.830 4.280 ;
        RECT 247.670 3.670 250.510 4.280 ;
        RECT 251.350 3.670 253.730 4.280 ;
        RECT 254.570 3.670 257.410 4.280 ;
        RECT 258.250 3.670 261.090 4.280 ;
        RECT 261.930 3.670 264.770 4.280 ;
        RECT 265.610 3.670 267.990 4.280 ;
        RECT 268.830 3.670 271.670 4.280 ;
        RECT 272.510 3.670 275.350 4.280 ;
        RECT 276.190 3.670 279.030 4.280 ;
        RECT 279.870 3.670 282.250 4.280 ;
        RECT 283.090 3.670 285.930 4.280 ;
        RECT 286.770 3.670 289.610 4.280 ;
        RECT 290.450 3.670 293.290 4.280 ;
        RECT 294.130 3.670 296.510 4.280 ;
        RECT 297.350 3.670 300.190 4.280 ;
        RECT 301.030 3.670 303.870 4.280 ;
        RECT 304.710 3.670 307.550 4.280 ;
        RECT 308.390 3.670 310.770 4.280 ;
        RECT 311.610 3.670 314.450 4.280 ;
        RECT 315.290 3.670 318.130 4.280 ;
        RECT 318.970 3.670 321.810 4.280 ;
        RECT 322.650 3.670 325.030 4.280 ;
        RECT 325.870 3.670 328.710 4.280 ;
        RECT 329.550 3.670 332.390 4.280 ;
        RECT 333.230 3.670 336.070 4.280 ;
        RECT 336.910 3.670 339.290 4.280 ;
        RECT 340.130 3.670 342.970 4.280 ;
        RECT 343.810 3.670 346.650 4.280 ;
        RECT 347.490 3.670 350.330 4.280 ;
        RECT 351.170 3.670 353.550 4.280 ;
        RECT 354.390 3.670 357.230 4.280 ;
        RECT 358.070 3.670 360.910 4.280 ;
        RECT 361.750 3.670 364.590 4.280 ;
        RECT 365.430 3.670 367.810 4.280 ;
        RECT 368.650 3.670 371.490 4.280 ;
        RECT 372.330 3.670 375.170 4.280 ;
        RECT 376.010 3.670 378.850 4.280 ;
        RECT 379.690 3.670 382.070 4.280 ;
        RECT 382.910 3.670 385.750 4.280 ;
        RECT 386.590 3.670 389.430 4.280 ;
        RECT 390.270 3.670 393.110 4.280 ;
        RECT 393.950 3.670 396.330 4.280 ;
        RECT 397.170 3.670 400.010 4.280 ;
        RECT 400.850 3.670 403.690 4.280 ;
        RECT 404.530 3.670 407.370 4.280 ;
        RECT 408.210 3.670 410.590 4.280 ;
        RECT 411.430 3.670 414.270 4.280 ;
        RECT 415.110 3.670 417.950 4.280 ;
        RECT 418.790 3.670 421.630 4.280 ;
        RECT 422.470 3.670 424.850 4.280 ;
        RECT 425.690 3.670 428.530 4.280 ;
        RECT 429.370 3.670 432.210 4.280 ;
        RECT 433.050 3.670 435.890 4.280 ;
        RECT 436.730 3.670 439.110 4.280 ;
        RECT 439.950 3.670 442.790 4.280 ;
        RECT 443.630 3.670 446.470 4.280 ;
        RECT 447.310 3.670 450.150 4.280 ;
        RECT 450.990 3.670 453.370 4.280 ;
        RECT 454.210 3.670 457.050 4.280 ;
        RECT 457.890 3.670 460.730 4.280 ;
        RECT 461.570 3.670 464.410 4.280 ;
        RECT 465.250 3.670 467.630 4.280 ;
        RECT 468.470 3.670 471.310 4.280 ;
        RECT 472.150 3.670 474.990 4.280 ;
        RECT 475.830 3.670 478.670 4.280 ;
        RECT 479.510 3.670 481.890 4.280 ;
        RECT 482.730 3.670 485.570 4.280 ;
        RECT 486.410 3.670 489.250 4.280 ;
        RECT 490.090 3.670 492.930 4.280 ;
        RECT 493.770 3.670 496.150 4.280 ;
        RECT 496.990 3.670 499.830 4.280 ;
        RECT 500.670 3.670 503.510 4.280 ;
        RECT 504.350 3.670 506.730 4.280 ;
        RECT 507.570 3.670 510.410 4.280 ;
        RECT 511.250 3.670 514.090 4.280 ;
        RECT 514.930 3.670 517.770 4.280 ;
        RECT 518.610 3.670 520.990 4.280 ;
        RECT 521.830 3.670 524.670 4.280 ;
        RECT 525.510 3.670 528.350 4.280 ;
        RECT 529.190 3.670 532.030 4.280 ;
        RECT 532.870 3.670 535.250 4.280 ;
        RECT 536.090 3.670 538.930 4.280 ;
        RECT 539.770 3.670 542.610 4.280 ;
        RECT 543.450 3.670 546.290 4.280 ;
        RECT 547.130 3.670 549.510 4.280 ;
        RECT 550.350 3.670 553.190 4.280 ;
        RECT 554.030 3.670 556.870 4.280 ;
        RECT 557.710 3.670 560.550 4.280 ;
        RECT 561.390 3.670 563.770 4.280 ;
        RECT 564.610 3.670 567.450 4.280 ;
        RECT 568.290 3.670 571.130 4.280 ;
        RECT 571.970 3.670 574.810 4.280 ;
        RECT 575.650 3.670 578.030 4.280 ;
        RECT 578.870 3.670 581.710 4.280 ;
        RECT 582.550 3.670 585.390 4.280 ;
        RECT 586.230 3.670 589.070 4.280 ;
        RECT 589.910 3.670 592.290 4.280 ;
        RECT 593.130 3.670 595.970 4.280 ;
        RECT 596.810 3.670 599.650 4.280 ;
        RECT 600.490 3.670 603.330 4.280 ;
        RECT 604.170 3.670 606.550 4.280 ;
        RECT 607.390 3.670 610.230 4.280 ;
        RECT 611.070 3.670 613.910 4.280 ;
        RECT 614.750 3.670 617.590 4.280 ;
        RECT 618.430 3.670 620.810 4.280 ;
        RECT 621.650 3.670 624.490 4.280 ;
        RECT 625.330 3.670 628.170 4.280 ;
        RECT 629.010 3.670 631.850 4.280 ;
        RECT 632.690 3.670 635.070 4.280 ;
        RECT 635.910 3.670 638.750 4.280 ;
        RECT 639.590 3.670 642.430 4.280 ;
        RECT 643.270 3.670 646.110 4.280 ;
        RECT 646.950 3.670 649.330 4.280 ;
        RECT 650.170 3.670 653.010 4.280 ;
        RECT 653.850 3.670 656.690 4.280 ;
        RECT 657.530 3.670 660.370 4.280 ;
        RECT 661.210 3.670 663.590 4.280 ;
        RECT 664.430 3.670 667.270 4.280 ;
        RECT 668.110 3.670 670.950 4.280 ;
        RECT 671.790 3.670 674.630 4.280 ;
        RECT 675.470 3.670 677.850 4.280 ;
        RECT 678.690 3.670 681.530 4.280 ;
        RECT 682.370 3.670 685.210 4.280 ;
        RECT 686.050 3.670 688.890 4.280 ;
        RECT 689.730 3.670 692.110 4.280 ;
        RECT 692.950 3.670 695.790 4.280 ;
        RECT 696.630 3.670 699.470 4.280 ;
        RECT 700.310 3.670 703.150 4.280 ;
        RECT 703.990 3.670 706.370 4.280 ;
        RECT 707.210 3.670 710.050 4.280 ;
        RECT 710.890 3.670 713.730 4.280 ;
        RECT 714.570 3.670 717.410 4.280 ;
        RECT 718.250 3.670 720.630 4.280 ;
        RECT 721.470 3.670 724.310 4.280 ;
        RECT 725.150 3.670 727.990 4.280 ;
        RECT 728.830 3.670 731.670 4.280 ;
        RECT 732.510 3.670 734.890 4.280 ;
        RECT 735.730 3.670 738.570 4.280 ;
        RECT 739.410 3.670 742.250 4.280 ;
        RECT 743.090 3.670 745.930 4.280 ;
        RECT 746.770 3.670 749.150 4.280 ;
        RECT 749.990 3.670 752.830 4.280 ;
        RECT 753.670 3.670 756.510 4.280 ;
        RECT 757.350 3.670 759.730 4.280 ;
        RECT 760.570 3.670 763.410 4.280 ;
        RECT 764.250 3.670 767.090 4.280 ;
        RECT 767.930 3.670 770.770 4.280 ;
        RECT 771.610 3.670 773.990 4.280 ;
        RECT 774.830 3.670 777.670 4.280 ;
        RECT 778.510 3.670 781.350 4.280 ;
        RECT 782.190 3.670 785.030 4.280 ;
        RECT 785.870 3.670 788.250 4.280 ;
        RECT 789.090 3.670 791.930 4.280 ;
        RECT 792.770 3.670 795.610 4.280 ;
        RECT 796.450 3.670 799.290 4.280 ;
        RECT 800.130 3.670 802.510 4.280 ;
        RECT 803.350 3.670 806.190 4.280 ;
        RECT 807.030 3.670 809.870 4.280 ;
        RECT 810.710 3.670 813.550 4.280 ;
        RECT 814.390 3.670 816.770 4.280 ;
        RECT 817.610 3.670 820.450 4.280 ;
        RECT 821.290 3.670 824.130 4.280 ;
        RECT 824.970 3.670 827.810 4.280 ;
        RECT 828.650 3.670 831.030 4.280 ;
        RECT 831.870 3.670 834.710 4.280 ;
        RECT 835.550 3.670 838.390 4.280 ;
        RECT 839.230 3.670 842.070 4.280 ;
        RECT 842.910 3.670 845.290 4.280 ;
        RECT 846.130 3.670 848.970 4.280 ;
        RECT 849.810 3.670 852.650 4.280 ;
        RECT 853.490 3.670 856.330 4.280 ;
        RECT 857.170 3.670 859.550 4.280 ;
        RECT 860.390 3.670 863.230 4.280 ;
        RECT 864.070 3.670 866.910 4.280 ;
        RECT 867.750 3.670 870.590 4.280 ;
        RECT 871.430 3.670 873.810 4.280 ;
        RECT 874.650 3.670 877.490 4.280 ;
        RECT 878.330 3.670 881.170 4.280 ;
        RECT 882.010 3.670 884.850 4.280 ;
        RECT 885.690 3.670 888.070 4.280 ;
        RECT 888.910 3.670 891.750 4.280 ;
        RECT 892.590 3.670 895.430 4.280 ;
        RECT 896.270 3.670 899.110 4.280 ;
        RECT 899.950 3.670 902.330 4.280 ;
        RECT 903.170 3.670 906.010 4.280 ;
        RECT 906.850 3.670 909.690 4.280 ;
        RECT 910.530 3.670 913.370 4.280 ;
        RECT 914.210 3.670 916.590 4.280 ;
        RECT 917.430 3.670 920.270 4.280 ;
        RECT 921.110 3.670 923.950 4.280 ;
        RECT 924.790 3.670 927.630 4.280 ;
        RECT 928.470 3.670 930.850 4.280 ;
        RECT 931.690 3.670 934.530 4.280 ;
        RECT 935.370 3.670 938.210 4.280 ;
        RECT 939.050 3.670 941.890 4.280 ;
        RECT 942.730 3.670 945.110 4.280 ;
        RECT 945.950 3.670 948.790 4.280 ;
        RECT 949.630 3.670 952.470 4.280 ;
        RECT 953.310 3.670 956.150 4.280 ;
        RECT 956.990 3.670 959.370 4.280 ;
        RECT 960.210 3.670 963.050 4.280 ;
        RECT 963.890 3.670 966.730 4.280 ;
        RECT 967.570 3.670 970.410 4.280 ;
        RECT 971.250 3.670 973.630 4.280 ;
        RECT 974.470 3.670 977.310 4.280 ;
        RECT 978.150 3.670 980.990 4.280 ;
        RECT 981.830 3.670 984.670 4.280 ;
        RECT 985.510 3.670 987.890 4.280 ;
        RECT 988.730 3.670 991.570 4.280 ;
        RECT 992.410 3.670 995.250 4.280 ;
        RECT 996.090 3.670 998.930 4.280 ;
        RECT 999.770 3.670 1002.150 4.280 ;
        RECT 1002.990 3.670 1005.830 4.280 ;
        RECT 1006.670 3.670 1009.510 4.280 ;
        RECT 1010.350 3.670 1012.730 4.280 ;
        RECT 1013.570 3.670 1016.410 4.280 ;
        RECT 1017.250 3.670 1020.090 4.280 ;
        RECT 1020.930 3.670 1023.770 4.280 ;
        RECT 1024.610 3.670 1026.990 4.280 ;
        RECT 1027.830 3.670 1030.670 4.280 ;
        RECT 1031.510 3.670 1034.350 4.280 ;
        RECT 1035.190 3.670 1038.030 4.280 ;
        RECT 1038.870 3.670 1041.250 4.280 ;
        RECT 1042.090 3.670 1044.930 4.280 ;
        RECT 1045.770 3.670 1048.610 4.280 ;
        RECT 1049.450 3.670 1052.290 4.280 ;
        RECT 1053.130 3.670 1055.510 4.280 ;
        RECT 1056.350 3.670 1059.190 4.280 ;
        RECT 1060.030 3.670 1062.870 4.280 ;
        RECT 1063.710 3.670 1066.550 4.280 ;
        RECT 1067.390 3.670 1069.770 4.280 ;
        RECT 1070.610 3.670 1073.450 4.280 ;
        RECT 1074.290 3.670 1077.130 4.280 ;
        RECT 1077.970 3.670 1080.810 4.280 ;
        RECT 1081.650 3.670 1084.030 4.280 ;
        RECT 1084.870 3.670 1087.710 4.280 ;
        RECT 1088.550 3.670 1091.390 4.280 ;
        RECT 1092.230 3.670 1095.070 4.280 ;
        RECT 1095.910 3.670 1098.290 4.280 ;
        RECT 1099.130 3.670 1101.970 4.280 ;
        RECT 1102.810 3.670 1105.650 4.280 ;
        RECT 1106.490 3.670 1109.330 4.280 ;
        RECT 1110.170 3.670 1112.550 4.280 ;
        RECT 1113.390 3.670 1116.230 4.280 ;
        RECT 1117.070 3.670 1119.910 4.280 ;
        RECT 1120.750 3.670 1123.590 4.280 ;
        RECT 1124.430 3.670 1126.810 4.280 ;
        RECT 1127.650 3.670 1130.490 4.280 ;
        RECT 1131.330 3.670 1134.170 4.280 ;
        RECT 1135.010 3.670 1137.850 4.280 ;
        RECT 1138.690 3.670 1141.070 4.280 ;
        RECT 1141.910 3.670 1144.750 4.280 ;
        RECT 1145.590 3.670 1148.430 4.280 ;
        RECT 1149.270 3.670 1152.110 4.280 ;
        RECT 1152.950 3.670 1155.330 4.280 ;
        RECT 1156.170 3.670 1159.010 4.280 ;
        RECT 1159.850 3.670 1162.690 4.280 ;
        RECT 1163.530 3.670 1166.370 4.280 ;
        RECT 1167.210 3.670 1169.590 4.280 ;
        RECT 1170.430 3.670 1173.270 4.280 ;
        RECT 1174.110 3.670 1176.950 4.280 ;
        RECT 1177.790 3.670 1180.630 4.280 ;
        RECT 1181.470 3.670 1183.850 4.280 ;
        RECT 1184.690 3.670 1187.530 4.280 ;
        RECT 1188.370 3.670 1191.210 4.280 ;
        RECT 1192.050 3.670 1194.890 4.280 ;
        RECT 1195.730 3.670 1198.110 4.280 ;
        RECT 1198.950 3.670 1201.790 4.280 ;
        RECT 1202.630 3.670 1205.470 4.280 ;
        RECT 1206.310 3.670 1209.150 4.280 ;
        RECT 1209.990 3.670 1212.370 4.280 ;
        RECT 1213.210 3.670 1216.050 4.280 ;
        RECT 1216.890 3.670 1219.730 4.280 ;
        RECT 1220.570 3.670 1223.410 4.280 ;
        RECT 1224.250 3.670 1226.630 4.280 ;
        RECT 1227.470 3.670 1230.310 4.280 ;
        RECT 1231.150 3.670 1233.990 4.280 ;
        RECT 1234.830 3.670 1237.670 4.280 ;
        RECT 1238.510 3.670 1240.890 4.280 ;
        RECT 1241.730 3.670 1244.570 4.280 ;
        RECT 1245.410 3.670 1248.250 4.280 ;
        RECT 1249.090 3.670 1251.930 4.280 ;
        RECT 1252.770 3.670 1255.150 4.280 ;
        RECT 1255.990 3.670 1258.830 4.280 ;
        RECT 1259.670 3.670 1262.510 4.280 ;
        RECT 1263.350 3.670 1265.730 4.280 ;
        RECT 1266.570 3.670 1269.410 4.280 ;
        RECT 1270.250 3.670 1273.090 4.280 ;
        RECT 1273.930 3.670 1276.770 4.280 ;
        RECT 1277.610 3.670 1279.990 4.280 ;
        RECT 1280.830 3.670 1283.670 4.280 ;
        RECT 1284.510 3.670 1287.350 4.280 ;
        RECT 1288.190 3.670 1291.030 4.280 ;
        RECT 1291.870 3.670 1294.250 4.280 ;
        RECT 1295.090 3.670 1297.930 4.280 ;
        RECT 1298.770 3.670 1301.610 4.280 ;
        RECT 1302.450 3.670 1305.290 4.280 ;
        RECT 1306.130 3.670 1308.510 4.280 ;
        RECT 1309.350 3.670 1312.190 4.280 ;
        RECT 1313.030 3.670 1315.870 4.280 ;
        RECT 1316.710 3.670 1319.550 4.280 ;
        RECT 1320.390 3.670 1322.770 4.280 ;
        RECT 1323.610 3.670 1326.450 4.280 ;
        RECT 1327.290 3.670 1330.130 4.280 ;
        RECT 1330.970 3.670 1333.810 4.280 ;
        RECT 1334.650 3.670 1337.030 4.280 ;
        RECT 1337.870 3.670 1340.710 4.280 ;
        RECT 1341.550 3.670 1344.390 4.280 ;
        RECT 1345.230 3.670 1348.070 4.280 ;
        RECT 1348.910 3.670 1351.290 4.280 ;
        RECT 1352.130 3.670 1354.970 4.280 ;
        RECT 1355.810 3.670 1358.650 4.280 ;
        RECT 1359.490 3.670 1362.330 4.280 ;
        RECT 1363.170 3.670 1365.550 4.280 ;
        RECT 1366.390 3.670 1369.230 4.280 ;
        RECT 1370.070 3.670 1372.910 4.280 ;
        RECT 1373.750 3.670 1376.590 4.280 ;
        RECT 1377.430 3.670 1379.810 4.280 ;
        RECT 1380.650 3.670 1383.490 4.280 ;
        RECT 1384.330 3.670 1387.170 4.280 ;
        RECT 1388.010 3.670 1390.850 4.280 ;
        RECT 1391.690 3.670 1394.070 4.280 ;
        RECT 1394.910 3.670 1397.750 4.280 ;
        RECT 1398.590 3.670 1401.430 4.280 ;
        RECT 1402.270 3.670 1405.110 4.280 ;
        RECT 1405.950 3.670 1408.330 4.280 ;
        RECT 1409.170 3.670 1412.010 4.280 ;
        RECT 1412.850 3.670 1415.690 4.280 ;
        RECT 1416.530 3.670 1419.370 4.280 ;
        RECT 1420.210 3.670 1422.590 4.280 ;
        RECT 1423.430 3.670 1426.270 4.280 ;
        RECT 1427.110 3.670 1429.950 4.280 ;
        RECT 1430.790 3.670 1433.630 4.280 ;
        RECT 1434.470 3.670 1436.850 4.280 ;
        RECT 1437.690 3.670 1440.530 4.280 ;
        RECT 1441.370 3.670 1444.210 4.280 ;
        RECT 1445.050 3.670 1447.890 4.280 ;
        RECT 1448.730 3.670 1451.110 4.280 ;
        RECT 1451.950 3.670 1454.790 4.280 ;
        RECT 1455.630 3.670 1458.470 4.280 ;
        RECT 1459.310 3.670 1462.150 4.280 ;
        RECT 1462.990 3.670 1465.370 4.280 ;
        RECT 1466.210 3.670 1469.050 4.280 ;
        RECT 1469.890 3.670 1472.730 4.280 ;
        RECT 1473.570 3.670 1476.410 4.280 ;
        RECT 1477.250 3.670 1479.630 4.280 ;
        RECT 1480.470 3.670 1483.310 4.280 ;
        RECT 1484.150 3.670 1486.990 4.280 ;
        RECT 1487.830 3.670 1490.670 4.280 ;
        RECT 1491.510 3.670 1493.890 4.280 ;
        RECT 1494.730 3.670 1497.570 4.280 ;
        RECT 1498.410 3.670 1501.250 4.280 ;
        RECT 1502.090 3.670 1504.930 4.280 ;
        RECT 1505.770 3.670 1508.150 4.280 ;
        RECT 1508.990 3.670 1511.830 4.280 ;
        RECT 1512.670 3.670 1515.510 4.280 ;
        RECT 1516.350 3.670 1518.730 4.280 ;
        RECT 1519.570 3.670 1522.410 4.280 ;
        RECT 1523.250 3.670 1526.090 4.280 ;
        RECT 1526.930 3.670 1529.770 4.280 ;
        RECT 1530.610 3.670 1532.990 4.280 ;
        RECT 1533.830 3.670 1536.670 4.280 ;
        RECT 1537.510 3.670 1540.350 4.280 ;
        RECT 1541.190 3.670 1544.030 4.280 ;
        RECT 1544.870 3.670 1547.250 4.280 ;
        RECT 1548.090 3.670 1550.930 4.280 ;
        RECT 1551.770 3.670 1554.610 4.280 ;
        RECT 1555.450 3.670 1558.290 4.280 ;
        RECT 1559.130 3.670 1561.510 4.280 ;
        RECT 1562.350 3.670 1565.190 4.280 ;
        RECT 1566.030 3.670 1568.870 4.280 ;
        RECT 1569.710 3.670 1572.550 4.280 ;
        RECT 1573.390 3.670 1575.770 4.280 ;
        RECT 1576.610 3.670 1579.450 4.280 ;
        RECT 1580.290 3.670 1583.130 4.280 ;
        RECT 1583.970 3.670 1586.810 4.280 ;
        RECT 1587.650 3.670 1590.030 4.280 ;
        RECT 1590.870 3.670 1593.710 4.280 ;
        RECT 1594.550 3.670 1597.390 4.280 ;
        RECT 1598.230 3.670 1601.070 4.280 ;
        RECT 1601.910 3.670 1604.290 4.280 ;
        RECT 1605.130 3.670 1607.970 4.280 ;
        RECT 1608.810 3.670 1611.650 4.280 ;
        RECT 1612.490 3.670 1615.330 4.280 ;
        RECT 1616.170 3.670 1618.550 4.280 ;
        RECT 1619.390 3.670 1622.230 4.280 ;
        RECT 1623.070 3.670 1625.910 4.280 ;
        RECT 1626.750 3.670 1629.590 4.280 ;
        RECT 1630.430 3.670 1632.810 4.280 ;
        RECT 1633.650 3.670 1636.490 4.280 ;
        RECT 1637.330 3.670 1640.170 4.280 ;
        RECT 1641.010 3.670 1643.850 4.280 ;
        RECT 1644.690 3.670 1647.070 4.280 ;
        RECT 1647.910 3.670 1650.750 4.280 ;
        RECT 1651.590 3.670 1654.430 4.280 ;
        RECT 1655.270 3.670 1658.110 4.280 ;
        RECT 1658.950 3.670 1661.330 4.280 ;
        RECT 1662.170 3.670 1665.010 4.280 ;
        RECT 1665.850 3.670 1668.690 4.280 ;
        RECT 1669.530 3.670 1672.370 4.280 ;
        RECT 1673.210 3.670 1675.590 4.280 ;
        RECT 1676.430 3.670 1679.270 4.280 ;
        RECT 1680.110 3.670 1682.950 4.280 ;
        RECT 1683.790 3.670 1686.630 4.280 ;
        RECT 1687.470 3.670 1689.850 4.280 ;
        RECT 1690.690 3.670 1693.530 4.280 ;
        RECT 1694.370 3.670 1697.210 4.280 ;
        RECT 1698.050 3.670 1700.890 4.280 ;
        RECT 1701.730 3.670 1704.110 4.280 ;
        RECT 1704.950 3.670 1707.790 4.280 ;
        RECT 1708.630 3.670 1711.470 4.280 ;
        RECT 1712.310 3.670 1715.150 4.280 ;
        RECT 1715.990 3.670 1718.370 4.280 ;
        RECT 1719.210 3.670 1722.050 4.280 ;
        RECT 1722.890 3.670 1725.730 4.280 ;
        RECT 1726.570 3.670 1729.410 4.280 ;
        RECT 1730.250 3.670 1732.630 4.280 ;
        RECT 1733.470 3.670 1736.310 4.280 ;
        RECT 1737.150 3.670 1739.990 4.280 ;
        RECT 1740.830 3.670 1743.670 4.280 ;
        RECT 1744.510 3.670 1746.890 4.280 ;
        RECT 1747.730 3.670 1750.570 4.280 ;
        RECT 1751.410 3.670 1754.250 4.280 ;
      LAYER met3 ;
        RECT 1.905 1763.600 1741.495 1767.145 ;
        RECT 4.400 1762.200 1741.495 1763.600 ;
        RECT 1.905 1756.120 1741.495 1762.200 ;
        RECT 4.400 1754.720 1741.495 1756.120 ;
        RECT 1.905 1747.960 1741.495 1754.720 ;
        RECT 4.400 1746.560 1741.495 1747.960 ;
        RECT 1.905 1740.480 1741.495 1746.560 ;
        RECT 4.400 1739.080 1741.495 1740.480 ;
        RECT 1.905 1732.320 1741.495 1739.080 ;
        RECT 4.400 1730.920 1741.495 1732.320 ;
        RECT 1.905 1724.840 1741.495 1730.920 ;
        RECT 4.400 1723.440 1741.495 1724.840 ;
        RECT 1.905 1716.680 1741.495 1723.440 ;
        RECT 4.400 1715.280 1741.495 1716.680 ;
        RECT 1.905 1709.200 1741.495 1715.280 ;
        RECT 4.400 1707.800 1741.495 1709.200 ;
        RECT 1.905 1701.040 1741.495 1707.800 ;
        RECT 4.400 1699.640 1741.495 1701.040 ;
        RECT 1.905 1693.560 1741.495 1699.640 ;
        RECT 4.400 1692.160 1741.495 1693.560 ;
        RECT 1.905 1685.400 1741.495 1692.160 ;
        RECT 4.400 1684.000 1741.495 1685.400 ;
        RECT 1.905 1677.920 1741.495 1684.000 ;
        RECT 4.400 1676.520 1741.495 1677.920 ;
        RECT 1.905 1669.760 1741.495 1676.520 ;
        RECT 4.400 1668.360 1741.495 1669.760 ;
        RECT 1.905 1662.280 1741.495 1668.360 ;
        RECT 4.400 1660.880 1741.495 1662.280 ;
        RECT 1.905 1654.120 1741.495 1660.880 ;
        RECT 4.400 1652.720 1741.495 1654.120 ;
        RECT 1.905 1646.640 1741.495 1652.720 ;
        RECT 4.400 1645.240 1741.495 1646.640 ;
        RECT 1.905 1638.480 1741.495 1645.240 ;
        RECT 4.400 1637.080 1741.495 1638.480 ;
        RECT 1.905 1631.000 1741.495 1637.080 ;
        RECT 4.400 1629.600 1741.495 1631.000 ;
        RECT 1.905 1622.840 1741.495 1629.600 ;
        RECT 4.400 1621.440 1741.495 1622.840 ;
        RECT 1.905 1615.360 1741.495 1621.440 ;
        RECT 4.400 1613.960 1741.495 1615.360 ;
        RECT 1.905 1607.200 1741.495 1613.960 ;
        RECT 4.400 1605.800 1741.495 1607.200 ;
        RECT 1.905 1599.720 1741.495 1605.800 ;
        RECT 4.400 1598.320 1741.495 1599.720 ;
        RECT 1.905 1591.560 1741.495 1598.320 ;
        RECT 4.400 1590.160 1741.495 1591.560 ;
        RECT 1.905 1584.080 1741.495 1590.160 ;
        RECT 4.400 1582.680 1741.495 1584.080 ;
        RECT 1.905 1575.920 1741.495 1582.680 ;
        RECT 4.400 1574.520 1741.495 1575.920 ;
        RECT 1.905 1568.440 1741.495 1574.520 ;
        RECT 4.400 1567.040 1741.495 1568.440 ;
        RECT 1.905 1560.280 1741.495 1567.040 ;
        RECT 4.400 1558.880 1741.495 1560.280 ;
        RECT 1.905 1552.800 1741.495 1558.880 ;
        RECT 4.400 1551.400 1741.495 1552.800 ;
        RECT 1.905 1544.640 1741.495 1551.400 ;
        RECT 4.400 1543.240 1741.495 1544.640 ;
        RECT 1.905 1537.160 1741.495 1543.240 ;
        RECT 4.400 1535.760 1741.495 1537.160 ;
        RECT 1.905 1529.000 1741.495 1535.760 ;
        RECT 4.400 1527.600 1741.495 1529.000 ;
        RECT 1.905 1521.520 1741.495 1527.600 ;
        RECT 4.400 1520.120 1741.495 1521.520 ;
        RECT 1.905 1513.360 1741.495 1520.120 ;
        RECT 4.400 1511.960 1741.495 1513.360 ;
        RECT 1.905 1505.880 1741.495 1511.960 ;
        RECT 4.400 1504.480 1741.495 1505.880 ;
        RECT 1.905 1497.720 1741.495 1504.480 ;
        RECT 4.400 1496.320 1741.495 1497.720 ;
        RECT 1.905 1490.240 1741.495 1496.320 ;
        RECT 4.400 1488.840 1741.495 1490.240 ;
        RECT 1.905 1482.080 1741.495 1488.840 ;
        RECT 4.400 1480.680 1741.495 1482.080 ;
        RECT 1.905 1474.600 1741.495 1480.680 ;
        RECT 4.400 1473.200 1741.495 1474.600 ;
        RECT 1.905 1466.440 1741.495 1473.200 ;
        RECT 4.400 1465.040 1741.495 1466.440 ;
        RECT 1.905 1458.960 1741.495 1465.040 ;
        RECT 4.400 1457.560 1741.495 1458.960 ;
        RECT 1.905 1450.800 1741.495 1457.560 ;
        RECT 4.400 1449.400 1741.495 1450.800 ;
        RECT 1.905 1443.320 1741.495 1449.400 ;
        RECT 4.400 1441.920 1741.495 1443.320 ;
        RECT 1.905 1435.160 1741.495 1441.920 ;
        RECT 4.400 1433.760 1741.495 1435.160 ;
        RECT 1.905 1427.680 1741.495 1433.760 ;
        RECT 4.400 1426.280 1741.495 1427.680 ;
        RECT 1.905 1419.520 1741.495 1426.280 ;
        RECT 4.400 1418.120 1741.495 1419.520 ;
        RECT 1.905 1412.040 1741.495 1418.120 ;
        RECT 4.400 1410.640 1741.495 1412.040 ;
        RECT 1.905 1403.880 1741.495 1410.640 ;
        RECT 4.400 1402.480 1741.495 1403.880 ;
        RECT 1.905 1396.400 1741.495 1402.480 ;
        RECT 4.400 1395.000 1741.495 1396.400 ;
        RECT 1.905 1388.240 1741.495 1395.000 ;
        RECT 4.400 1386.840 1741.495 1388.240 ;
        RECT 1.905 1380.760 1741.495 1386.840 ;
        RECT 4.400 1379.360 1741.495 1380.760 ;
        RECT 1.905 1372.600 1741.495 1379.360 ;
        RECT 4.400 1371.200 1741.495 1372.600 ;
        RECT 1.905 1365.120 1741.495 1371.200 ;
        RECT 4.400 1363.720 1741.495 1365.120 ;
        RECT 1.905 1356.960 1741.495 1363.720 ;
        RECT 4.400 1355.560 1741.495 1356.960 ;
        RECT 1.905 1349.480 1741.495 1355.560 ;
        RECT 4.400 1348.080 1741.495 1349.480 ;
        RECT 1.905 1341.320 1741.495 1348.080 ;
        RECT 4.400 1339.920 1741.495 1341.320 ;
        RECT 1.905 1333.840 1741.495 1339.920 ;
        RECT 4.400 1332.440 1741.495 1333.840 ;
        RECT 1.905 1325.680 1741.495 1332.440 ;
        RECT 4.400 1324.280 1741.495 1325.680 ;
        RECT 1.905 1318.200 1741.495 1324.280 ;
        RECT 4.400 1316.800 1741.495 1318.200 ;
        RECT 1.905 1310.040 1741.495 1316.800 ;
        RECT 4.400 1308.640 1741.495 1310.040 ;
        RECT 1.905 1302.560 1741.495 1308.640 ;
        RECT 4.400 1301.160 1741.495 1302.560 ;
        RECT 1.905 1294.400 1741.495 1301.160 ;
        RECT 4.400 1293.000 1741.495 1294.400 ;
        RECT 1.905 1286.920 1741.495 1293.000 ;
        RECT 4.400 1285.520 1741.495 1286.920 ;
        RECT 1.905 1278.760 1741.495 1285.520 ;
        RECT 4.400 1277.360 1741.495 1278.760 ;
        RECT 1.905 1271.280 1741.495 1277.360 ;
        RECT 4.400 1269.880 1741.495 1271.280 ;
        RECT 1.905 1263.120 1741.495 1269.880 ;
        RECT 4.400 1261.720 1741.495 1263.120 ;
        RECT 1.905 1255.640 1741.495 1261.720 ;
        RECT 4.400 1254.240 1741.495 1255.640 ;
        RECT 1.905 1247.480 1741.495 1254.240 ;
        RECT 4.400 1246.080 1741.495 1247.480 ;
        RECT 1.905 1240.000 1741.495 1246.080 ;
        RECT 4.400 1238.600 1741.495 1240.000 ;
        RECT 1.905 1231.840 1741.495 1238.600 ;
        RECT 4.400 1230.440 1741.495 1231.840 ;
        RECT 1.905 1224.360 1741.495 1230.440 ;
        RECT 4.400 1222.960 1741.495 1224.360 ;
        RECT 1.905 1216.200 1741.495 1222.960 ;
        RECT 4.400 1214.800 1741.495 1216.200 ;
        RECT 1.905 1208.720 1741.495 1214.800 ;
        RECT 4.400 1207.320 1741.495 1208.720 ;
        RECT 1.905 1200.560 1741.495 1207.320 ;
        RECT 4.400 1199.160 1741.495 1200.560 ;
        RECT 1.905 1193.080 1741.495 1199.160 ;
        RECT 4.400 1191.680 1741.495 1193.080 ;
        RECT 1.905 1184.920 1741.495 1191.680 ;
        RECT 4.400 1183.520 1741.495 1184.920 ;
        RECT 1.905 1177.440 1741.495 1183.520 ;
        RECT 4.400 1176.040 1741.495 1177.440 ;
        RECT 1.905 1169.280 1741.495 1176.040 ;
        RECT 4.400 1167.880 1741.495 1169.280 ;
        RECT 1.905 1161.800 1741.495 1167.880 ;
        RECT 4.400 1160.400 1741.495 1161.800 ;
        RECT 1.905 1153.640 1741.495 1160.400 ;
        RECT 4.400 1152.240 1741.495 1153.640 ;
        RECT 1.905 1146.160 1741.495 1152.240 ;
        RECT 4.400 1144.760 1741.495 1146.160 ;
        RECT 1.905 1138.000 1741.495 1144.760 ;
        RECT 4.400 1136.600 1741.495 1138.000 ;
        RECT 1.905 1130.520 1741.495 1136.600 ;
        RECT 4.400 1129.120 1741.495 1130.520 ;
        RECT 1.905 1122.360 1741.495 1129.120 ;
        RECT 4.400 1120.960 1741.495 1122.360 ;
        RECT 1.905 1114.880 1741.495 1120.960 ;
        RECT 4.400 1113.480 1741.495 1114.880 ;
        RECT 1.905 1106.720 1741.495 1113.480 ;
        RECT 4.400 1105.320 1741.495 1106.720 ;
        RECT 1.905 1099.240 1741.495 1105.320 ;
        RECT 4.400 1097.840 1741.495 1099.240 ;
        RECT 1.905 1091.080 1741.495 1097.840 ;
        RECT 4.400 1089.680 1741.495 1091.080 ;
        RECT 1.905 1083.600 1741.495 1089.680 ;
        RECT 4.400 1082.200 1741.495 1083.600 ;
        RECT 1.905 1075.440 1741.495 1082.200 ;
        RECT 4.400 1074.040 1741.495 1075.440 ;
        RECT 1.905 1067.960 1741.495 1074.040 ;
        RECT 4.400 1066.560 1741.495 1067.960 ;
        RECT 1.905 1059.800 1741.495 1066.560 ;
        RECT 4.400 1058.400 1741.495 1059.800 ;
        RECT 1.905 1052.320 1741.495 1058.400 ;
        RECT 4.400 1050.920 1741.495 1052.320 ;
        RECT 1.905 1044.160 1741.495 1050.920 ;
        RECT 4.400 1042.760 1741.495 1044.160 ;
        RECT 1.905 1036.680 1741.495 1042.760 ;
        RECT 4.400 1035.280 1741.495 1036.680 ;
        RECT 1.905 1028.520 1741.495 1035.280 ;
        RECT 4.400 1027.120 1741.495 1028.520 ;
        RECT 1.905 1021.040 1741.495 1027.120 ;
        RECT 4.400 1019.640 1741.495 1021.040 ;
        RECT 1.905 1012.880 1741.495 1019.640 ;
        RECT 4.400 1011.480 1741.495 1012.880 ;
        RECT 1.905 1005.400 1741.495 1011.480 ;
        RECT 4.400 1004.000 1741.495 1005.400 ;
        RECT 1.905 997.240 1741.495 1004.000 ;
        RECT 4.400 995.840 1741.495 997.240 ;
        RECT 1.905 989.760 1741.495 995.840 ;
        RECT 4.400 988.360 1741.495 989.760 ;
        RECT 1.905 981.600 1741.495 988.360 ;
        RECT 4.400 980.200 1741.495 981.600 ;
        RECT 1.905 974.120 1741.495 980.200 ;
        RECT 4.400 972.720 1741.495 974.120 ;
        RECT 1.905 965.960 1741.495 972.720 ;
        RECT 4.400 964.560 1741.495 965.960 ;
        RECT 1.905 958.480 1741.495 964.560 ;
        RECT 4.400 957.080 1741.495 958.480 ;
        RECT 1.905 950.320 1741.495 957.080 ;
        RECT 4.400 948.920 1741.495 950.320 ;
        RECT 1.905 942.840 1741.495 948.920 ;
        RECT 4.400 941.440 1741.495 942.840 ;
        RECT 1.905 934.680 1741.495 941.440 ;
        RECT 4.400 933.280 1741.495 934.680 ;
        RECT 1.905 927.200 1741.495 933.280 ;
        RECT 4.400 925.800 1741.495 927.200 ;
        RECT 1.905 919.040 1741.495 925.800 ;
        RECT 4.400 917.640 1741.495 919.040 ;
        RECT 1.905 911.560 1741.495 917.640 ;
        RECT 4.400 910.160 1741.495 911.560 ;
        RECT 1.905 903.400 1741.495 910.160 ;
        RECT 4.400 902.000 1741.495 903.400 ;
        RECT 1.905 895.920 1741.495 902.000 ;
        RECT 4.400 894.520 1741.495 895.920 ;
        RECT 1.905 887.760 1741.495 894.520 ;
        RECT 4.400 886.360 1741.495 887.760 ;
        RECT 1.905 880.280 1741.495 886.360 ;
        RECT 4.400 878.880 1741.495 880.280 ;
        RECT 1.905 872.120 1741.495 878.880 ;
        RECT 4.400 870.720 1741.495 872.120 ;
        RECT 1.905 864.640 1741.495 870.720 ;
        RECT 4.400 863.240 1741.495 864.640 ;
        RECT 1.905 856.480 1741.495 863.240 ;
        RECT 4.400 855.080 1741.495 856.480 ;
        RECT 1.905 849.000 1741.495 855.080 ;
        RECT 4.400 847.600 1741.495 849.000 ;
        RECT 1.905 840.840 1741.495 847.600 ;
        RECT 4.400 839.440 1741.495 840.840 ;
        RECT 1.905 833.360 1741.495 839.440 ;
        RECT 4.400 831.960 1741.495 833.360 ;
        RECT 1.905 825.200 1741.495 831.960 ;
        RECT 4.400 823.800 1741.495 825.200 ;
        RECT 1.905 817.720 1741.495 823.800 ;
        RECT 4.400 816.320 1741.495 817.720 ;
        RECT 1.905 809.560 1741.495 816.320 ;
        RECT 4.400 808.160 1741.495 809.560 ;
        RECT 1.905 802.080 1741.495 808.160 ;
        RECT 4.400 800.680 1741.495 802.080 ;
        RECT 1.905 793.920 1741.495 800.680 ;
        RECT 4.400 792.520 1741.495 793.920 ;
        RECT 1.905 786.440 1741.495 792.520 ;
        RECT 4.400 785.040 1741.495 786.440 ;
        RECT 1.905 778.280 1741.495 785.040 ;
        RECT 4.400 776.880 1741.495 778.280 ;
        RECT 1.905 770.800 1741.495 776.880 ;
        RECT 4.400 769.400 1741.495 770.800 ;
        RECT 1.905 762.640 1741.495 769.400 ;
        RECT 4.400 761.240 1741.495 762.640 ;
        RECT 1.905 755.160 1741.495 761.240 ;
        RECT 4.400 753.760 1741.495 755.160 ;
        RECT 1.905 747.000 1741.495 753.760 ;
        RECT 4.400 745.600 1741.495 747.000 ;
        RECT 1.905 739.520 1741.495 745.600 ;
        RECT 4.400 738.120 1741.495 739.520 ;
        RECT 1.905 731.360 1741.495 738.120 ;
        RECT 4.400 729.960 1741.495 731.360 ;
        RECT 1.905 723.880 1741.495 729.960 ;
        RECT 4.400 722.480 1741.495 723.880 ;
        RECT 1.905 715.720 1741.495 722.480 ;
        RECT 4.400 714.320 1741.495 715.720 ;
        RECT 1.905 708.240 1741.495 714.320 ;
        RECT 4.400 706.840 1741.495 708.240 ;
        RECT 1.905 700.080 1741.495 706.840 ;
        RECT 4.400 698.680 1741.495 700.080 ;
        RECT 1.905 692.600 1741.495 698.680 ;
        RECT 4.400 691.200 1741.495 692.600 ;
        RECT 1.905 684.440 1741.495 691.200 ;
        RECT 4.400 683.040 1741.495 684.440 ;
        RECT 1.905 676.960 1741.495 683.040 ;
        RECT 4.400 675.560 1741.495 676.960 ;
        RECT 1.905 668.800 1741.495 675.560 ;
        RECT 4.400 667.400 1741.495 668.800 ;
        RECT 1.905 661.320 1741.495 667.400 ;
        RECT 4.400 659.920 1741.495 661.320 ;
        RECT 1.905 653.160 1741.495 659.920 ;
        RECT 4.400 651.760 1741.495 653.160 ;
        RECT 1.905 645.680 1741.495 651.760 ;
        RECT 4.400 644.280 1741.495 645.680 ;
        RECT 1.905 637.520 1741.495 644.280 ;
        RECT 4.400 636.120 1741.495 637.520 ;
        RECT 1.905 630.040 1741.495 636.120 ;
        RECT 4.400 628.640 1741.495 630.040 ;
        RECT 1.905 621.880 1741.495 628.640 ;
        RECT 4.400 620.480 1741.495 621.880 ;
        RECT 1.905 614.400 1741.495 620.480 ;
        RECT 4.400 613.000 1741.495 614.400 ;
        RECT 1.905 606.240 1741.495 613.000 ;
        RECT 4.400 604.840 1741.495 606.240 ;
        RECT 1.905 598.760 1741.495 604.840 ;
        RECT 4.400 597.360 1741.495 598.760 ;
        RECT 1.905 590.600 1741.495 597.360 ;
        RECT 4.400 589.200 1741.495 590.600 ;
        RECT 1.905 583.120 1741.495 589.200 ;
        RECT 4.400 581.720 1741.495 583.120 ;
        RECT 1.905 574.960 1741.495 581.720 ;
        RECT 4.400 573.560 1741.495 574.960 ;
        RECT 1.905 567.480 1741.495 573.560 ;
        RECT 4.400 566.080 1741.495 567.480 ;
        RECT 1.905 559.320 1741.495 566.080 ;
        RECT 4.400 557.920 1741.495 559.320 ;
        RECT 1.905 551.840 1741.495 557.920 ;
        RECT 4.400 550.440 1741.495 551.840 ;
        RECT 1.905 543.680 1741.495 550.440 ;
        RECT 4.400 542.280 1741.495 543.680 ;
        RECT 1.905 536.200 1741.495 542.280 ;
        RECT 4.400 534.800 1741.495 536.200 ;
        RECT 1.905 528.040 1741.495 534.800 ;
        RECT 4.400 526.640 1741.495 528.040 ;
        RECT 1.905 520.560 1741.495 526.640 ;
        RECT 4.400 519.160 1741.495 520.560 ;
        RECT 1.905 512.400 1741.495 519.160 ;
        RECT 4.400 511.000 1741.495 512.400 ;
        RECT 1.905 504.920 1741.495 511.000 ;
        RECT 4.400 503.520 1741.495 504.920 ;
        RECT 1.905 496.760 1741.495 503.520 ;
        RECT 4.400 495.360 1741.495 496.760 ;
        RECT 1.905 489.280 1741.495 495.360 ;
        RECT 4.400 487.880 1741.495 489.280 ;
        RECT 1.905 481.120 1741.495 487.880 ;
        RECT 4.400 479.720 1741.495 481.120 ;
        RECT 1.905 473.640 1741.495 479.720 ;
        RECT 4.400 472.240 1741.495 473.640 ;
        RECT 1.905 465.480 1741.495 472.240 ;
        RECT 4.400 464.080 1741.495 465.480 ;
        RECT 1.905 458.000 1741.495 464.080 ;
        RECT 4.400 456.600 1741.495 458.000 ;
        RECT 1.905 449.840 1741.495 456.600 ;
        RECT 4.400 448.440 1741.495 449.840 ;
        RECT 1.905 442.360 1741.495 448.440 ;
        RECT 4.400 440.960 1741.495 442.360 ;
        RECT 1.905 434.200 1741.495 440.960 ;
        RECT 4.400 432.800 1741.495 434.200 ;
        RECT 1.905 426.720 1741.495 432.800 ;
        RECT 4.400 425.320 1741.495 426.720 ;
        RECT 1.905 418.560 1741.495 425.320 ;
        RECT 4.400 417.160 1741.495 418.560 ;
        RECT 1.905 411.080 1741.495 417.160 ;
        RECT 4.400 409.680 1741.495 411.080 ;
        RECT 1.905 402.920 1741.495 409.680 ;
        RECT 4.400 401.520 1741.495 402.920 ;
        RECT 1.905 395.440 1741.495 401.520 ;
        RECT 4.400 394.040 1741.495 395.440 ;
        RECT 1.905 387.280 1741.495 394.040 ;
        RECT 4.400 385.880 1741.495 387.280 ;
        RECT 1.905 379.800 1741.495 385.880 ;
        RECT 4.400 378.400 1741.495 379.800 ;
        RECT 1.905 371.640 1741.495 378.400 ;
        RECT 4.400 370.240 1741.495 371.640 ;
        RECT 1.905 364.160 1741.495 370.240 ;
        RECT 4.400 362.760 1741.495 364.160 ;
        RECT 1.905 356.000 1741.495 362.760 ;
        RECT 4.400 354.600 1741.495 356.000 ;
        RECT 1.905 348.520 1741.495 354.600 ;
        RECT 4.400 347.120 1741.495 348.520 ;
        RECT 1.905 340.360 1741.495 347.120 ;
        RECT 4.400 338.960 1741.495 340.360 ;
        RECT 1.905 332.880 1741.495 338.960 ;
        RECT 4.400 331.480 1741.495 332.880 ;
        RECT 1.905 324.720 1741.495 331.480 ;
        RECT 4.400 323.320 1741.495 324.720 ;
        RECT 1.905 317.240 1741.495 323.320 ;
        RECT 4.400 315.840 1741.495 317.240 ;
        RECT 1.905 309.080 1741.495 315.840 ;
        RECT 4.400 307.680 1741.495 309.080 ;
        RECT 1.905 301.600 1741.495 307.680 ;
        RECT 4.400 300.200 1741.495 301.600 ;
        RECT 1.905 293.440 1741.495 300.200 ;
        RECT 4.400 292.040 1741.495 293.440 ;
        RECT 1.905 285.960 1741.495 292.040 ;
        RECT 4.400 284.560 1741.495 285.960 ;
        RECT 1.905 277.800 1741.495 284.560 ;
        RECT 4.400 276.400 1741.495 277.800 ;
        RECT 1.905 270.320 1741.495 276.400 ;
        RECT 4.400 268.920 1741.495 270.320 ;
        RECT 1.905 262.160 1741.495 268.920 ;
        RECT 4.400 260.760 1741.495 262.160 ;
        RECT 1.905 254.680 1741.495 260.760 ;
        RECT 4.400 253.280 1741.495 254.680 ;
        RECT 1.905 246.520 1741.495 253.280 ;
        RECT 4.400 245.120 1741.495 246.520 ;
        RECT 1.905 239.040 1741.495 245.120 ;
        RECT 4.400 237.640 1741.495 239.040 ;
        RECT 1.905 230.880 1741.495 237.640 ;
        RECT 4.400 229.480 1741.495 230.880 ;
        RECT 1.905 223.400 1741.495 229.480 ;
        RECT 4.400 222.000 1741.495 223.400 ;
        RECT 1.905 215.240 1741.495 222.000 ;
        RECT 4.400 213.840 1741.495 215.240 ;
        RECT 1.905 207.760 1741.495 213.840 ;
        RECT 4.400 206.360 1741.495 207.760 ;
        RECT 1.905 199.600 1741.495 206.360 ;
        RECT 4.400 198.200 1741.495 199.600 ;
        RECT 1.905 192.120 1741.495 198.200 ;
        RECT 4.400 190.720 1741.495 192.120 ;
        RECT 1.905 183.960 1741.495 190.720 ;
        RECT 4.400 182.560 1741.495 183.960 ;
        RECT 1.905 176.480 1741.495 182.560 ;
        RECT 4.400 175.080 1741.495 176.480 ;
        RECT 1.905 168.320 1741.495 175.080 ;
        RECT 4.400 166.920 1741.495 168.320 ;
        RECT 1.905 160.840 1741.495 166.920 ;
        RECT 4.400 159.440 1741.495 160.840 ;
        RECT 1.905 152.680 1741.495 159.440 ;
        RECT 4.400 151.280 1741.495 152.680 ;
        RECT 1.905 145.200 1741.495 151.280 ;
        RECT 4.400 143.800 1741.495 145.200 ;
        RECT 1.905 137.040 1741.495 143.800 ;
        RECT 4.400 135.640 1741.495 137.040 ;
        RECT 1.905 129.560 1741.495 135.640 ;
        RECT 4.400 128.160 1741.495 129.560 ;
        RECT 1.905 121.400 1741.495 128.160 ;
        RECT 4.400 120.000 1741.495 121.400 ;
        RECT 1.905 113.920 1741.495 120.000 ;
        RECT 4.400 112.520 1741.495 113.920 ;
        RECT 1.905 105.760 1741.495 112.520 ;
        RECT 4.400 104.360 1741.495 105.760 ;
        RECT 1.905 98.280 1741.495 104.360 ;
        RECT 4.400 96.880 1741.495 98.280 ;
        RECT 1.905 90.120 1741.495 96.880 ;
        RECT 4.400 88.720 1741.495 90.120 ;
        RECT 1.905 82.640 1741.495 88.720 ;
        RECT 4.400 81.240 1741.495 82.640 ;
        RECT 1.905 74.480 1741.495 81.240 ;
        RECT 4.400 73.080 1741.495 74.480 ;
        RECT 1.905 67.000 1741.495 73.080 ;
        RECT 4.400 65.600 1741.495 67.000 ;
        RECT 1.905 58.840 1741.495 65.600 ;
        RECT 4.400 57.440 1741.495 58.840 ;
        RECT 1.905 51.360 1741.495 57.440 ;
        RECT 4.400 49.960 1741.495 51.360 ;
        RECT 1.905 43.200 1741.495 49.960 ;
        RECT 4.400 41.800 1741.495 43.200 ;
        RECT 1.905 35.720 1741.495 41.800 ;
        RECT 4.400 34.320 1741.495 35.720 ;
        RECT 1.905 27.560 1741.495 34.320 ;
        RECT 4.400 26.160 1741.495 27.560 ;
        RECT 1.905 20.080 1741.495 26.160 ;
        RECT 4.400 18.680 1741.495 20.080 ;
        RECT 1.905 11.920 1741.495 18.680 ;
        RECT 4.400 10.520 1741.495 11.920 ;
        RECT 1.905 4.440 1741.495 10.520 ;
        RECT 4.400 3.590 1741.495 4.440 ;
      LAYER met4 ;
        RECT 2.135 1755.040 1733.905 1767.145 ;
        RECT 2.135 11.735 20.640 1755.040 ;
        RECT 23.040 11.735 97.440 1755.040 ;
        RECT 99.840 11.735 174.240 1755.040 ;
        RECT 176.640 11.735 251.040 1755.040 ;
        RECT 253.440 11.735 327.840 1755.040 ;
        RECT 330.240 11.735 404.640 1755.040 ;
        RECT 407.040 11.735 481.440 1755.040 ;
        RECT 483.840 11.735 558.240 1755.040 ;
        RECT 560.640 11.735 635.040 1755.040 ;
        RECT 637.440 11.735 711.840 1755.040 ;
        RECT 714.240 11.735 788.640 1755.040 ;
        RECT 791.040 11.735 865.440 1755.040 ;
        RECT 867.840 11.735 942.240 1755.040 ;
        RECT 944.640 11.735 1019.040 1755.040 ;
        RECT 1021.440 11.735 1095.840 1755.040 ;
        RECT 1098.240 11.735 1172.640 1755.040 ;
        RECT 1175.040 11.735 1249.440 1755.040 ;
        RECT 1251.840 11.735 1326.240 1755.040 ;
        RECT 1328.640 11.735 1403.040 1755.040 ;
        RECT 1405.440 11.735 1479.840 1755.040 ;
        RECT 1482.240 11.735 1556.640 1755.040 ;
        RECT 1559.040 11.735 1633.440 1755.040 ;
        RECT 1635.840 11.735 1710.240 1755.040 ;
        RECT 1712.640 11.735 1733.905 1755.040 ;
  END
END Marmot
END LIBRARY

