magic
tech sky130A
magscale 1 2
timestamp 1647763611
<< obsli1 >>
rect 1104 2159 352360 353073
<< obsm1 >>
rect 290 309448 353520 353796
rect 290 309148 353524 309448
rect 290 261848 353520 309148
rect 290 261480 353524 261848
rect 290 960 353520 261480
<< metal2 >>
rect 1490 354864 1546 355664
rect 4526 354864 4582 355664
rect 7654 354864 7710 355664
rect 10782 354864 10838 355664
rect 13818 354864 13874 355664
rect 16946 354864 17002 355664
rect 20074 354864 20130 355664
rect 23110 354864 23166 355664
rect 26238 354864 26294 355664
rect 29366 354864 29422 355664
rect 32494 354864 32550 355664
rect 35530 354864 35586 355664
rect 38658 354864 38714 355664
rect 41786 354864 41842 355664
rect 44822 354864 44878 355664
rect 47950 354864 48006 355664
rect 51078 354864 51134 355664
rect 54206 354864 54262 355664
rect 57242 354864 57298 355664
rect 60370 354864 60426 355664
rect 63498 354864 63554 355664
rect 66534 354864 66590 355664
rect 69662 354864 69718 355664
rect 72790 354864 72846 355664
rect 75918 354864 75974 355664
rect 78954 354864 79010 355664
rect 82082 354864 82138 355664
rect 85210 354864 85266 355664
rect 88246 354864 88302 355664
rect 91374 354864 91430 355664
rect 94502 354864 94558 355664
rect 97630 354864 97686 355664
rect 100666 354864 100722 355664
rect 103794 354864 103850 355664
rect 106922 354864 106978 355664
rect 109958 354864 110014 355664
rect 113086 354864 113142 355664
rect 116214 354864 116270 355664
rect 119342 354864 119398 355664
rect 122378 354864 122434 355664
rect 125506 354864 125562 355664
rect 128634 354864 128690 355664
rect 131670 354864 131726 355664
rect 134798 354864 134854 355664
rect 137926 354864 137982 355664
rect 140962 354864 141018 355664
rect 144090 354864 144146 355664
rect 147218 354864 147274 355664
rect 150346 354864 150402 355664
rect 153382 354864 153438 355664
rect 156510 354864 156566 355664
rect 159638 354864 159694 355664
rect 162674 354864 162730 355664
rect 165802 354864 165858 355664
rect 168930 354864 168986 355664
rect 172058 354864 172114 355664
rect 175094 354864 175150 355664
rect 178222 354864 178278 355664
rect 181350 354864 181406 355664
rect 184386 354864 184442 355664
rect 187514 354864 187570 355664
rect 190642 354864 190698 355664
rect 193770 354864 193826 355664
rect 196806 354864 196862 355664
rect 199934 354864 199990 355664
rect 203062 354864 203118 355664
rect 206098 354864 206154 355664
rect 209226 354864 209282 355664
rect 212354 354864 212410 355664
rect 215482 354864 215538 355664
rect 218518 354864 218574 355664
rect 221646 354864 221702 355664
rect 224774 354864 224830 355664
rect 227810 354864 227866 355664
rect 230938 354864 230994 355664
rect 234066 354864 234122 355664
rect 237194 354864 237250 355664
rect 240230 354864 240286 355664
rect 243358 354864 243414 355664
rect 246486 354864 246542 355664
rect 249522 354864 249578 355664
rect 252650 354864 252706 355664
rect 255778 354864 255834 355664
rect 258814 354864 258870 355664
rect 261942 354864 261998 355664
rect 265070 354864 265126 355664
rect 268198 354864 268254 355664
rect 271234 354864 271290 355664
rect 274362 354864 274418 355664
rect 277490 354864 277546 355664
rect 280526 354864 280582 355664
rect 283654 354864 283710 355664
rect 286782 354864 286838 355664
rect 289910 354864 289966 355664
rect 292946 354864 293002 355664
rect 296074 354864 296130 355664
rect 299202 354864 299258 355664
rect 302238 354864 302294 355664
rect 305366 354864 305422 355664
rect 308494 354864 308550 355664
rect 311622 354864 311678 355664
rect 314658 354864 314714 355664
rect 317786 354864 317842 355664
rect 320914 354864 320970 355664
rect 323950 354864 324006 355664
rect 327078 354864 327134 355664
rect 330206 354864 330262 355664
rect 333334 354864 333390 355664
rect 336370 354864 336426 355664
rect 339498 354864 339554 355664
rect 342626 354864 342682 355664
rect 345662 354864 345718 355664
rect 348790 354864 348846 355664
rect 351918 354864 351974 355664
rect 294 0 350 800
rect 938 0 994 800
rect 1674 0 1730 800
rect 2410 0 2466 800
rect 3146 0 3202 800
rect 3790 0 3846 800
rect 4526 0 4582 800
rect 5262 0 5318 800
rect 5998 0 6054 800
rect 6734 0 6790 800
rect 7378 0 7434 800
rect 8114 0 8170 800
rect 8850 0 8906 800
rect 9586 0 9642 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11702 0 11758 800
rect 12438 0 12494 800
rect 13174 0 13230 800
rect 13910 0 13966 800
rect 14554 0 14610 800
rect 15290 0 15346 800
rect 16026 0 16082 800
rect 16762 0 16818 800
rect 17498 0 17554 800
rect 18142 0 18198 800
rect 18878 0 18934 800
rect 19614 0 19670 800
rect 20350 0 20406 800
rect 21086 0 21142 800
rect 21730 0 21786 800
rect 22466 0 22522 800
rect 23202 0 23258 800
rect 23938 0 23994 800
rect 24674 0 24730 800
rect 25318 0 25374 800
rect 26054 0 26110 800
rect 26790 0 26846 800
rect 27526 0 27582 800
rect 28262 0 28318 800
rect 28906 0 28962 800
rect 29642 0 29698 800
rect 30378 0 30434 800
rect 31114 0 31170 800
rect 31758 0 31814 800
rect 32494 0 32550 800
rect 33230 0 33286 800
rect 33966 0 34022 800
rect 34702 0 34758 800
rect 35346 0 35402 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37554 0 37610 800
rect 38290 0 38346 800
rect 38934 0 38990 800
rect 39670 0 39726 800
rect 40406 0 40462 800
rect 41142 0 41198 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43258 0 43314 800
rect 43994 0 44050 800
rect 44730 0 44786 800
rect 45466 0 45522 800
rect 46110 0 46166 800
rect 46846 0 46902 800
rect 47582 0 47638 800
rect 48318 0 48374 800
rect 49054 0 49110 800
rect 49698 0 49754 800
rect 50434 0 50490 800
rect 51170 0 51226 800
rect 51906 0 51962 800
rect 52642 0 52698 800
rect 53286 0 53342 800
rect 54022 0 54078 800
rect 54758 0 54814 800
rect 55494 0 55550 800
rect 56230 0 56286 800
rect 56874 0 56930 800
rect 57610 0 57666 800
rect 58346 0 58402 800
rect 59082 0 59138 800
rect 59726 0 59782 800
rect 60462 0 60518 800
rect 61198 0 61254 800
rect 61934 0 61990 800
rect 62670 0 62726 800
rect 63314 0 63370 800
rect 64050 0 64106 800
rect 64786 0 64842 800
rect 65522 0 65578 800
rect 66258 0 66314 800
rect 66902 0 66958 800
rect 67638 0 67694 800
rect 68374 0 68430 800
rect 69110 0 69166 800
rect 69846 0 69902 800
rect 70490 0 70546 800
rect 71226 0 71282 800
rect 71962 0 72018 800
rect 72698 0 72754 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74814 0 74870 800
rect 75550 0 75606 800
rect 76286 0 76342 800
rect 77022 0 77078 800
rect 77666 0 77722 800
rect 78402 0 78458 800
rect 79138 0 79194 800
rect 79874 0 79930 800
rect 80610 0 80666 800
rect 81254 0 81310 800
rect 81990 0 82046 800
rect 82726 0 82782 800
rect 83462 0 83518 800
rect 84198 0 84254 800
rect 84842 0 84898 800
rect 85578 0 85634 800
rect 86314 0 86370 800
rect 87050 0 87106 800
rect 87786 0 87842 800
rect 88430 0 88486 800
rect 89166 0 89222 800
rect 89902 0 89958 800
rect 90638 0 90694 800
rect 91282 0 91338 800
rect 92018 0 92074 800
rect 92754 0 92810 800
rect 93490 0 93546 800
rect 94226 0 94282 800
rect 94870 0 94926 800
rect 95606 0 95662 800
rect 96342 0 96398 800
rect 97078 0 97134 800
rect 97814 0 97870 800
rect 98458 0 98514 800
rect 99194 0 99250 800
rect 99930 0 99986 800
rect 100666 0 100722 800
rect 101402 0 101458 800
rect 102046 0 102102 800
rect 102782 0 102838 800
rect 103518 0 103574 800
rect 104254 0 104310 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106370 0 106426 800
rect 107106 0 107162 800
rect 107842 0 107898 800
rect 108578 0 108634 800
rect 109222 0 109278 800
rect 109958 0 110014 800
rect 110694 0 110750 800
rect 111430 0 111486 800
rect 112166 0 112222 800
rect 112810 0 112866 800
rect 113546 0 113602 800
rect 114282 0 114338 800
rect 115018 0 115074 800
rect 115754 0 115810 800
rect 116398 0 116454 800
rect 117134 0 117190 800
rect 117870 0 117926 800
rect 118606 0 118662 800
rect 119250 0 119306 800
rect 119986 0 120042 800
rect 120722 0 120778 800
rect 121458 0 121514 800
rect 122194 0 122250 800
rect 122838 0 122894 800
rect 123574 0 123630 800
rect 124310 0 124366 800
rect 125046 0 125102 800
rect 125782 0 125838 800
rect 126426 0 126482 800
rect 127162 0 127218 800
rect 127898 0 127954 800
rect 128634 0 128690 800
rect 129370 0 129426 800
rect 130014 0 130070 800
rect 130750 0 130806 800
rect 131486 0 131542 800
rect 132222 0 132278 800
rect 132958 0 133014 800
rect 133602 0 133658 800
rect 134338 0 134394 800
rect 135074 0 135130 800
rect 135810 0 135866 800
rect 136546 0 136602 800
rect 137190 0 137246 800
rect 137926 0 137982 800
rect 138662 0 138718 800
rect 139398 0 139454 800
rect 140134 0 140190 800
rect 140778 0 140834 800
rect 141514 0 141570 800
rect 142250 0 142306 800
rect 142986 0 143042 800
rect 143722 0 143778 800
rect 144366 0 144422 800
rect 145102 0 145158 800
rect 145838 0 145894 800
rect 146574 0 146630 800
rect 147310 0 147366 800
rect 147954 0 148010 800
rect 148690 0 148746 800
rect 149426 0 149482 800
rect 150162 0 150218 800
rect 150806 0 150862 800
rect 151542 0 151598 800
rect 152278 0 152334 800
rect 153014 0 153070 800
rect 153750 0 153806 800
rect 154394 0 154450 800
rect 155130 0 155186 800
rect 155866 0 155922 800
rect 156602 0 156658 800
rect 157338 0 157394 800
rect 157982 0 158038 800
rect 158718 0 158774 800
rect 159454 0 159510 800
rect 160190 0 160246 800
rect 160926 0 160982 800
rect 161570 0 161626 800
rect 162306 0 162362 800
rect 163042 0 163098 800
rect 163778 0 163834 800
rect 164514 0 164570 800
rect 165158 0 165214 800
rect 165894 0 165950 800
rect 166630 0 166686 800
rect 167366 0 167422 800
rect 168102 0 168158 800
rect 168746 0 168802 800
rect 169482 0 169538 800
rect 170218 0 170274 800
rect 170954 0 171010 800
rect 171690 0 171746 800
rect 172334 0 172390 800
rect 173070 0 173126 800
rect 173806 0 173862 800
rect 174542 0 174598 800
rect 175278 0 175334 800
rect 175922 0 175978 800
rect 176658 0 176714 800
rect 177394 0 177450 800
rect 178130 0 178186 800
rect 178774 0 178830 800
rect 179510 0 179566 800
rect 180246 0 180302 800
rect 180982 0 181038 800
rect 181718 0 181774 800
rect 182362 0 182418 800
rect 183098 0 183154 800
rect 183834 0 183890 800
rect 184570 0 184626 800
rect 185306 0 185362 800
rect 185950 0 186006 800
rect 186686 0 186742 800
rect 187422 0 187478 800
rect 188158 0 188214 800
rect 188894 0 188950 800
rect 189538 0 189594 800
rect 190274 0 190330 800
rect 191010 0 191066 800
rect 191746 0 191802 800
rect 192482 0 192538 800
rect 193126 0 193182 800
rect 193862 0 193918 800
rect 194598 0 194654 800
rect 195334 0 195390 800
rect 196070 0 196126 800
rect 196714 0 196770 800
rect 197450 0 197506 800
rect 198186 0 198242 800
rect 198922 0 198978 800
rect 199658 0 199714 800
rect 200302 0 200358 800
rect 201038 0 201094 800
rect 201774 0 201830 800
rect 202510 0 202566 800
rect 203246 0 203302 800
rect 203890 0 203946 800
rect 204626 0 204682 800
rect 205362 0 205418 800
rect 206098 0 206154 800
rect 206742 0 206798 800
rect 207478 0 207534 800
rect 208214 0 208270 800
rect 208950 0 209006 800
rect 209686 0 209742 800
rect 210330 0 210386 800
rect 211066 0 211122 800
rect 211802 0 211858 800
rect 212538 0 212594 800
rect 213274 0 213330 800
rect 213918 0 213974 800
rect 214654 0 214710 800
rect 215390 0 215446 800
rect 216126 0 216182 800
rect 216862 0 216918 800
rect 217506 0 217562 800
rect 218242 0 218298 800
rect 218978 0 219034 800
rect 219714 0 219770 800
rect 220450 0 220506 800
rect 221094 0 221150 800
rect 221830 0 221886 800
rect 222566 0 222622 800
rect 223302 0 223358 800
rect 224038 0 224094 800
rect 224682 0 224738 800
rect 225418 0 225474 800
rect 226154 0 226210 800
rect 226890 0 226946 800
rect 227626 0 227682 800
rect 228270 0 228326 800
rect 229006 0 229062 800
rect 229742 0 229798 800
rect 230478 0 230534 800
rect 231214 0 231270 800
rect 231858 0 231914 800
rect 232594 0 232650 800
rect 233330 0 233386 800
rect 234066 0 234122 800
rect 234802 0 234858 800
rect 235446 0 235502 800
rect 236182 0 236238 800
rect 236918 0 236974 800
rect 237654 0 237710 800
rect 238298 0 238354 800
rect 239034 0 239090 800
rect 239770 0 239826 800
rect 240506 0 240562 800
rect 241242 0 241298 800
rect 241886 0 241942 800
rect 242622 0 242678 800
rect 243358 0 243414 800
rect 244094 0 244150 800
rect 244830 0 244886 800
rect 245474 0 245530 800
rect 246210 0 246266 800
rect 246946 0 247002 800
rect 247682 0 247738 800
rect 248418 0 248474 800
rect 249062 0 249118 800
rect 249798 0 249854 800
rect 250534 0 250590 800
rect 251270 0 251326 800
rect 252006 0 252062 800
rect 252650 0 252706 800
rect 253386 0 253442 800
rect 254122 0 254178 800
rect 254858 0 254914 800
rect 255594 0 255650 800
rect 256238 0 256294 800
rect 256974 0 257030 800
rect 257710 0 257766 800
rect 258446 0 258502 800
rect 259182 0 259238 800
rect 259826 0 259882 800
rect 260562 0 260618 800
rect 261298 0 261354 800
rect 262034 0 262090 800
rect 262770 0 262826 800
rect 263414 0 263470 800
rect 264150 0 264206 800
rect 264886 0 264942 800
rect 265622 0 265678 800
rect 266266 0 266322 800
rect 267002 0 267058 800
rect 267738 0 267794 800
rect 268474 0 268530 800
rect 269210 0 269266 800
rect 269854 0 269910 800
rect 270590 0 270646 800
rect 271326 0 271382 800
rect 272062 0 272118 800
rect 272798 0 272854 800
rect 273442 0 273498 800
rect 274178 0 274234 800
rect 274914 0 274970 800
rect 275650 0 275706 800
rect 276386 0 276442 800
rect 277030 0 277086 800
rect 277766 0 277822 800
rect 278502 0 278558 800
rect 279238 0 279294 800
rect 279974 0 280030 800
rect 280618 0 280674 800
rect 281354 0 281410 800
rect 282090 0 282146 800
rect 282826 0 282882 800
rect 283562 0 283618 800
rect 284206 0 284262 800
rect 284942 0 284998 800
rect 285678 0 285734 800
rect 286414 0 286470 800
rect 287150 0 287206 800
rect 287794 0 287850 800
rect 288530 0 288586 800
rect 289266 0 289322 800
rect 290002 0 290058 800
rect 290738 0 290794 800
rect 291382 0 291438 800
rect 292118 0 292174 800
rect 292854 0 292910 800
rect 293590 0 293646 800
rect 294326 0 294382 800
rect 294970 0 295026 800
rect 295706 0 295762 800
rect 296442 0 296498 800
rect 297178 0 297234 800
rect 297822 0 297878 800
rect 298558 0 298614 800
rect 299294 0 299350 800
rect 300030 0 300086 800
rect 300766 0 300822 800
rect 301410 0 301466 800
rect 302146 0 302202 800
rect 302882 0 302938 800
rect 303618 0 303674 800
rect 304354 0 304410 800
rect 304998 0 305054 800
rect 305734 0 305790 800
rect 306470 0 306526 800
rect 307206 0 307262 800
rect 307942 0 307998 800
rect 308586 0 308642 800
rect 309322 0 309378 800
rect 310058 0 310114 800
rect 310794 0 310850 800
rect 311530 0 311586 800
rect 312174 0 312230 800
rect 312910 0 312966 800
rect 313646 0 313702 800
rect 314382 0 314438 800
rect 315118 0 315174 800
rect 315762 0 315818 800
rect 316498 0 316554 800
rect 317234 0 317290 800
rect 317970 0 318026 800
rect 318706 0 318762 800
rect 319350 0 319406 800
rect 320086 0 320142 800
rect 320822 0 320878 800
rect 321558 0 321614 800
rect 322294 0 322350 800
rect 322938 0 322994 800
rect 323674 0 323730 800
rect 324410 0 324466 800
rect 325146 0 325202 800
rect 325790 0 325846 800
rect 326526 0 326582 800
rect 327262 0 327318 800
rect 327998 0 328054 800
rect 328734 0 328790 800
rect 329378 0 329434 800
rect 330114 0 330170 800
rect 330850 0 330906 800
rect 331586 0 331642 800
rect 332322 0 332378 800
rect 332966 0 333022 800
rect 333702 0 333758 800
rect 334438 0 334494 800
rect 335174 0 335230 800
rect 335910 0 335966 800
rect 336554 0 336610 800
rect 337290 0 337346 800
rect 338026 0 338082 800
rect 338762 0 338818 800
rect 339498 0 339554 800
rect 340142 0 340198 800
rect 340878 0 340934 800
rect 341614 0 341670 800
rect 342350 0 342406 800
rect 343086 0 343142 800
rect 343730 0 343786 800
rect 344466 0 344522 800
rect 345202 0 345258 800
rect 345938 0 345994 800
rect 346674 0 346730 800
rect 347318 0 347374 800
rect 348054 0 348110 800
rect 348790 0 348846 800
rect 349526 0 349582 800
rect 350262 0 350318 800
rect 350906 0 350962 800
rect 351642 0 351698 800
rect 352378 0 352434 800
rect 353114 0 353170 800
<< obsm2 >>
rect 294 354808 1434 355065
rect 1602 354808 4470 355065
rect 4638 354808 7598 355065
rect 7766 354808 10726 355065
rect 10894 354808 13762 355065
rect 13930 354808 16890 355065
rect 17058 354808 20018 355065
rect 20186 354808 23054 355065
rect 23222 354808 26182 355065
rect 26350 354808 29310 355065
rect 29478 354808 32438 355065
rect 32606 354808 35474 355065
rect 35642 354808 38602 355065
rect 38770 354808 41730 355065
rect 41898 354808 44766 355065
rect 44934 354808 47894 355065
rect 48062 354808 51022 355065
rect 51190 354808 54150 355065
rect 54318 354808 57186 355065
rect 57354 354808 60314 355065
rect 60482 354808 63442 355065
rect 63610 354808 66478 355065
rect 66646 354808 69606 355065
rect 69774 354808 72734 355065
rect 72902 354808 75862 355065
rect 76030 354808 78898 355065
rect 79066 354808 82026 355065
rect 82194 354808 85154 355065
rect 85322 354808 88190 355065
rect 88358 354808 91318 355065
rect 91486 354808 94446 355065
rect 94614 354808 97574 355065
rect 97742 354808 100610 355065
rect 100778 354808 103738 355065
rect 103906 354808 106866 355065
rect 107034 354808 109902 355065
rect 110070 354808 113030 355065
rect 113198 354808 116158 355065
rect 116326 354808 119286 355065
rect 119454 354808 122322 355065
rect 122490 354808 125450 355065
rect 125618 354808 128578 355065
rect 128746 354808 131614 355065
rect 131782 354808 134742 355065
rect 134910 354808 137870 355065
rect 138038 354808 140906 355065
rect 141074 354808 144034 355065
rect 144202 354808 147162 355065
rect 147330 354808 150290 355065
rect 150458 354808 153326 355065
rect 153494 354808 156454 355065
rect 156622 354808 159582 355065
rect 159750 354808 162618 355065
rect 162786 354808 165746 355065
rect 165914 354808 168874 355065
rect 169042 354808 172002 355065
rect 172170 354808 175038 355065
rect 175206 354808 178166 355065
rect 178334 354808 181294 355065
rect 181462 354808 184330 355065
rect 184498 354808 187458 355065
rect 187626 354808 190586 355065
rect 190754 354808 193714 355065
rect 193882 354808 196750 355065
rect 196918 354808 199878 355065
rect 200046 354808 203006 355065
rect 203174 354808 206042 355065
rect 206210 354808 209170 355065
rect 209338 354808 212298 355065
rect 212466 354808 215426 355065
rect 215594 354808 218462 355065
rect 218630 354808 221590 355065
rect 221758 354808 224718 355065
rect 224886 354808 227754 355065
rect 227922 354808 230882 355065
rect 231050 354808 234010 355065
rect 234178 354808 237138 355065
rect 237306 354808 240174 355065
rect 240342 354808 243302 355065
rect 243470 354808 246430 355065
rect 246598 354808 249466 355065
rect 249634 354808 252594 355065
rect 252762 354808 255722 355065
rect 255890 354808 258758 355065
rect 258926 354808 261886 355065
rect 262054 354808 265014 355065
rect 265182 354808 268142 355065
rect 268310 354808 271178 355065
rect 271346 354808 274306 355065
rect 274474 354808 277434 355065
rect 277602 354808 280470 355065
rect 280638 354808 283598 355065
rect 283766 354808 286726 355065
rect 286894 354808 289854 355065
rect 290022 354808 292890 355065
rect 293058 354808 296018 355065
rect 296186 354808 299146 355065
rect 299314 354808 302182 355065
rect 302350 354808 305310 355065
rect 305478 354808 308438 355065
rect 308606 354808 311566 355065
rect 311734 354808 314602 355065
rect 314770 354808 317730 355065
rect 317898 354808 320858 355065
rect 321026 354808 323894 355065
rect 324062 354808 327022 355065
rect 327190 354808 330150 355065
rect 330318 354808 333278 355065
rect 333446 354808 336314 355065
rect 336482 354808 339442 355065
rect 339610 354808 342570 355065
rect 342738 354808 345606 355065
rect 345774 354808 348734 355065
rect 348902 354808 351862 355065
rect 352030 354808 353520 355065
rect 294 318866 353520 354808
rect 294 287388 353524 318866
rect 294 278774 353520 287388
rect 294 261582 353524 278774
rect 294 162364 353520 261582
rect 294 148532 353524 162364
rect 294 144914 353520 148532
rect 294 143500 353524 144914
rect 294 143392 353520 143500
rect 294 132960 353524 143392
rect 294 130778 353520 132960
rect 294 119360 353524 130778
rect 294 119218 353520 119360
rect 294 114328 353524 119218
rect 294 108372 353520 114328
rect 294 84166 353524 108372
rect 294 856 353520 84166
rect 406 303 882 856
rect 1050 303 1618 856
rect 1786 303 2354 856
rect 2522 303 3090 856
rect 3258 303 3734 856
rect 3902 303 4470 856
rect 4638 303 5206 856
rect 5374 303 5942 856
rect 6110 303 6678 856
rect 6846 303 7322 856
rect 7490 303 8058 856
rect 8226 303 8794 856
rect 8962 303 9530 856
rect 9698 303 10266 856
rect 10434 303 10910 856
rect 11078 303 11646 856
rect 11814 303 12382 856
rect 12550 303 13118 856
rect 13286 303 13854 856
rect 14022 303 14498 856
rect 14666 303 15234 856
rect 15402 303 15970 856
rect 16138 303 16706 856
rect 16874 303 17442 856
rect 17610 303 18086 856
rect 18254 303 18822 856
rect 18990 303 19558 856
rect 19726 303 20294 856
rect 20462 303 21030 856
rect 21198 303 21674 856
rect 21842 303 22410 856
rect 22578 303 23146 856
rect 23314 303 23882 856
rect 24050 303 24618 856
rect 24786 303 25262 856
rect 25430 303 25998 856
rect 26166 303 26734 856
rect 26902 303 27470 856
rect 27638 303 28206 856
rect 28374 303 28850 856
rect 29018 303 29586 856
rect 29754 303 30322 856
rect 30490 303 31058 856
rect 31226 303 31702 856
rect 31870 303 32438 856
rect 32606 303 33174 856
rect 33342 303 33910 856
rect 34078 303 34646 856
rect 34814 303 35290 856
rect 35458 303 36026 856
rect 36194 303 36762 856
rect 36930 303 37498 856
rect 37666 303 38234 856
rect 38402 303 38878 856
rect 39046 303 39614 856
rect 39782 303 40350 856
rect 40518 303 41086 856
rect 41254 303 41822 856
rect 41990 303 42466 856
rect 42634 303 43202 856
rect 43370 303 43938 856
rect 44106 303 44674 856
rect 44842 303 45410 856
rect 45578 303 46054 856
rect 46222 303 46790 856
rect 46958 303 47526 856
rect 47694 303 48262 856
rect 48430 303 48998 856
rect 49166 303 49642 856
rect 49810 303 50378 856
rect 50546 303 51114 856
rect 51282 303 51850 856
rect 52018 303 52586 856
rect 52754 303 53230 856
rect 53398 303 53966 856
rect 54134 303 54702 856
rect 54870 303 55438 856
rect 55606 303 56174 856
rect 56342 303 56818 856
rect 56986 303 57554 856
rect 57722 303 58290 856
rect 58458 303 59026 856
rect 59194 303 59670 856
rect 59838 303 60406 856
rect 60574 303 61142 856
rect 61310 303 61878 856
rect 62046 303 62614 856
rect 62782 303 63258 856
rect 63426 303 63994 856
rect 64162 303 64730 856
rect 64898 303 65466 856
rect 65634 303 66202 856
rect 66370 303 66846 856
rect 67014 303 67582 856
rect 67750 303 68318 856
rect 68486 303 69054 856
rect 69222 303 69790 856
rect 69958 303 70434 856
rect 70602 303 71170 856
rect 71338 303 71906 856
rect 72074 303 72642 856
rect 72810 303 73378 856
rect 73546 303 74022 856
rect 74190 303 74758 856
rect 74926 303 75494 856
rect 75662 303 76230 856
rect 76398 303 76966 856
rect 77134 303 77610 856
rect 77778 303 78346 856
rect 78514 303 79082 856
rect 79250 303 79818 856
rect 79986 303 80554 856
rect 80722 303 81198 856
rect 81366 303 81934 856
rect 82102 303 82670 856
rect 82838 303 83406 856
rect 83574 303 84142 856
rect 84310 303 84786 856
rect 84954 303 85522 856
rect 85690 303 86258 856
rect 86426 303 86994 856
rect 87162 303 87730 856
rect 87898 303 88374 856
rect 88542 303 89110 856
rect 89278 303 89846 856
rect 90014 303 90582 856
rect 90750 303 91226 856
rect 91394 303 91962 856
rect 92130 303 92698 856
rect 92866 303 93434 856
rect 93602 303 94170 856
rect 94338 303 94814 856
rect 94982 303 95550 856
rect 95718 303 96286 856
rect 96454 303 97022 856
rect 97190 303 97758 856
rect 97926 303 98402 856
rect 98570 303 99138 856
rect 99306 303 99874 856
rect 100042 303 100610 856
rect 100778 303 101346 856
rect 101514 303 101990 856
rect 102158 303 102726 856
rect 102894 303 103462 856
rect 103630 303 104198 856
rect 104366 303 104934 856
rect 105102 303 105578 856
rect 105746 303 106314 856
rect 106482 303 107050 856
rect 107218 303 107786 856
rect 107954 303 108522 856
rect 108690 303 109166 856
rect 109334 303 109902 856
rect 110070 303 110638 856
rect 110806 303 111374 856
rect 111542 303 112110 856
rect 112278 303 112754 856
rect 112922 303 113490 856
rect 113658 303 114226 856
rect 114394 303 114962 856
rect 115130 303 115698 856
rect 115866 303 116342 856
rect 116510 303 117078 856
rect 117246 303 117814 856
rect 117982 303 118550 856
rect 118718 303 119194 856
rect 119362 303 119930 856
rect 120098 303 120666 856
rect 120834 303 121402 856
rect 121570 303 122138 856
rect 122306 303 122782 856
rect 122950 303 123518 856
rect 123686 303 124254 856
rect 124422 303 124990 856
rect 125158 303 125726 856
rect 125894 303 126370 856
rect 126538 303 127106 856
rect 127274 303 127842 856
rect 128010 303 128578 856
rect 128746 303 129314 856
rect 129482 303 129958 856
rect 130126 303 130694 856
rect 130862 303 131430 856
rect 131598 303 132166 856
rect 132334 303 132902 856
rect 133070 303 133546 856
rect 133714 303 134282 856
rect 134450 303 135018 856
rect 135186 303 135754 856
rect 135922 303 136490 856
rect 136658 303 137134 856
rect 137302 303 137870 856
rect 138038 303 138606 856
rect 138774 303 139342 856
rect 139510 303 140078 856
rect 140246 303 140722 856
rect 140890 303 141458 856
rect 141626 303 142194 856
rect 142362 303 142930 856
rect 143098 303 143666 856
rect 143834 303 144310 856
rect 144478 303 145046 856
rect 145214 303 145782 856
rect 145950 303 146518 856
rect 146686 303 147254 856
rect 147422 303 147898 856
rect 148066 303 148634 856
rect 148802 303 149370 856
rect 149538 303 150106 856
rect 150274 303 150750 856
rect 150918 303 151486 856
rect 151654 303 152222 856
rect 152390 303 152958 856
rect 153126 303 153694 856
rect 153862 303 154338 856
rect 154506 303 155074 856
rect 155242 303 155810 856
rect 155978 303 156546 856
rect 156714 303 157282 856
rect 157450 303 157926 856
rect 158094 303 158662 856
rect 158830 303 159398 856
rect 159566 303 160134 856
rect 160302 303 160870 856
rect 161038 303 161514 856
rect 161682 303 162250 856
rect 162418 303 162986 856
rect 163154 303 163722 856
rect 163890 303 164458 856
rect 164626 303 165102 856
rect 165270 303 165838 856
rect 166006 303 166574 856
rect 166742 303 167310 856
rect 167478 303 168046 856
rect 168214 303 168690 856
rect 168858 303 169426 856
rect 169594 303 170162 856
rect 170330 303 170898 856
rect 171066 303 171634 856
rect 171802 303 172278 856
rect 172446 303 173014 856
rect 173182 303 173750 856
rect 173918 303 174486 856
rect 174654 303 175222 856
rect 175390 303 175866 856
rect 176034 303 176602 856
rect 176770 303 177338 856
rect 177506 303 178074 856
rect 178242 303 178718 856
rect 178886 303 179454 856
rect 179622 303 180190 856
rect 180358 303 180926 856
rect 181094 303 181662 856
rect 181830 303 182306 856
rect 182474 303 183042 856
rect 183210 303 183778 856
rect 183946 303 184514 856
rect 184682 303 185250 856
rect 185418 303 185894 856
rect 186062 303 186630 856
rect 186798 303 187366 856
rect 187534 303 188102 856
rect 188270 303 188838 856
rect 189006 303 189482 856
rect 189650 303 190218 856
rect 190386 303 190954 856
rect 191122 303 191690 856
rect 191858 303 192426 856
rect 192594 303 193070 856
rect 193238 303 193806 856
rect 193974 303 194542 856
rect 194710 303 195278 856
rect 195446 303 196014 856
rect 196182 303 196658 856
rect 196826 303 197394 856
rect 197562 303 198130 856
rect 198298 303 198866 856
rect 199034 303 199602 856
rect 199770 303 200246 856
rect 200414 303 200982 856
rect 201150 303 201718 856
rect 201886 303 202454 856
rect 202622 303 203190 856
rect 203358 303 203834 856
rect 204002 303 204570 856
rect 204738 303 205306 856
rect 205474 303 206042 856
rect 206210 303 206686 856
rect 206854 303 207422 856
rect 207590 303 208158 856
rect 208326 303 208894 856
rect 209062 303 209630 856
rect 209798 303 210274 856
rect 210442 303 211010 856
rect 211178 303 211746 856
rect 211914 303 212482 856
rect 212650 303 213218 856
rect 213386 303 213862 856
rect 214030 303 214598 856
rect 214766 303 215334 856
rect 215502 303 216070 856
rect 216238 303 216806 856
rect 216974 303 217450 856
rect 217618 303 218186 856
rect 218354 303 218922 856
rect 219090 303 219658 856
rect 219826 303 220394 856
rect 220562 303 221038 856
rect 221206 303 221774 856
rect 221942 303 222510 856
rect 222678 303 223246 856
rect 223414 303 223982 856
rect 224150 303 224626 856
rect 224794 303 225362 856
rect 225530 303 226098 856
rect 226266 303 226834 856
rect 227002 303 227570 856
rect 227738 303 228214 856
rect 228382 303 228950 856
rect 229118 303 229686 856
rect 229854 303 230422 856
rect 230590 303 231158 856
rect 231326 303 231802 856
rect 231970 303 232538 856
rect 232706 303 233274 856
rect 233442 303 234010 856
rect 234178 303 234746 856
rect 234914 303 235390 856
rect 235558 303 236126 856
rect 236294 303 236862 856
rect 237030 303 237598 856
rect 237766 303 238242 856
rect 238410 303 238978 856
rect 239146 303 239714 856
rect 239882 303 240450 856
rect 240618 303 241186 856
rect 241354 303 241830 856
rect 241998 303 242566 856
rect 242734 303 243302 856
rect 243470 303 244038 856
rect 244206 303 244774 856
rect 244942 303 245418 856
rect 245586 303 246154 856
rect 246322 303 246890 856
rect 247058 303 247626 856
rect 247794 303 248362 856
rect 248530 303 249006 856
rect 249174 303 249742 856
rect 249910 303 250478 856
rect 250646 303 251214 856
rect 251382 303 251950 856
rect 252118 303 252594 856
rect 252762 303 253330 856
rect 253498 303 254066 856
rect 254234 303 254802 856
rect 254970 303 255538 856
rect 255706 303 256182 856
rect 256350 303 256918 856
rect 257086 303 257654 856
rect 257822 303 258390 856
rect 258558 303 259126 856
rect 259294 303 259770 856
rect 259938 303 260506 856
rect 260674 303 261242 856
rect 261410 303 261978 856
rect 262146 303 262714 856
rect 262882 303 263358 856
rect 263526 303 264094 856
rect 264262 303 264830 856
rect 264998 303 265566 856
rect 265734 303 266210 856
rect 266378 303 266946 856
rect 267114 303 267682 856
rect 267850 303 268418 856
rect 268586 303 269154 856
rect 269322 303 269798 856
rect 269966 303 270534 856
rect 270702 303 271270 856
rect 271438 303 272006 856
rect 272174 303 272742 856
rect 272910 303 273386 856
rect 273554 303 274122 856
rect 274290 303 274858 856
rect 275026 303 275594 856
rect 275762 303 276330 856
rect 276498 303 276974 856
rect 277142 303 277710 856
rect 277878 303 278446 856
rect 278614 303 279182 856
rect 279350 303 279918 856
rect 280086 303 280562 856
rect 280730 303 281298 856
rect 281466 303 282034 856
rect 282202 303 282770 856
rect 282938 303 283506 856
rect 283674 303 284150 856
rect 284318 303 284886 856
rect 285054 303 285622 856
rect 285790 303 286358 856
rect 286526 303 287094 856
rect 287262 303 287738 856
rect 287906 303 288474 856
rect 288642 303 289210 856
rect 289378 303 289946 856
rect 290114 303 290682 856
rect 290850 303 291326 856
rect 291494 303 292062 856
rect 292230 303 292798 856
rect 292966 303 293534 856
rect 293702 303 294270 856
rect 294438 303 294914 856
rect 295082 303 295650 856
rect 295818 303 296386 856
rect 296554 303 297122 856
rect 297290 303 297766 856
rect 297934 303 298502 856
rect 298670 303 299238 856
rect 299406 303 299974 856
rect 300142 303 300710 856
rect 300878 303 301354 856
rect 301522 303 302090 856
rect 302258 303 302826 856
rect 302994 303 303562 856
rect 303730 303 304298 856
rect 304466 303 304942 856
rect 305110 303 305678 856
rect 305846 303 306414 856
rect 306582 303 307150 856
rect 307318 303 307886 856
rect 308054 303 308530 856
rect 308698 303 309266 856
rect 309434 303 310002 856
rect 310170 303 310738 856
rect 310906 303 311474 856
rect 311642 303 312118 856
rect 312286 303 312854 856
rect 313022 303 313590 856
rect 313758 303 314326 856
rect 314494 303 315062 856
rect 315230 303 315706 856
rect 315874 303 316442 856
rect 316610 303 317178 856
rect 317346 303 317914 856
rect 318082 303 318650 856
rect 318818 303 319294 856
rect 319462 303 320030 856
rect 320198 303 320766 856
rect 320934 303 321502 856
rect 321670 303 322238 856
rect 322406 303 322882 856
rect 323050 303 323618 856
rect 323786 303 324354 856
rect 324522 303 325090 856
rect 325258 303 325734 856
rect 325902 303 326470 856
rect 326638 303 327206 856
rect 327374 303 327942 856
rect 328110 303 328678 856
rect 328846 303 329322 856
rect 329490 303 330058 856
rect 330226 303 330794 856
rect 330962 303 331530 856
rect 331698 303 332266 856
rect 332434 303 332910 856
rect 333078 303 333646 856
rect 333814 303 334382 856
rect 334550 303 335118 856
rect 335286 303 335854 856
rect 336022 303 336498 856
rect 336666 303 337234 856
rect 337402 303 337970 856
rect 338138 303 338706 856
rect 338874 303 339442 856
rect 339610 303 340086 856
rect 340254 303 340822 856
rect 340990 303 341558 856
rect 341726 303 342294 856
rect 342462 303 343030 856
rect 343198 303 343674 856
rect 343842 303 344410 856
rect 344578 303 345146 856
rect 345314 303 345882 856
rect 346050 303 346618 856
rect 346786 303 347262 856
rect 347430 303 347998 856
rect 348166 303 348734 856
rect 348902 303 349470 856
rect 349638 303 350206 856
rect 350374 303 350850 856
rect 351018 303 351586 856
rect 351754 303 352322 856
rect 352490 303 353058 856
rect 353226 303 353520 856
<< metal3 >>
rect 0 355104 800 355224
rect 352720 354968 353520 355088
rect 0 354424 800 354544
rect 0 353744 800 353864
rect 352720 353880 353520 354000
rect 0 353064 800 353184
rect 352720 352792 353520 352912
rect 0 352384 800 352504
rect 0 351568 800 351688
rect 352720 351704 353520 351824
rect 0 350888 800 351008
rect 352720 350616 353520 350736
rect 0 350208 800 350328
rect 0 349528 800 349648
rect 352720 349528 353520 349648
rect 0 348848 800 348968
rect 352720 348440 353520 348560
rect 0 348168 800 348288
rect 0 347352 800 347472
rect 352720 347352 353520 347472
rect 0 346672 800 346792
rect 352720 346264 353520 346384
rect 0 345992 800 346112
rect 0 345312 800 345432
rect 352720 345176 353520 345296
rect 0 344632 800 344752
rect 352720 344088 353520 344208
rect 0 343816 800 343936
rect 0 343136 800 343256
rect 352720 343000 353520 343120
rect 0 342456 800 342576
rect 0 341776 800 341896
rect 352720 341912 353520 342032
rect 0 341096 800 341216
rect 352720 340824 353520 340944
rect 0 340416 800 340536
rect 0 339600 800 339720
rect 352720 339736 353520 339856
rect 0 338920 800 339040
rect 352720 338648 353520 338768
rect 0 338240 800 338360
rect 0 337560 800 337680
rect 352720 337560 353520 337680
rect 0 336880 800 337000
rect 352720 336472 353520 336592
rect 0 336200 800 336320
rect 0 335384 800 335504
rect 352720 335384 353520 335504
rect 0 334704 800 334824
rect 352720 334296 353520 334416
rect 0 334024 800 334144
rect 0 333344 800 333464
rect 352720 333208 353520 333328
rect 0 332664 800 332784
rect 352720 332120 353520 332240
rect 0 331848 800 331968
rect 0 331168 800 331288
rect 352720 331032 353520 331152
rect 0 330488 800 330608
rect 0 329808 800 329928
rect 352720 329944 353520 330064
rect 0 329128 800 329248
rect 352720 328856 353520 328976
rect 0 328448 800 328568
rect 0 327632 800 327752
rect 352720 327768 353520 327888
rect 0 326952 800 327072
rect 352720 326680 353520 326800
rect 0 326272 800 326392
rect 0 325592 800 325712
rect 352720 325592 353520 325712
rect 0 324912 800 325032
rect 352720 324504 353520 324624
rect 0 324096 800 324216
rect 0 323416 800 323536
rect 352720 323416 353520 323536
rect 0 322736 800 322856
rect 352720 322328 353520 322448
rect 0 322056 800 322176
rect 0 321376 800 321496
rect 352720 321240 353520 321360
rect 0 320696 800 320816
rect 352720 320152 353520 320272
rect 0 319880 800 320000
rect 0 319200 800 319320
rect 352720 319064 353520 319184
rect 0 318520 800 318640
rect 0 317840 800 317960
rect 352720 317976 353520 318096
rect 0 317160 800 317280
rect 352720 316888 353520 317008
rect 0 316480 800 316600
rect 352720 315936 353520 316056
rect 0 315664 800 315784
rect 0 314984 800 315104
rect 352720 314848 353520 314968
rect 0 314304 800 314424
rect 0 313624 800 313744
rect 352720 313760 353520 313880
rect 0 312944 800 313064
rect 352720 312672 353520 312792
rect 0 312128 800 312248
rect 0 311448 800 311568
rect 352720 311584 353520 311704
rect 0 310768 800 310888
rect 352720 310496 353520 310616
rect 0 310088 800 310208
rect 0 309408 800 309528
rect 352720 309408 353520 309528
rect 0 308728 800 308848
rect 352720 308320 353520 308440
rect 0 307912 800 308032
rect 0 307232 800 307352
rect 352720 307232 353520 307352
rect 0 306552 800 306672
rect 352720 306144 353520 306264
rect 0 305872 800 305992
rect 0 305192 800 305312
rect 352720 305056 353520 305176
rect 0 304376 800 304496
rect 352720 303968 353520 304088
rect 0 303696 800 303816
rect 0 303016 800 303136
rect 352720 302880 353520 303000
rect 0 302336 800 302456
rect 0 301656 800 301776
rect 352720 301792 353520 301912
rect 0 300976 800 301096
rect 352720 300704 353520 300824
rect 0 300160 800 300280
rect 0 299480 800 299600
rect 352720 299616 353520 299736
rect 0 298800 800 298920
rect 352720 298528 353520 298648
rect 0 298120 800 298240
rect 0 297440 800 297560
rect 352720 297440 353520 297560
rect 0 296760 800 296880
rect 352720 296352 353520 296472
rect 0 295944 800 296064
rect 0 295264 800 295384
rect 352720 295264 353520 295384
rect 0 294584 800 294704
rect 352720 294176 353520 294296
rect 0 293904 800 294024
rect 0 293224 800 293344
rect 352720 293088 353520 293208
rect 0 292408 800 292528
rect 352720 292000 353520 292120
rect 0 291728 800 291848
rect 0 291048 800 291168
rect 352720 290912 353520 291032
rect 0 290368 800 290488
rect 0 289688 800 289808
rect 352720 289824 353520 289944
rect 0 289008 800 289128
rect 352720 288736 353520 288856
rect 0 288192 800 288312
rect 0 287512 800 287632
rect 352720 287648 353520 287768
rect 0 286832 800 286952
rect 352720 286560 353520 286680
rect 0 286152 800 286272
rect 0 285472 800 285592
rect 352720 285472 353520 285592
rect 0 284792 800 284912
rect 352720 284384 353520 284504
rect 0 283976 800 284096
rect 0 283296 800 283416
rect 352720 283296 353520 283416
rect 0 282616 800 282736
rect 352720 282208 353520 282328
rect 0 281936 800 282056
rect 0 281256 800 281376
rect 352720 281120 353520 281240
rect 0 280440 800 280560
rect 352720 280032 353520 280152
rect 0 279760 800 279880
rect 0 279080 800 279200
rect 352720 278944 353520 279064
rect 0 278400 800 278520
rect 0 277720 800 277840
rect 352720 277856 353520 277976
rect 0 277040 800 277160
rect 352720 276904 353520 277024
rect 0 276224 800 276344
rect 352720 275816 353520 275936
rect 0 275544 800 275664
rect 0 274864 800 274984
rect 352720 274728 353520 274848
rect 0 274184 800 274304
rect 0 273504 800 273624
rect 352720 273640 353520 273760
rect 0 272688 800 272808
rect 352720 272552 353520 272672
rect 0 272008 800 272128
rect 0 271328 800 271448
rect 352720 271464 353520 271584
rect 0 270648 800 270768
rect 352720 270376 353520 270496
rect 0 269968 800 270088
rect 0 269288 800 269408
rect 352720 269288 353520 269408
rect 0 268472 800 268592
rect 352720 268200 353520 268320
rect 0 267792 800 267912
rect 0 267112 800 267232
rect 352720 267112 353520 267232
rect 0 266432 800 266552
rect 352720 266024 353520 266144
rect 0 265752 800 265872
rect 0 265072 800 265192
rect 352720 264936 353520 265056
rect 0 264256 800 264376
rect 352720 263848 353520 263968
rect 0 263576 800 263696
rect 0 262896 800 263016
rect 352720 262760 353520 262880
rect 0 262216 800 262336
rect 0 261536 800 261656
rect 352720 261672 353520 261792
rect 0 260720 800 260840
rect 352720 260584 353520 260704
rect 0 260040 800 260160
rect 0 259360 800 259480
rect 352720 259496 353520 259616
rect 0 258680 800 258800
rect 352720 258408 353520 258528
rect 0 258000 800 258120
rect 0 257320 800 257440
rect 352720 257320 353520 257440
rect 0 256504 800 256624
rect 352720 256232 353520 256352
rect 0 255824 800 255944
rect 0 255144 800 255264
rect 352720 255144 353520 255264
rect 0 254464 800 254584
rect 352720 254056 353520 254176
rect 0 253784 800 253904
rect 0 252968 800 253088
rect 352720 252968 353520 253088
rect 0 252288 800 252408
rect 352720 251880 353520 252000
rect 0 251608 800 251728
rect 0 250928 800 251048
rect 352720 250792 353520 250912
rect 0 250248 800 250368
rect 0 249568 800 249688
rect 352720 249704 353520 249824
rect 0 248752 800 248872
rect 352720 248616 353520 248736
rect 0 248072 800 248192
rect 0 247392 800 247512
rect 352720 247528 353520 247648
rect 0 246712 800 246832
rect 352720 246440 353520 246560
rect 0 246032 800 246152
rect 0 245352 800 245472
rect 352720 245352 353520 245472
rect 0 244536 800 244656
rect 352720 244264 353520 244384
rect 0 243856 800 243976
rect 0 243176 800 243296
rect 352720 243176 353520 243296
rect 0 242496 800 242616
rect 352720 242088 353520 242208
rect 0 241816 800 241936
rect 0 241000 800 241120
rect 352720 241000 353520 241120
rect 0 240320 800 240440
rect 352720 239912 353520 240032
rect 0 239640 800 239760
rect 0 238960 800 239080
rect 352720 238824 353520 238944
rect 0 238280 800 238400
rect 0 237600 800 237720
rect 352720 237736 353520 237856
rect 0 236784 800 236904
rect 352720 236784 353520 236904
rect 0 236104 800 236224
rect 352720 235696 353520 235816
rect 0 235424 800 235544
rect 0 234744 800 234864
rect 352720 234608 353520 234728
rect 0 234064 800 234184
rect 352720 233520 353520 233640
rect 0 233248 800 233368
rect 0 232568 800 232688
rect 352720 232432 353520 232552
rect 0 231888 800 232008
rect 0 231208 800 231328
rect 352720 231344 353520 231464
rect 0 230528 800 230648
rect 352720 230256 353520 230376
rect 0 229848 800 229968
rect 0 229032 800 229152
rect 352720 229168 353520 229288
rect 0 228352 800 228472
rect 352720 228080 353520 228200
rect 0 227672 800 227792
rect 0 226992 800 227112
rect 352720 226992 353520 227112
rect 0 226312 800 226432
rect 352720 225904 353520 226024
rect 0 225632 800 225752
rect 0 224816 800 224936
rect 352720 224816 353520 224936
rect 0 224136 800 224256
rect 352720 223728 353520 223848
rect 0 223456 800 223576
rect 0 222776 800 222896
rect 352720 222640 353520 222760
rect 0 222096 800 222216
rect 352720 221552 353520 221672
rect 0 221280 800 221400
rect 0 220600 800 220720
rect 352720 220464 353520 220584
rect 0 219920 800 220040
rect 0 219240 800 219360
rect 352720 219376 353520 219496
rect 0 218560 800 218680
rect 352720 218288 353520 218408
rect 0 217880 800 218000
rect 0 217064 800 217184
rect 352720 217200 353520 217320
rect 0 216384 800 216504
rect 352720 216112 353520 216232
rect 0 215704 800 215824
rect 0 215024 800 215144
rect 352720 215024 353520 215144
rect 0 214344 800 214464
rect 352720 213936 353520 214056
rect 0 213664 800 213784
rect 0 212848 800 212968
rect 352720 212848 353520 212968
rect 0 212168 800 212288
rect 352720 211760 353520 211880
rect 0 211488 800 211608
rect 0 210808 800 210928
rect 352720 210672 353520 210792
rect 0 210128 800 210248
rect 352720 209584 353520 209704
rect 0 209312 800 209432
rect 0 208632 800 208752
rect 352720 208496 353520 208616
rect 0 207952 800 208072
rect 0 207272 800 207392
rect 352720 207408 353520 207528
rect 0 206592 800 206712
rect 352720 206320 353520 206440
rect 0 205912 800 206032
rect 0 205096 800 205216
rect 352720 205232 353520 205352
rect 0 204416 800 204536
rect 352720 204144 353520 204264
rect 0 203736 800 203856
rect 0 203056 800 203176
rect 352720 203056 353520 203176
rect 0 202376 800 202496
rect 352720 201968 353520 202088
rect 0 201560 800 201680
rect 0 200880 800 201000
rect 352720 200880 353520 201000
rect 0 200200 800 200320
rect 352720 199792 353520 199912
rect 0 199520 800 199640
rect 0 198840 800 198960
rect 352720 198704 353520 198824
rect 0 198160 800 198280
rect 352720 197752 353520 197872
rect 0 197344 800 197464
rect 0 196664 800 196784
rect 352720 196664 353520 196784
rect 0 195984 800 196104
rect 352720 195576 353520 195696
rect 0 195304 800 195424
rect 0 194624 800 194744
rect 352720 194488 353520 194608
rect 0 193944 800 194064
rect 352720 193400 353520 193520
rect 0 193128 800 193248
rect 0 192448 800 192568
rect 352720 192312 353520 192432
rect 0 191768 800 191888
rect 0 191088 800 191208
rect 352720 191224 353520 191344
rect 0 190408 800 190528
rect 352720 190136 353520 190256
rect 0 189592 800 189712
rect 0 188912 800 189032
rect 352720 189048 353520 189168
rect 0 188232 800 188352
rect 352720 187960 353520 188080
rect 0 187552 800 187672
rect 0 186872 800 186992
rect 352720 186872 353520 186992
rect 0 186192 800 186312
rect 352720 185784 353520 185904
rect 0 185376 800 185496
rect 0 184696 800 184816
rect 352720 184696 353520 184816
rect 0 184016 800 184136
rect 352720 183608 353520 183728
rect 0 183336 800 183456
rect 0 182656 800 182776
rect 352720 182520 353520 182640
rect 0 181840 800 181960
rect 352720 181432 353520 181552
rect 0 181160 800 181280
rect 0 180480 800 180600
rect 352720 180344 353520 180464
rect 0 179800 800 179920
rect 0 179120 800 179240
rect 352720 179256 353520 179376
rect 0 178440 800 178560
rect 352720 178168 353520 178288
rect 0 177624 800 177744
rect 0 176944 800 177064
rect 352720 177080 353520 177200
rect 0 176264 800 176384
rect 352720 175992 353520 176112
rect 0 175584 800 175704
rect 0 174904 800 175024
rect 352720 174904 353520 175024
rect 0 174224 800 174344
rect 352720 173816 353520 173936
rect 0 173408 800 173528
rect 0 172728 800 172848
rect 352720 172728 353520 172848
rect 0 172048 800 172168
rect 352720 171640 353520 171760
rect 0 171368 800 171488
rect 0 170688 800 170808
rect 352720 170552 353520 170672
rect 0 169872 800 169992
rect 352720 169464 353520 169584
rect 0 169192 800 169312
rect 0 168512 800 168632
rect 352720 168376 353520 168496
rect 0 167832 800 167952
rect 0 167152 800 167272
rect 352720 167288 353520 167408
rect 0 166472 800 166592
rect 352720 166200 353520 166320
rect 0 165656 800 165776
rect 0 164976 800 165096
rect 352720 165112 353520 165232
rect 0 164296 800 164416
rect 352720 164024 353520 164144
rect 0 163616 800 163736
rect 0 162936 800 163056
rect 352720 162936 353520 163056
rect 0 162120 800 162240
rect 352720 161848 353520 161968
rect 0 161440 800 161560
rect 0 160760 800 160880
rect 352720 160760 353520 160880
rect 0 160080 800 160200
rect 352720 159672 353520 159792
rect 0 159400 800 159520
rect 0 158720 800 158840
rect 352720 158584 353520 158704
rect 0 157904 800 158024
rect 352720 157632 353520 157752
rect 0 157224 800 157344
rect 0 156544 800 156664
rect 352720 156544 353520 156664
rect 0 155864 800 155984
rect 352720 155456 353520 155576
rect 0 155184 800 155304
rect 0 154504 800 154624
rect 352720 154368 353520 154488
rect 0 153688 800 153808
rect 352720 153280 353520 153400
rect 0 153008 800 153128
rect 0 152328 800 152448
rect 352720 152192 353520 152312
rect 0 151648 800 151768
rect 0 150968 800 151088
rect 352720 151104 353520 151224
rect 0 150152 800 150272
rect 352720 150016 353520 150136
rect 0 149472 800 149592
rect 0 148792 800 148912
rect 352720 148928 353520 149048
rect 0 148112 800 148232
rect 352720 147840 353520 147960
rect 0 147432 800 147552
rect 0 146752 800 146872
rect 352720 146752 353520 146872
rect 0 145936 800 146056
rect 352720 145664 353520 145784
rect 0 145256 800 145376
rect 0 144576 800 144696
rect 352720 144576 353520 144696
rect 0 143896 800 144016
rect 352720 143488 353520 143608
rect 0 143216 800 143336
rect 0 142536 800 142656
rect 352720 142400 353520 142520
rect 0 141720 800 141840
rect 352720 141312 353520 141432
rect 0 141040 800 141160
rect 0 140360 800 140480
rect 352720 140224 353520 140344
rect 0 139680 800 139800
rect 0 139000 800 139120
rect 352720 139136 353520 139256
rect 0 138184 800 138304
rect 352720 138048 353520 138168
rect 0 137504 800 137624
rect 0 136824 800 136944
rect 352720 136960 353520 137080
rect 0 136144 800 136264
rect 352720 135872 353520 135992
rect 0 135464 800 135584
rect 0 134784 800 134904
rect 352720 134784 353520 134904
rect 0 133968 800 134088
rect 352720 133696 353520 133816
rect 0 133288 800 133408
rect 0 132608 800 132728
rect 352720 132608 353520 132728
rect 0 131928 800 132048
rect 352720 131520 353520 131640
rect 0 131248 800 131368
rect 0 130432 800 130552
rect 352720 130432 353520 130552
rect 0 129752 800 129872
rect 352720 129344 353520 129464
rect 0 129072 800 129192
rect 0 128392 800 128512
rect 352720 128256 353520 128376
rect 0 127712 800 127832
rect 0 127032 800 127152
rect 352720 127168 353520 127288
rect 0 126216 800 126336
rect 352720 126080 353520 126200
rect 0 125536 800 125656
rect 0 124856 800 124976
rect 352720 124992 353520 125112
rect 0 124176 800 124296
rect 352720 123904 353520 124024
rect 0 123496 800 123616
rect 0 122816 800 122936
rect 352720 122816 353520 122936
rect 0 122000 800 122120
rect 352720 121728 353520 121848
rect 0 121320 800 121440
rect 0 120640 800 120760
rect 352720 120640 353520 120760
rect 0 119960 800 120080
rect 352720 119552 353520 119672
rect 0 119280 800 119400
rect 0 118464 800 118584
rect 352720 118600 353520 118720
rect 0 117784 800 117904
rect 352720 117512 353520 117632
rect 0 117104 800 117224
rect 0 116424 800 116544
rect 352720 116424 353520 116544
rect 0 115744 800 115864
rect 352720 115336 353520 115456
rect 0 115064 800 115184
rect 0 114248 800 114368
rect 352720 114248 353520 114368
rect 0 113568 800 113688
rect 352720 113160 353520 113280
rect 0 112888 800 113008
rect 0 112208 800 112328
rect 352720 112072 353520 112192
rect 0 111528 800 111648
rect 352720 110984 353520 111104
rect 0 110712 800 110832
rect 0 110032 800 110152
rect 352720 109896 353520 110016
rect 0 109352 800 109472
rect 0 108672 800 108792
rect 352720 108808 353520 108928
rect 0 107992 800 108112
rect 352720 107720 353520 107840
rect 0 107312 800 107432
rect 0 106496 800 106616
rect 352720 106632 353520 106752
rect 0 105816 800 105936
rect 352720 105544 353520 105664
rect 0 105136 800 105256
rect 0 104456 800 104576
rect 352720 104456 353520 104576
rect 0 103776 800 103896
rect 352720 103368 353520 103488
rect 0 103096 800 103216
rect 0 102280 800 102400
rect 352720 102280 353520 102400
rect 0 101600 800 101720
rect 352720 101192 353520 101312
rect 0 100920 800 101040
rect 0 100240 800 100360
rect 352720 100104 353520 100224
rect 0 99560 800 99680
rect 352720 99016 353520 99136
rect 0 98744 800 98864
rect 0 98064 800 98184
rect 352720 97928 353520 98048
rect 0 97384 800 97504
rect 0 96704 800 96824
rect 352720 96840 353520 96960
rect 0 96024 800 96144
rect 352720 95752 353520 95872
rect 0 95344 800 95464
rect 0 94528 800 94648
rect 352720 94664 353520 94784
rect 0 93848 800 93968
rect 352720 93576 353520 93696
rect 0 93168 800 93288
rect 0 92488 800 92608
rect 352720 92488 353520 92608
rect 0 91808 800 91928
rect 352720 91400 353520 91520
rect 0 90992 800 91112
rect 0 90312 800 90432
rect 352720 90312 353520 90432
rect 0 89632 800 89752
rect 352720 89224 353520 89344
rect 0 88952 800 89072
rect 0 88272 800 88392
rect 352720 88136 353520 88256
rect 0 87592 800 87712
rect 352720 87048 353520 87168
rect 0 86776 800 86896
rect 0 86096 800 86216
rect 352720 85960 353520 86080
rect 0 85416 800 85536
rect 0 84736 800 84856
rect 352720 84872 353520 84992
rect 0 84056 800 84176
rect 352720 83784 353520 83904
rect 0 83376 800 83496
rect 0 82560 800 82680
rect 352720 82696 353520 82816
rect 0 81880 800 82000
rect 352720 81608 353520 81728
rect 0 81200 800 81320
rect 0 80520 800 80640
rect 352720 80520 353520 80640
rect 0 79840 800 79960
rect 352720 79432 353520 79552
rect 0 79024 800 79144
rect 0 78344 800 78464
rect 352720 78480 353520 78600
rect 0 77664 800 77784
rect 352720 77392 353520 77512
rect 0 76984 800 77104
rect 0 76304 800 76424
rect 352720 76304 353520 76424
rect 0 75624 800 75744
rect 352720 75216 353520 75336
rect 0 74808 800 74928
rect 0 74128 800 74248
rect 352720 74128 353520 74248
rect 0 73448 800 73568
rect 352720 73040 353520 73160
rect 0 72768 800 72888
rect 0 72088 800 72208
rect 352720 71952 353520 72072
rect 0 71408 800 71528
rect 352720 70864 353520 70984
rect 0 70592 800 70712
rect 0 69912 800 70032
rect 352720 69776 353520 69896
rect 0 69232 800 69352
rect 0 68552 800 68672
rect 352720 68688 353520 68808
rect 0 67872 800 67992
rect 352720 67600 353520 67720
rect 0 67056 800 67176
rect 0 66376 800 66496
rect 352720 66512 353520 66632
rect 0 65696 800 65816
rect 352720 65424 353520 65544
rect 0 65016 800 65136
rect 0 64336 800 64456
rect 352720 64336 353520 64456
rect 0 63656 800 63776
rect 352720 63248 353520 63368
rect 0 62840 800 62960
rect 0 62160 800 62280
rect 352720 62160 353520 62280
rect 0 61480 800 61600
rect 352720 61072 353520 61192
rect 0 60800 800 60920
rect 0 60120 800 60240
rect 352720 59984 353520 60104
rect 0 59304 800 59424
rect 352720 58896 353520 59016
rect 0 58624 800 58744
rect 0 57944 800 58064
rect 352720 57808 353520 57928
rect 0 57264 800 57384
rect 0 56584 800 56704
rect 352720 56720 353520 56840
rect 0 55904 800 56024
rect 352720 55632 353520 55752
rect 0 55088 800 55208
rect 0 54408 800 54528
rect 352720 54544 353520 54664
rect 0 53728 800 53848
rect 352720 53456 353520 53576
rect 0 53048 800 53168
rect 0 52368 800 52488
rect 352720 52368 353520 52488
rect 0 51688 800 51808
rect 352720 51280 353520 51400
rect 0 50872 800 50992
rect 0 50192 800 50312
rect 352720 50192 353520 50312
rect 0 49512 800 49632
rect 352720 49104 353520 49224
rect 0 48832 800 48952
rect 0 48152 800 48272
rect 352720 48016 353520 48136
rect 0 47336 800 47456
rect 352720 46928 353520 47048
rect 0 46656 800 46776
rect 0 45976 800 46096
rect 352720 45840 353520 45960
rect 0 45296 800 45416
rect 0 44616 800 44736
rect 352720 44752 353520 44872
rect 0 43936 800 44056
rect 352720 43664 353520 43784
rect 0 43120 800 43240
rect 0 42440 800 42560
rect 352720 42576 353520 42696
rect 0 41760 800 41880
rect 352720 41488 353520 41608
rect 0 41080 800 41200
rect 0 40400 800 40520
rect 352720 40400 353520 40520
rect 0 39584 800 39704
rect 352720 39448 353520 39568
rect 0 38904 800 39024
rect 0 38224 800 38344
rect 352720 38360 353520 38480
rect 0 37544 800 37664
rect 352720 37272 353520 37392
rect 0 36864 800 36984
rect 0 36184 800 36304
rect 352720 36184 353520 36304
rect 0 35368 800 35488
rect 352720 35096 353520 35216
rect 0 34688 800 34808
rect 0 34008 800 34128
rect 352720 34008 353520 34128
rect 0 33328 800 33448
rect 352720 32920 353520 33040
rect 0 32648 800 32768
rect 0 31968 800 32088
rect 352720 31832 353520 31952
rect 0 31152 800 31272
rect 352720 30744 353520 30864
rect 0 30472 800 30592
rect 0 29792 800 29912
rect 352720 29656 353520 29776
rect 0 29112 800 29232
rect 0 28432 800 28552
rect 352720 28568 353520 28688
rect 0 27616 800 27736
rect 352720 27480 353520 27600
rect 0 26936 800 27056
rect 0 26256 800 26376
rect 352720 26392 353520 26512
rect 0 25576 800 25696
rect 352720 25304 353520 25424
rect 0 24896 800 25016
rect 0 24216 800 24336
rect 352720 24216 353520 24336
rect 0 23400 800 23520
rect 352720 23128 353520 23248
rect 0 22720 800 22840
rect 0 22040 800 22160
rect 352720 22040 353520 22160
rect 0 21360 800 21480
rect 352720 20952 353520 21072
rect 0 20680 800 20800
rect 0 19864 800 19984
rect 352720 19864 353520 19984
rect 0 19184 800 19304
rect 352720 18776 353520 18896
rect 0 18504 800 18624
rect 0 17824 800 17944
rect 352720 17688 353520 17808
rect 0 17144 800 17264
rect 0 16464 800 16584
rect 352720 16600 353520 16720
rect 0 15648 800 15768
rect 352720 15512 353520 15632
rect 0 14968 800 15088
rect 0 14288 800 14408
rect 352720 14424 353520 14544
rect 0 13608 800 13728
rect 352720 13336 353520 13456
rect 0 12928 800 13048
rect 0 12248 800 12368
rect 352720 12248 353520 12368
rect 0 11432 800 11552
rect 352720 11160 353520 11280
rect 0 10752 800 10872
rect 0 10072 800 10192
rect 352720 10072 353520 10192
rect 0 9392 800 9512
rect 352720 8984 353520 9104
rect 0 8712 800 8832
rect 0 7896 800 8016
rect 352720 7896 353520 8016
rect 0 7216 800 7336
rect 352720 6808 353520 6928
rect 0 6536 800 6656
rect 0 5856 800 5976
rect 352720 5720 353520 5840
rect 0 5176 800 5296
rect 0 4496 800 4616
rect 352720 4632 353520 4752
rect 0 3680 800 3800
rect 352720 3544 353520 3664
rect 0 3000 800 3120
rect 0 2320 800 2440
rect 352720 2456 353520 2576
rect 0 1640 800 1760
rect 352720 1368 353520 1488
rect 0 960 800 1080
rect 0 280 800 400
rect 352720 416 353520 536
<< obsm3 >>
rect 880 355024 352640 355061
rect 289 354888 352640 355024
rect 289 354624 353451 354888
rect 880 354344 353451 354624
rect 289 354080 353451 354344
rect 289 353944 352640 354080
rect 880 353800 352640 353944
rect 880 353664 353451 353800
rect 289 353264 353451 353664
rect 880 352992 353451 353264
rect 880 352984 352640 352992
rect 289 352712 352640 352984
rect 289 352584 353451 352712
rect 880 352304 353451 352584
rect 289 351904 353451 352304
rect 289 351768 352640 351904
rect 880 351624 352640 351768
rect 880 351488 353451 351624
rect 289 351088 353451 351488
rect 880 350816 353451 351088
rect 880 350808 352640 350816
rect 289 350536 352640 350808
rect 289 350408 353451 350536
rect 880 350128 353451 350408
rect 289 349728 353451 350128
rect 880 349448 352640 349728
rect 289 349048 353451 349448
rect 880 348768 353451 349048
rect 289 348640 353451 348768
rect 289 348368 352640 348640
rect 880 348360 352640 348368
rect 880 348088 353451 348360
rect 289 347552 353451 348088
rect 880 347272 352640 347552
rect 289 346872 353451 347272
rect 880 346592 353451 346872
rect 289 346464 353451 346592
rect 289 346192 352640 346464
rect 880 346184 352640 346192
rect 880 345912 353451 346184
rect 289 345512 353451 345912
rect 880 345376 353451 345512
rect 880 345232 352640 345376
rect 289 345096 352640 345232
rect 289 344832 353451 345096
rect 880 344552 353451 344832
rect 289 344288 353451 344552
rect 289 344016 352640 344288
rect 880 344008 352640 344016
rect 880 343736 353451 344008
rect 289 343336 353451 343736
rect 880 343200 353451 343336
rect 880 343056 352640 343200
rect 289 342920 352640 343056
rect 289 342656 353451 342920
rect 880 342376 353451 342656
rect 289 342112 353451 342376
rect 289 341976 352640 342112
rect 880 341832 352640 341976
rect 880 341696 353451 341832
rect 289 341296 353451 341696
rect 880 341024 353451 341296
rect 880 341016 352640 341024
rect 289 340744 352640 341016
rect 289 340616 353451 340744
rect 880 340336 353451 340616
rect 289 339936 353451 340336
rect 289 339800 352640 339936
rect 880 339656 352640 339800
rect 880 339520 353451 339656
rect 289 339120 353451 339520
rect 880 338848 353451 339120
rect 880 338840 352640 338848
rect 289 338568 352640 338840
rect 289 338440 353451 338568
rect 880 338160 353451 338440
rect 289 337760 353451 338160
rect 880 337480 352640 337760
rect 289 337080 353451 337480
rect 880 336800 353451 337080
rect 289 336672 353451 336800
rect 289 336400 352640 336672
rect 880 336392 352640 336400
rect 880 336120 353451 336392
rect 289 335584 353451 336120
rect 880 335304 352640 335584
rect 289 334904 353451 335304
rect 880 334624 353451 334904
rect 289 334496 353451 334624
rect 289 334224 352640 334496
rect 880 334216 352640 334224
rect 880 333944 353451 334216
rect 289 333544 353451 333944
rect 880 333408 353451 333544
rect 880 333264 352640 333408
rect 289 333128 352640 333264
rect 289 332864 353451 333128
rect 880 332584 353451 332864
rect 289 332320 353451 332584
rect 289 332048 352640 332320
rect 880 332040 352640 332048
rect 880 331768 353451 332040
rect 289 331368 353451 331768
rect 880 331232 353451 331368
rect 880 331088 352640 331232
rect 289 330952 352640 331088
rect 289 330688 353451 330952
rect 880 330408 353451 330688
rect 289 330144 353451 330408
rect 289 330008 352640 330144
rect 880 329864 352640 330008
rect 880 329728 353451 329864
rect 289 329328 353451 329728
rect 880 329056 353451 329328
rect 880 329048 352640 329056
rect 289 328776 352640 329048
rect 289 328648 353451 328776
rect 880 328368 353451 328648
rect 289 327968 353451 328368
rect 289 327832 352640 327968
rect 880 327688 352640 327832
rect 880 327552 353451 327688
rect 289 327152 353451 327552
rect 880 326880 353451 327152
rect 880 326872 352640 326880
rect 289 326600 352640 326872
rect 289 326472 353451 326600
rect 880 326192 353451 326472
rect 289 325792 353451 326192
rect 880 325512 352640 325792
rect 289 325112 353451 325512
rect 880 324832 353451 325112
rect 289 324704 353451 324832
rect 289 324424 352640 324704
rect 289 324296 353451 324424
rect 880 324016 353451 324296
rect 289 323616 353451 324016
rect 880 323336 352640 323616
rect 289 322936 353451 323336
rect 880 322656 353451 322936
rect 289 322528 353451 322656
rect 289 322256 352640 322528
rect 880 322248 352640 322256
rect 880 321976 353451 322248
rect 289 321576 353451 321976
rect 880 321440 353451 321576
rect 880 321296 352640 321440
rect 289 321160 352640 321296
rect 289 320896 353451 321160
rect 880 320616 353451 320896
rect 289 320352 353451 320616
rect 289 320080 352640 320352
rect 880 320072 352640 320080
rect 880 319800 353451 320072
rect 289 319400 353451 319800
rect 880 319264 353451 319400
rect 880 319120 352640 319264
rect 289 318984 352640 319120
rect 289 318720 353451 318984
rect 880 318440 353451 318720
rect 289 318176 353451 318440
rect 289 318040 352640 318176
rect 880 317896 352640 318040
rect 880 317760 353451 317896
rect 289 317360 353451 317760
rect 880 317088 353451 317360
rect 880 317080 352640 317088
rect 289 316808 352640 317080
rect 289 316680 353451 316808
rect 880 316400 353451 316680
rect 289 316136 353451 316400
rect 289 315864 352640 316136
rect 880 315856 352640 315864
rect 880 315584 353451 315856
rect 289 315184 353451 315584
rect 880 315048 353451 315184
rect 880 314904 352640 315048
rect 289 314768 352640 314904
rect 289 314504 353451 314768
rect 880 314224 353451 314504
rect 289 313960 353451 314224
rect 289 313824 352640 313960
rect 880 313680 352640 313824
rect 880 313544 353451 313680
rect 289 313144 353451 313544
rect 880 312872 353451 313144
rect 880 312864 352640 312872
rect 289 312592 352640 312864
rect 289 312328 353451 312592
rect 880 312048 353451 312328
rect 289 311784 353451 312048
rect 289 311648 352640 311784
rect 880 311504 352640 311648
rect 880 311368 353451 311504
rect 289 310968 353451 311368
rect 880 310696 353451 310968
rect 880 310688 352640 310696
rect 289 310416 352640 310688
rect 289 310288 353451 310416
rect 880 310008 353451 310288
rect 289 309608 353451 310008
rect 880 309328 352640 309608
rect 289 308928 353451 309328
rect 880 308648 353451 308928
rect 289 308520 353451 308648
rect 289 308240 352640 308520
rect 289 308112 353451 308240
rect 880 307832 353451 308112
rect 289 307432 353451 307832
rect 880 307152 352640 307432
rect 289 306752 353451 307152
rect 880 306472 353451 306752
rect 289 306344 353451 306472
rect 289 306072 352640 306344
rect 880 306064 352640 306072
rect 880 305792 353451 306064
rect 289 305392 353451 305792
rect 880 305256 353451 305392
rect 880 305112 352640 305256
rect 289 304976 352640 305112
rect 289 304576 353451 304976
rect 880 304296 353451 304576
rect 289 304168 353451 304296
rect 289 303896 352640 304168
rect 880 303888 352640 303896
rect 880 303616 353451 303888
rect 289 303216 353451 303616
rect 880 303080 353451 303216
rect 880 302936 352640 303080
rect 289 302800 352640 302936
rect 289 302536 353451 302800
rect 880 302256 353451 302536
rect 289 301992 353451 302256
rect 289 301856 352640 301992
rect 880 301712 352640 301856
rect 880 301576 353451 301712
rect 289 301176 353451 301576
rect 880 300904 353451 301176
rect 880 300896 352640 300904
rect 289 300624 352640 300896
rect 289 300360 353451 300624
rect 880 300080 353451 300360
rect 289 299816 353451 300080
rect 289 299680 352640 299816
rect 880 299536 352640 299680
rect 880 299400 353451 299536
rect 289 299000 353451 299400
rect 880 298728 353451 299000
rect 880 298720 352640 298728
rect 289 298448 352640 298720
rect 289 298320 353451 298448
rect 880 298040 353451 298320
rect 289 297640 353451 298040
rect 880 297360 352640 297640
rect 289 296960 353451 297360
rect 880 296680 353451 296960
rect 289 296552 353451 296680
rect 289 296272 352640 296552
rect 289 296144 353451 296272
rect 880 295864 353451 296144
rect 289 295464 353451 295864
rect 880 295184 352640 295464
rect 289 294784 353451 295184
rect 880 294504 353451 294784
rect 289 294376 353451 294504
rect 289 294104 352640 294376
rect 880 294096 352640 294104
rect 880 293824 353451 294096
rect 289 293424 353451 293824
rect 880 293288 353451 293424
rect 880 293144 352640 293288
rect 289 293008 352640 293144
rect 289 292608 353451 293008
rect 880 292328 353451 292608
rect 289 292200 353451 292328
rect 289 291928 352640 292200
rect 880 291920 352640 291928
rect 880 291648 353451 291920
rect 289 291248 353451 291648
rect 880 291112 353451 291248
rect 880 290968 352640 291112
rect 289 290832 352640 290968
rect 289 290568 353451 290832
rect 880 290288 353451 290568
rect 289 290024 353451 290288
rect 289 289888 352640 290024
rect 880 289744 352640 289888
rect 880 289608 353451 289744
rect 289 289208 353451 289608
rect 880 288936 353451 289208
rect 880 288928 352640 288936
rect 289 288656 352640 288928
rect 289 288392 353451 288656
rect 880 288112 353451 288392
rect 289 287848 353451 288112
rect 289 287712 352640 287848
rect 880 287568 352640 287712
rect 880 287432 353451 287568
rect 289 287032 353451 287432
rect 880 286760 353451 287032
rect 880 286752 352640 286760
rect 289 286480 352640 286752
rect 289 286352 353451 286480
rect 880 286072 353451 286352
rect 289 285672 353451 286072
rect 880 285392 352640 285672
rect 289 284992 353451 285392
rect 880 284712 353451 284992
rect 289 284584 353451 284712
rect 289 284304 352640 284584
rect 289 284176 353451 284304
rect 880 283896 353451 284176
rect 289 283496 353451 283896
rect 880 283216 352640 283496
rect 289 282816 353451 283216
rect 880 282536 353451 282816
rect 289 282408 353451 282536
rect 289 282136 352640 282408
rect 880 282128 352640 282136
rect 880 281856 353451 282128
rect 289 281456 353451 281856
rect 880 281320 353451 281456
rect 880 281176 352640 281320
rect 289 281040 352640 281176
rect 289 280640 353451 281040
rect 880 280360 353451 280640
rect 289 280232 353451 280360
rect 289 279960 352640 280232
rect 880 279952 352640 279960
rect 880 279680 353451 279952
rect 289 279280 353451 279680
rect 880 279144 353451 279280
rect 880 279000 352640 279144
rect 289 278864 352640 279000
rect 289 278600 353451 278864
rect 880 278320 353451 278600
rect 289 278056 353451 278320
rect 289 277920 352640 278056
rect 880 277776 352640 277920
rect 880 277640 353451 277776
rect 289 277240 353451 277640
rect 880 277104 353451 277240
rect 880 276960 352640 277104
rect 289 276824 352640 276960
rect 289 276424 353451 276824
rect 880 276144 353451 276424
rect 289 276016 353451 276144
rect 289 275744 352640 276016
rect 880 275736 352640 275744
rect 880 275464 353451 275736
rect 289 275064 353451 275464
rect 880 274928 353451 275064
rect 880 274784 352640 274928
rect 289 274648 352640 274784
rect 289 274384 353451 274648
rect 880 274104 353451 274384
rect 289 273840 353451 274104
rect 289 273704 352640 273840
rect 880 273560 352640 273704
rect 880 273424 353451 273560
rect 289 272888 353451 273424
rect 880 272752 353451 272888
rect 880 272608 352640 272752
rect 289 272472 352640 272608
rect 289 272208 353451 272472
rect 880 271928 353451 272208
rect 289 271664 353451 271928
rect 289 271528 352640 271664
rect 880 271384 352640 271528
rect 880 271248 353451 271384
rect 289 270848 353451 271248
rect 880 270576 353451 270848
rect 880 270568 352640 270576
rect 289 270296 352640 270568
rect 289 270168 353451 270296
rect 880 269888 353451 270168
rect 289 269488 353451 269888
rect 880 269208 352640 269488
rect 289 268672 353451 269208
rect 880 268400 353451 268672
rect 880 268392 352640 268400
rect 289 268120 352640 268392
rect 289 267992 353451 268120
rect 880 267712 353451 267992
rect 289 267312 353451 267712
rect 880 267032 352640 267312
rect 289 266632 353451 267032
rect 880 266352 353451 266632
rect 289 266224 353451 266352
rect 289 265952 352640 266224
rect 880 265944 352640 265952
rect 880 265672 353451 265944
rect 289 265272 353451 265672
rect 880 265136 353451 265272
rect 880 264992 352640 265136
rect 289 264856 352640 264992
rect 289 264456 353451 264856
rect 880 264176 353451 264456
rect 289 264048 353451 264176
rect 289 263776 352640 264048
rect 880 263768 352640 263776
rect 880 263496 353451 263768
rect 289 263096 353451 263496
rect 880 262960 353451 263096
rect 880 262816 352640 262960
rect 289 262680 352640 262816
rect 289 262416 353451 262680
rect 880 262136 353451 262416
rect 289 261872 353451 262136
rect 289 261736 352640 261872
rect 880 261592 352640 261736
rect 880 261456 353451 261592
rect 289 260920 353451 261456
rect 880 260784 353451 260920
rect 880 260640 352640 260784
rect 289 260504 352640 260640
rect 289 260240 353451 260504
rect 880 259960 353451 260240
rect 289 259696 353451 259960
rect 289 259560 352640 259696
rect 880 259416 352640 259560
rect 880 259280 353451 259416
rect 289 258880 353451 259280
rect 880 258608 353451 258880
rect 880 258600 352640 258608
rect 289 258328 352640 258600
rect 289 258200 353451 258328
rect 880 257920 353451 258200
rect 289 257520 353451 257920
rect 880 257240 352640 257520
rect 289 256704 353451 257240
rect 880 256432 353451 256704
rect 880 256424 352640 256432
rect 289 256152 352640 256424
rect 289 256024 353451 256152
rect 880 255744 353451 256024
rect 289 255344 353451 255744
rect 880 255064 352640 255344
rect 289 254664 353451 255064
rect 880 254384 353451 254664
rect 289 254256 353451 254384
rect 289 253984 352640 254256
rect 880 253976 352640 253984
rect 880 253704 353451 253976
rect 289 253168 353451 253704
rect 880 252888 352640 253168
rect 289 252488 353451 252888
rect 880 252208 353451 252488
rect 289 252080 353451 252208
rect 289 251808 352640 252080
rect 880 251800 352640 251808
rect 880 251528 353451 251800
rect 289 251128 353451 251528
rect 880 250992 353451 251128
rect 880 250848 352640 250992
rect 289 250712 352640 250848
rect 289 250448 353451 250712
rect 880 250168 353451 250448
rect 289 249904 353451 250168
rect 289 249768 352640 249904
rect 880 249624 352640 249768
rect 880 249488 353451 249624
rect 289 248952 353451 249488
rect 880 248816 353451 248952
rect 880 248672 352640 248816
rect 289 248536 352640 248672
rect 289 248272 353451 248536
rect 880 247992 353451 248272
rect 289 247728 353451 247992
rect 289 247592 352640 247728
rect 880 247448 352640 247592
rect 880 247312 353451 247448
rect 289 246912 353451 247312
rect 880 246640 353451 246912
rect 880 246632 352640 246640
rect 289 246360 352640 246632
rect 289 246232 353451 246360
rect 880 245952 353451 246232
rect 289 245552 353451 245952
rect 880 245272 352640 245552
rect 289 244736 353451 245272
rect 880 244464 353451 244736
rect 880 244456 352640 244464
rect 289 244184 352640 244456
rect 289 244056 353451 244184
rect 880 243776 353451 244056
rect 289 243376 353451 243776
rect 880 243096 352640 243376
rect 289 242696 353451 243096
rect 880 242416 353451 242696
rect 289 242288 353451 242416
rect 289 242016 352640 242288
rect 880 242008 352640 242016
rect 880 241736 353451 242008
rect 289 241200 353451 241736
rect 880 240920 352640 241200
rect 289 240520 353451 240920
rect 880 240240 353451 240520
rect 289 240112 353451 240240
rect 289 239840 352640 240112
rect 880 239832 352640 239840
rect 880 239560 353451 239832
rect 289 239160 353451 239560
rect 880 239024 353451 239160
rect 880 238880 352640 239024
rect 289 238744 352640 238880
rect 289 238480 353451 238744
rect 880 238200 353451 238480
rect 289 237936 353451 238200
rect 289 237800 352640 237936
rect 880 237656 352640 237800
rect 880 237520 353451 237656
rect 289 236984 353451 237520
rect 880 236704 352640 236984
rect 289 236304 353451 236704
rect 880 236024 353451 236304
rect 289 235896 353451 236024
rect 289 235624 352640 235896
rect 880 235616 352640 235624
rect 880 235344 353451 235616
rect 289 234944 353451 235344
rect 880 234808 353451 234944
rect 880 234664 352640 234808
rect 289 234528 352640 234664
rect 289 234264 353451 234528
rect 880 233984 353451 234264
rect 289 233720 353451 233984
rect 289 233448 352640 233720
rect 880 233440 352640 233448
rect 880 233168 353451 233440
rect 289 232768 353451 233168
rect 880 232632 353451 232768
rect 880 232488 352640 232632
rect 289 232352 352640 232488
rect 289 232088 353451 232352
rect 880 231808 353451 232088
rect 289 231544 353451 231808
rect 289 231408 352640 231544
rect 880 231264 352640 231408
rect 880 231128 353451 231264
rect 289 230728 353451 231128
rect 880 230456 353451 230728
rect 880 230448 352640 230456
rect 289 230176 352640 230448
rect 289 230048 353451 230176
rect 880 229768 353451 230048
rect 289 229368 353451 229768
rect 289 229232 352640 229368
rect 880 229088 352640 229232
rect 880 228952 353451 229088
rect 289 228552 353451 228952
rect 880 228280 353451 228552
rect 880 228272 352640 228280
rect 289 228000 352640 228272
rect 289 227872 353451 228000
rect 880 227592 353451 227872
rect 289 227192 353451 227592
rect 880 226912 352640 227192
rect 289 226512 353451 226912
rect 880 226232 353451 226512
rect 289 226104 353451 226232
rect 289 225832 352640 226104
rect 880 225824 352640 225832
rect 880 225552 353451 225824
rect 289 225016 353451 225552
rect 880 224736 352640 225016
rect 289 224336 353451 224736
rect 880 224056 353451 224336
rect 289 223928 353451 224056
rect 289 223656 352640 223928
rect 880 223648 352640 223656
rect 880 223376 353451 223648
rect 289 222976 353451 223376
rect 880 222840 353451 222976
rect 880 222696 352640 222840
rect 289 222560 352640 222696
rect 289 222296 353451 222560
rect 880 222016 353451 222296
rect 289 221752 353451 222016
rect 289 221480 352640 221752
rect 880 221472 352640 221480
rect 880 221200 353451 221472
rect 289 220800 353451 221200
rect 880 220664 353451 220800
rect 880 220520 352640 220664
rect 289 220384 352640 220520
rect 289 220120 353451 220384
rect 880 219840 353451 220120
rect 289 219576 353451 219840
rect 289 219440 352640 219576
rect 880 219296 352640 219440
rect 880 219160 353451 219296
rect 289 218760 353451 219160
rect 880 218488 353451 218760
rect 880 218480 352640 218488
rect 289 218208 352640 218480
rect 289 218080 353451 218208
rect 880 217800 353451 218080
rect 289 217400 353451 217800
rect 289 217264 352640 217400
rect 880 217120 352640 217264
rect 880 216984 353451 217120
rect 289 216584 353451 216984
rect 880 216312 353451 216584
rect 880 216304 352640 216312
rect 289 216032 352640 216304
rect 289 215904 353451 216032
rect 880 215624 353451 215904
rect 289 215224 353451 215624
rect 880 214944 352640 215224
rect 289 214544 353451 214944
rect 880 214264 353451 214544
rect 289 214136 353451 214264
rect 289 213864 352640 214136
rect 880 213856 352640 213864
rect 880 213584 353451 213856
rect 289 213048 353451 213584
rect 880 212768 352640 213048
rect 289 212368 353451 212768
rect 880 212088 353451 212368
rect 289 211960 353451 212088
rect 289 211688 352640 211960
rect 880 211680 352640 211688
rect 880 211408 353451 211680
rect 289 211008 353451 211408
rect 880 210872 353451 211008
rect 880 210728 352640 210872
rect 289 210592 352640 210728
rect 289 210328 353451 210592
rect 880 210048 353451 210328
rect 289 209784 353451 210048
rect 289 209512 352640 209784
rect 880 209504 352640 209512
rect 880 209232 353451 209504
rect 289 208832 353451 209232
rect 880 208696 353451 208832
rect 880 208552 352640 208696
rect 289 208416 352640 208552
rect 289 208152 353451 208416
rect 880 207872 353451 208152
rect 289 207608 353451 207872
rect 289 207472 352640 207608
rect 880 207328 352640 207472
rect 880 207192 353451 207328
rect 289 206792 353451 207192
rect 880 206520 353451 206792
rect 880 206512 352640 206520
rect 289 206240 352640 206512
rect 289 206112 353451 206240
rect 880 205832 353451 206112
rect 289 205432 353451 205832
rect 289 205296 352640 205432
rect 880 205152 352640 205296
rect 880 205016 353451 205152
rect 289 204616 353451 205016
rect 880 204344 353451 204616
rect 880 204336 352640 204344
rect 289 204064 352640 204336
rect 289 203936 353451 204064
rect 880 203656 353451 203936
rect 289 203256 353451 203656
rect 880 202976 352640 203256
rect 289 202576 353451 202976
rect 880 202296 353451 202576
rect 289 202168 353451 202296
rect 289 201888 352640 202168
rect 289 201760 353451 201888
rect 880 201480 353451 201760
rect 289 201080 353451 201480
rect 880 200800 352640 201080
rect 289 200400 353451 200800
rect 880 200120 353451 200400
rect 289 199992 353451 200120
rect 289 199720 352640 199992
rect 880 199712 352640 199720
rect 880 199440 353451 199712
rect 289 199040 353451 199440
rect 880 198904 353451 199040
rect 880 198760 352640 198904
rect 289 198624 352640 198760
rect 289 198360 353451 198624
rect 880 198080 353451 198360
rect 289 197952 353451 198080
rect 289 197672 352640 197952
rect 289 197544 353451 197672
rect 880 197264 353451 197544
rect 289 196864 353451 197264
rect 880 196584 352640 196864
rect 289 196184 353451 196584
rect 880 195904 353451 196184
rect 289 195776 353451 195904
rect 289 195504 352640 195776
rect 880 195496 352640 195504
rect 880 195224 353451 195496
rect 289 194824 353451 195224
rect 880 194688 353451 194824
rect 880 194544 352640 194688
rect 289 194408 352640 194544
rect 289 194144 353451 194408
rect 880 193864 353451 194144
rect 289 193600 353451 193864
rect 289 193328 352640 193600
rect 880 193320 352640 193328
rect 880 193048 353451 193320
rect 289 192648 353451 193048
rect 880 192512 353451 192648
rect 880 192368 352640 192512
rect 289 192232 352640 192368
rect 289 191968 353451 192232
rect 880 191688 353451 191968
rect 289 191424 353451 191688
rect 289 191288 352640 191424
rect 880 191144 352640 191288
rect 880 191008 353451 191144
rect 289 190608 353451 191008
rect 880 190336 353451 190608
rect 880 190328 352640 190336
rect 289 190056 352640 190328
rect 289 189792 353451 190056
rect 880 189512 353451 189792
rect 289 189248 353451 189512
rect 289 189112 352640 189248
rect 880 188968 352640 189112
rect 880 188832 353451 188968
rect 289 188432 353451 188832
rect 880 188160 353451 188432
rect 880 188152 352640 188160
rect 289 187880 352640 188152
rect 289 187752 353451 187880
rect 880 187472 353451 187752
rect 289 187072 353451 187472
rect 880 186792 352640 187072
rect 289 186392 353451 186792
rect 880 186112 353451 186392
rect 289 185984 353451 186112
rect 289 185704 352640 185984
rect 289 185576 353451 185704
rect 880 185296 353451 185576
rect 289 184896 353451 185296
rect 880 184616 352640 184896
rect 289 184216 353451 184616
rect 880 183936 353451 184216
rect 289 183808 353451 183936
rect 289 183536 352640 183808
rect 880 183528 352640 183536
rect 880 183256 353451 183528
rect 289 182856 353451 183256
rect 880 182720 353451 182856
rect 880 182576 352640 182720
rect 289 182440 352640 182576
rect 289 182040 353451 182440
rect 880 181760 353451 182040
rect 289 181632 353451 181760
rect 289 181360 352640 181632
rect 880 181352 352640 181360
rect 880 181080 353451 181352
rect 289 180680 353451 181080
rect 880 180544 353451 180680
rect 880 180400 352640 180544
rect 289 180264 352640 180400
rect 289 180000 353451 180264
rect 880 179720 353451 180000
rect 289 179456 353451 179720
rect 289 179320 352640 179456
rect 880 179176 352640 179320
rect 880 179040 353451 179176
rect 289 178640 353451 179040
rect 880 178368 353451 178640
rect 880 178360 352640 178368
rect 289 178088 352640 178360
rect 289 177824 353451 178088
rect 880 177544 353451 177824
rect 289 177280 353451 177544
rect 289 177144 352640 177280
rect 880 177000 352640 177144
rect 880 176864 353451 177000
rect 289 176464 353451 176864
rect 880 176192 353451 176464
rect 880 176184 352640 176192
rect 289 175912 352640 176184
rect 289 175784 353451 175912
rect 880 175504 353451 175784
rect 289 175104 353451 175504
rect 880 174824 352640 175104
rect 289 174424 353451 174824
rect 880 174144 353451 174424
rect 289 174016 353451 174144
rect 289 173736 352640 174016
rect 289 173608 353451 173736
rect 880 173328 353451 173608
rect 289 172928 353451 173328
rect 880 172648 352640 172928
rect 289 172248 353451 172648
rect 880 171968 353451 172248
rect 289 171840 353451 171968
rect 289 171568 352640 171840
rect 880 171560 352640 171568
rect 880 171288 353451 171560
rect 289 170888 353451 171288
rect 880 170752 353451 170888
rect 880 170608 352640 170752
rect 289 170472 352640 170608
rect 289 170072 353451 170472
rect 880 169792 353451 170072
rect 289 169664 353451 169792
rect 289 169392 352640 169664
rect 880 169384 352640 169392
rect 880 169112 353451 169384
rect 289 168712 353451 169112
rect 880 168576 353451 168712
rect 880 168432 352640 168576
rect 289 168296 352640 168432
rect 289 168032 353451 168296
rect 880 167752 353451 168032
rect 289 167488 353451 167752
rect 289 167352 352640 167488
rect 880 167208 352640 167352
rect 880 167072 353451 167208
rect 289 166672 353451 167072
rect 880 166400 353451 166672
rect 880 166392 352640 166400
rect 289 166120 352640 166392
rect 289 165856 353451 166120
rect 880 165576 353451 165856
rect 289 165312 353451 165576
rect 289 165176 352640 165312
rect 880 165032 352640 165176
rect 880 164896 353451 165032
rect 289 164496 353451 164896
rect 880 164224 353451 164496
rect 880 164216 352640 164224
rect 289 163944 352640 164216
rect 289 163816 353451 163944
rect 880 163536 353451 163816
rect 289 163136 353451 163536
rect 880 162856 352640 163136
rect 289 162320 353451 162856
rect 880 162048 353451 162320
rect 880 162040 352640 162048
rect 289 161768 352640 162040
rect 289 161640 353451 161768
rect 880 161360 353451 161640
rect 289 160960 353451 161360
rect 880 160680 352640 160960
rect 289 160280 353451 160680
rect 880 160000 353451 160280
rect 289 159872 353451 160000
rect 289 159600 352640 159872
rect 880 159592 352640 159600
rect 880 159320 353451 159592
rect 289 158920 353451 159320
rect 880 158784 353451 158920
rect 880 158640 352640 158784
rect 289 158504 352640 158640
rect 289 158104 353451 158504
rect 880 157832 353451 158104
rect 880 157824 352640 157832
rect 289 157552 352640 157824
rect 289 157424 353451 157552
rect 880 157144 353451 157424
rect 289 156744 353451 157144
rect 880 156464 352640 156744
rect 289 156064 353451 156464
rect 880 155784 353451 156064
rect 289 155656 353451 155784
rect 289 155384 352640 155656
rect 880 155376 352640 155384
rect 880 155104 353451 155376
rect 289 154704 353451 155104
rect 880 154568 353451 154704
rect 880 154424 352640 154568
rect 289 154288 352640 154424
rect 289 153888 353451 154288
rect 880 153608 353451 153888
rect 289 153480 353451 153608
rect 289 153208 352640 153480
rect 880 153200 352640 153208
rect 880 152928 353451 153200
rect 289 152528 353451 152928
rect 880 152392 353451 152528
rect 880 152248 352640 152392
rect 289 152112 352640 152248
rect 289 151848 353451 152112
rect 880 151568 353451 151848
rect 289 151304 353451 151568
rect 289 151168 352640 151304
rect 880 151024 352640 151168
rect 880 150888 353451 151024
rect 289 150352 353451 150888
rect 880 150216 353451 150352
rect 880 150072 352640 150216
rect 289 149936 352640 150072
rect 289 149672 353451 149936
rect 880 149392 353451 149672
rect 289 149128 353451 149392
rect 289 148992 352640 149128
rect 880 148848 352640 148992
rect 880 148712 353451 148848
rect 289 148312 353451 148712
rect 880 148040 353451 148312
rect 880 148032 352640 148040
rect 289 147760 352640 148032
rect 289 147632 353451 147760
rect 880 147352 353451 147632
rect 289 146952 353451 147352
rect 880 146672 352640 146952
rect 289 146136 353451 146672
rect 880 145864 353451 146136
rect 880 145856 352640 145864
rect 289 145584 352640 145856
rect 289 145456 353451 145584
rect 880 145176 353451 145456
rect 289 144776 353451 145176
rect 880 144496 352640 144776
rect 289 144096 353451 144496
rect 880 143816 353451 144096
rect 289 143688 353451 143816
rect 289 143416 352640 143688
rect 880 143408 352640 143416
rect 880 143136 353451 143408
rect 289 142736 353451 143136
rect 880 142600 353451 142736
rect 880 142456 352640 142600
rect 289 142320 352640 142456
rect 289 141920 353451 142320
rect 880 141640 353451 141920
rect 289 141512 353451 141640
rect 289 141240 352640 141512
rect 880 141232 352640 141240
rect 880 140960 353451 141232
rect 289 140560 353451 140960
rect 880 140424 353451 140560
rect 880 140280 352640 140424
rect 289 140144 352640 140280
rect 289 139880 353451 140144
rect 880 139600 353451 139880
rect 289 139336 353451 139600
rect 289 139200 352640 139336
rect 880 139056 352640 139200
rect 880 138920 353451 139056
rect 289 138384 353451 138920
rect 880 138248 353451 138384
rect 880 138104 352640 138248
rect 289 137968 352640 138104
rect 289 137704 353451 137968
rect 880 137424 353451 137704
rect 289 137160 353451 137424
rect 289 137024 352640 137160
rect 880 136880 352640 137024
rect 880 136744 353451 136880
rect 289 136344 353451 136744
rect 880 136072 353451 136344
rect 880 136064 352640 136072
rect 289 135792 352640 136064
rect 289 135664 353451 135792
rect 880 135384 353451 135664
rect 289 134984 353451 135384
rect 880 134704 352640 134984
rect 289 134168 353451 134704
rect 880 133896 353451 134168
rect 880 133888 352640 133896
rect 289 133616 352640 133888
rect 289 133488 353451 133616
rect 880 133208 353451 133488
rect 289 132808 353451 133208
rect 880 132528 352640 132808
rect 289 132128 353451 132528
rect 880 131848 353451 132128
rect 289 131720 353451 131848
rect 289 131448 352640 131720
rect 880 131440 352640 131448
rect 880 131168 353451 131440
rect 289 130632 353451 131168
rect 880 130352 352640 130632
rect 289 129952 353451 130352
rect 880 129672 353451 129952
rect 289 129544 353451 129672
rect 289 129272 352640 129544
rect 880 129264 352640 129272
rect 880 128992 353451 129264
rect 289 128592 353451 128992
rect 880 128456 353451 128592
rect 880 128312 352640 128456
rect 289 128176 352640 128312
rect 289 127912 353451 128176
rect 880 127632 353451 127912
rect 289 127368 353451 127632
rect 289 127232 352640 127368
rect 880 127088 352640 127232
rect 880 126952 353451 127088
rect 289 126416 353451 126952
rect 880 126280 353451 126416
rect 880 126136 352640 126280
rect 289 126000 352640 126136
rect 289 125736 353451 126000
rect 880 125456 353451 125736
rect 289 125192 353451 125456
rect 289 125056 352640 125192
rect 880 124912 352640 125056
rect 880 124776 353451 124912
rect 289 124376 353451 124776
rect 880 124104 353451 124376
rect 880 124096 352640 124104
rect 289 123824 352640 124096
rect 289 123696 353451 123824
rect 880 123416 353451 123696
rect 289 123016 353451 123416
rect 880 122736 352640 123016
rect 289 122200 353451 122736
rect 880 121928 353451 122200
rect 880 121920 352640 121928
rect 289 121648 352640 121920
rect 289 121520 353451 121648
rect 880 121240 353451 121520
rect 289 120840 353451 121240
rect 880 120560 352640 120840
rect 289 120160 353451 120560
rect 880 119880 353451 120160
rect 289 119752 353451 119880
rect 289 119480 352640 119752
rect 880 119472 352640 119480
rect 880 119200 353451 119472
rect 289 118800 353451 119200
rect 289 118664 352640 118800
rect 880 118520 352640 118664
rect 880 118384 353451 118520
rect 289 117984 353451 118384
rect 880 117712 353451 117984
rect 880 117704 352640 117712
rect 289 117432 352640 117704
rect 289 117304 353451 117432
rect 880 117024 353451 117304
rect 289 116624 353451 117024
rect 880 116344 352640 116624
rect 289 115944 353451 116344
rect 880 115664 353451 115944
rect 289 115536 353451 115664
rect 289 115264 352640 115536
rect 880 115256 352640 115264
rect 880 114984 353451 115256
rect 289 114448 353451 114984
rect 880 114168 352640 114448
rect 289 113768 353451 114168
rect 880 113488 353451 113768
rect 289 113360 353451 113488
rect 289 113088 352640 113360
rect 880 113080 352640 113088
rect 880 112808 353451 113080
rect 289 112408 353451 112808
rect 880 112272 353451 112408
rect 880 112128 352640 112272
rect 289 111992 352640 112128
rect 289 111728 353451 111992
rect 880 111448 353451 111728
rect 289 111184 353451 111448
rect 289 110912 352640 111184
rect 880 110904 352640 110912
rect 880 110632 353451 110904
rect 289 110232 353451 110632
rect 880 110096 353451 110232
rect 880 109952 352640 110096
rect 289 109816 352640 109952
rect 289 109552 353451 109816
rect 880 109272 353451 109552
rect 289 109008 353451 109272
rect 289 108872 352640 109008
rect 880 108728 352640 108872
rect 880 108592 353451 108728
rect 289 108192 353451 108592
rect 880 107920 353451 108192
rect 880 107912 352640 107920
rect 289 107640 352640 107912
rect 289 107512 353451 107640
rect 880 107232 353451 107512
rect 289 106832 353451 107232
rect 289 106696 352640 106832
rect 880 106552 352640 106696
rect 880 106416 353451 106552
rect 289 106016 353451 106416
rect 880 105744 353451 106016
rect 880 105736 352640 105744
rect 289 105464 352640 105736
rect 289 105336 353451 105464
rect 880 105056 353451 105336
rect 289 104656 353451 105056
rect 880 104376 352640 104656
rect 289 103976 353451 104376
rect 880 103696 353451 103976
rect 289 103568 353451 103696
rect 289 103296 352640 103568
rect 880 103288 352640 103296
rect 880 103016 353451 103288
rect 289 102480 353451 103016
rect 880 102200 352640 102480
rect 289 101800 353451 102200
rect 880 101520 353451 101800
rect 289 101392 353451 101520
rect 289 101120 352640 101392
rect 880 101112 352640 101120
rect 880 100840 353451 101112
rect 289 100440 353451 100840
rect 880 100304 353451 100440
rect 880 100160 352640 100304
rect 289 100024 352640 100160
rect 289 99760 353451 100024
rect 880 99480 353451 99760
rect 289 99216 353451 99480
rect 289 98944 352640 99216
rect 880 98936 352640 98944
rect 880 98664 353451 98936
rect 289 98264 353451 98664
rect 880 98128 353451 98264
rect 880 97984 352640 98128
rect 289 97848 352640 97984
rect 289 97584 353451 97848
rect 880 97304 353451 97584
rect 289 97040 353451 97304
rect 289 96904 352640 97040
rect 880 96760 352640 96904
rect 880 96624 353451 96760
rect 289 96224 353451 96624
rect 880 95952 353451 96224
rect 880 95944 352640 95952
rect 289 95672 352640 95944
rect 289 95544 353451 95672
rect 880 95264 353451 95544
rect 289 94864 353451 95264
rect 289 94728 352640 94864
rect 880 94584 352640 94728
rect 880 94448 353451 94584
rect 289 94048 353451 94448
rect 880 93776 353451 94048
rect 880 93768 352640 93776
rect 289 93496 352640 93768
rect 289 93368 353451 93496
rect 880 93088 353451 93368
rect 289 92688 353451 93088
rect 880 92408 352640 92688
rect 289 92008 353451 92408
rect 880 91728 353451 92008
rect 289 91600 353451 91728
rect 289 91320 352640 91600
rect 289 91192 353451 91320
rect 880 90912 353451 91192
rect 289 90512 353451 90912
rect 880 90232 352640 90512
rect 289 89832 353451 90232
rect 880 89552 353451 89832
rect 289 89424 353451 89552
rect 289 89152 352640 89424
rect 880 89144 352640 89152
rect 880 88872 353451 89144
rect 289 88472 353451 88872
rect 880 88336 353451 88472
rect 880 88192 352640 88336
rect 289 88056 352640 88192
rect 289 87792 353451 88056
rect 880 87512 353451 87792
rect 289 87248 353451 87512
rect 289 86976 352640 87248
rect 880 86968 352640 86976
rect 880 86696 353451 86968
rect 289 86296 353451 86696
rect 880 86160 353451 86296
rect 880 86016 352640 86160
rect 289 85880 352640 86016
rect 289 85616 353451 85880
rect 880 85336 353451 85616
rect 289 85072 353451 85336
rect 289 84936 352640 85072
rect 880 84792 352640 84936
rect 880 84656 353451 84792
rect 289 84256 353451 84656
rect 880 83984 353451 84256
rect 880 83976 352640 83984
rect 289 83704 352640 83976
rect 289 83576 353451 83704
rect 880 83296 353451 83576
rect 289 82896 353451 83296
rect 289 82760 352640 82896
rect 880 82616 352640 82760
rect 880 82480 353451 82616
rect 289 82080 353451 82480
rect 880 81808 353451 82080
rect 880 81800 352640 81808
rect 289 81528 352640 81800
rect 289 81400 353451 81528
rect 880 81120 353451 81400
rect 289 80720 353451 81120
rect 880 80440 352640 80720
rect 289 80040 353451 80440
rect 880 79760 353451 80040
rect 289 79632 353451 79760
rect 289 79352 352640 79632
rect 289 79224 353451 79352
rect 880 78944 353451 79224
rect 289 78680 353451 78944
rect 289 78544 352640 78680
rect 880 78400 352640 78544
rect 880 78264 353451 78400
rect 289 77864 353451 78264
rect 880 77592 353451 77864
rect 880 77584 352640 77592
rect 289 77312 352640 77584
rect 289 77184 353451 77312
rect 880 76904 353451 77184
rect 289 76504 353451 76904
rect 880 76224 352640 76504
rect 289 75824 353451 76224
rect 880 75544 353451 75824
rect 289 75416 353451 75544
rect 289 75136 352640 75416
rect 289 75008 353451 75136
rect 880 74728 353451 75008
rect 289 74328 353451 74728
rect 880 74048 352640 74328
rect 289 73648 353451 74048
rect 880 73368 353451 73648
rect 289 73240 353451 73368
rect 289 72968 352640 73240
rect 880 72960 352640 72968
rect 880 72688 353451 72960
rect 289 72288 353451 72688
rect 880 72152 353451 72288
rect 880 72008 352640 72152
rect 289 71872 352640 72008
rect 289 71608 353451 71872
rect 880 71328 353451 71608
rect 289 71064 353451 71328
rect 289 70792 352640 71064
rect 880 70784 352640 70792
rect 880 70512 353451 70784
rect 289 70112 353451 70512
rect 880 69976 353451 70112
rect 880 69832 352640 69976
rect 289 69696 352640 69832
rect 289 69432 353451 69696
rect 880 69152 353451 69432
rect 289 68888 353451 69152
rect 289 68752 352640 68888
rect 880 68608 352640 68752
rect 880 68472 353451 68608
rect 289 68072 353451 68472
rect 880 67800 353451 68072
rect 880 67792 352640 67800
rect 289 67520 352640 67792
rect 289 67256 353451 67520
rect 880 66976 353451 67256
rect 289 66712 353451 66976
rect 289 66576 352640 66712
rect 880 66432 352640 66576
rect 880 66296 353451 66432
rect 289 65896 353451 66296
rect 880 65624 353451 65896
rect 880 65616 352640 65624
rect 289 65344 352640 65616
rect 289 65216 353451 65344
rect 880 64936 353451 65216
rect 289 64536 353451 64936
rect 880 64256 352640 64536
rect 289 63856 353451 64256
rect 880 63576 353451 63856
rect 289 63448 353451 63576
rect 289 63168 352640 63448
rect 289 63040 353451 63168
rect 880 62760 353451 63040
rect 289 62360 353451 62760
rect 880 62080 352640 62360
rect 289 61680 353451 62080
rect 880 61400 353451 61680
rect 289 61272 353451 61400
rect 289 61000 352640 61272
rect 880 60992 352640 61000
rect 880 60720 353451 60992
rect 289 60320 353451 60720
rect 880 60184 353451 60320
rect 880 60040 352640 60184
rect 289 59904 352640 60040
rect 289 59504 353451 59904
rect 880 59224 353451 59504
rect 289 59096 353451 59224
rect 289 58824 352640 59096
rect 880 58816 352640 58824
rect 880 58544 353451 58816
rect 289 58144 353451 58544
rect 880 58008 353451 58144
rect 880 57864 352640 58008
rect 289 57728 352640 57864
rect 289 57464 353451 57728
rect 880 57184 353451 57464
rect 289 56920 353451 57184
rect 289 56784 352640 56920
rect 880 56640 352640 56784
rect 880 56504 353451 56640
rect 289 56104 353451 56504
rect 880 55832 353451 56104
rect 880 55824 352640 55832
rect 289 55552 352640 55824
rect 289 55288 353451 55552
rect 880 55008 353451 55288
rect 289 54744 353451 55008
rect 289 54608 352640 54744
rect 880 54464 352640 54608
rect 880 54328 353451 54464
rect 289 53928 353451 54328
rect 880 53656 353451 53928
rect 880 53648 352640 53656
rect 289 53376 352640 53648
rect 289 53248 353451 53376
rect 880 52968 353451 53248
rect 289 52568 353451 52968
rect 880 52288 352640 52568
rect 289 51888 353451 52288
rect 880 51608 353451 51888
rect 289 51480 353451 51608
rect 289 51200 352640 51480
rect 289 51072 353451 51200
rect 880 50792 353451 51072
rect 289 50392 353451 50792
rect 880 50112 352640 50392
rect 289 49712 353451 50112
rect 880 49432 353451 49712
rect 289 49304 353451 49432
rect 289 49032 352640 49304
rect 880 49024 352640 49032
rect 880 48752 353451 49024
rect 289 48352 353451 48752
rect 880 48216 353451 48352
rect 880 48072 352640 48216
rect 289 47936 352640 48072
rect 289 47536 353451 47936
rect 880 47256 353451 47536
rect 289 47128 353451 47256
rect 289 46856 352640 47128
rect 880 46848 352640 46856
rect 880 46576 353451 46848
rect 289 46176 353451 46576
rect 880 46040 353451 46176
rect 880 45896 352640 46040
rect 289 45760 352640 45896
rect 289 45496 353451 45760
rect 880 45216 353451 45496
rect 289 44952 353451 45216
rect 289 44816 352640 44952
rect 880 44672 352640 44816
rect 880 44536 353451 44672
rect 289 44136 353451 44536
rect 880 43864 353451 44136
rect 880 43856 352640 43864
rect 289 43584 352640 43856
rect 289 43320 353451 43584
rect 880 43040 353451 43320
rect 289 42776 353451 43040
rect 289 42640 352640 42776
rect 880 42496 352640 42640
rect 880 42360 353451 42496
rect 289 41960 353451 42360
rect 880 41688 353451 41960
rect 880 41680 352640 41688
rect 289 41408 352640 41680
rect 289 41280 353451 41408
rect 880 41000 353451 41280
rect 289 40600 353451 41000
rect 880 40320 352640 40600
rect 289 39784 353451 40320
rect 880 39648 353451 39784
rect 880 39504 352640 39648
rect 289 39368 352640 39504
rect 289 39104 353451 39368
rect 880 38824 353451 39104
rect 289 38560 353451 38824
rect 289 38424 352640 38560
rect 880 38280 352640 38424
rect 880 38144 353451 38280
rect 289 37744 353451 38144
rect 880 37472 353451 37744
rect 880 37464 352640 37472
rect 289 37192 352640 37464
rect 289 37064 353451 37192
rect 880 36784 353451 37064
rect 289 36384 353451 36784
rect 880 36104 352640 36384
rect 289 35568 353451 36104
rect 880 35296 353451 35568
rect 880 35288 352640 35296
rect 289 35016 352640 35288
rect 289 34888 353451 35016
rect 880 34608 353451 34888
rect 289 34208 353451 34608
rect 880 33928 352640 34208
rect 289 33528 353451 33928
rect 880 33248 353451 33528
rect 289 33120 353451 33248
rect 289 32848 352640 33120
rect 880 32840 352640 32848
rect 880 32568 353451 32840
rect 289 32168 353451 32568
rect 880 32032 353451 32168
rect 880 31888 352640 32032
rect 289 31752 352640 31888
rect 289 31352 353451 31752
rect 880 31072 353451 31352
rect 289 30944 353451 31072
rect 289 30672 352640 30944
rect 880 30664 352640 30672
rect 880 30392 353451 30664
rect 289 29992 353451 30392
rect 880 29856 353451 29992
rect 880 29712 352640 29856
rect 289 29576 352640 29712
rect 289 29312 353451 29576
rect 880 29032 353451 29312
rect 289 28768 353451 29032
rect 289 28632 352640 28768
rect 880 28488 352640 28632
rect 880 28352 353451 28488
rect 289 27816 353451 28352
rect 880 27680 353451 27816
rect 880 27536 352640 27680
rect 289 27400 352640 27536
rect 289 27136 353451 27400
rect 880 26856 353451 27136
rect 289 26592 353451 26856
rect 289 26456 352640 26592
rect 880 26312 352640 26456
rect 880 26176 353451 26312
rect 289 25776 353451 26176
rect 880 25504 353451 25776
rect 880 25496 352640 25504
rect 289 25224 352640 25496
rect 289 25096 353451 25224
rect 880 24816 353451 25096
rect 289 24416 353451 24816
rect 880 24136 352640 24416
rect 289 23600 353451 24136
rect 880 23328 353451 23600
rect 880 23320 352640 23328
rect 289 23048 352640 23320
rect 289 22920 353451 23048
rect 880 22640 353451 22920
rect 289 22240 353451 22640
rect 880 21960 352640 22240
rect 289 21560 353451 21960
rect 880 21280 353451 21560
rect 289 21152 353451 21280
rect 289 20880 352640 21152
rect 880 20872 352640 20880
rect 880 20600 353451 20872
rect 289 20064 353451 20600
rect 880 19784 352640 20064
rect 289 19384 353451 19784
rect 880 19104 353451 19384
rect 289 18976 353451 19104
rect 289 18704 352640 18976
rect 880 18696 352640 18704
rect 880 18424 353451 18696
rect 289 18024 353451 18424
rect 880 17888 353451 18024
rect 880 17744 352640 17888
rect 289 17608 352640 17744
rect 289 17344 353451 17608
rect 880 17064 353451 17344
rect 289 16800 353451 17064
rect 289 16664 352640 16800
rect 880 16520 352640 16664
rect 880 16384 353451 16520
rect 289 15848 353451 16384
rect 880 15712 353451 15848
rect 880 15568 352640 15712
rect 289 15432 352640 15568
rect 289 15168 353451 15432
rect 880 14888 353451 15168
rect 289 14624 353451 14888
rect 289 14488 352640 14624
rect 880 14344 352640 14488
rect 880 14208 353451 14344
rect 289 13808 353451 14208
rect 880 13536 353451 13808
rect 880 13528 352640 13536
rect 289 13256 352640 13528
rect 289 13128 353451 13256
rect 880 12848 353451 13128
rect 289 12448 353451 12848
rect 880 12168 352640 12448
rect 289 11632 353451 12168
rect 880 11360 353451 11632
rect 880 11352 352640 11360
rect 289 11080 352640 11352
rect 289 10952 353451 11080
rect 880 10672 353451 10952
rect 289 10272 353451 10672
rect 880 9992 352640 10272
rect 289 9592 353451 9992
rect 880 9312 353451 9592
rect 289 9184 353451 9312
rect 289 8912 352640 9184
rect 880 8904 352640 8912
rect 880 8632 353451 8904
rect 289 8096 353451 8632
rect 880 7816 352640 8096
rect 289 7416 353451 7816
rect 880 7136 353451 7416
rect 289 7008 353451 7136
rect 289 6736 352640 7008
rect 880 6728 352640 6736
rect 880 6456 353451 6728
rect 289 6056 353451 6456
rect 880 5920 353451 6056
rect 880 5776 352640 5920
rect 289 5640 352640 5776
rect 289 5376 353451 5640
rect 880 5096 353451 5376
rect 289 4832 353451 5096
rect 289 4696 352640 4832
rect 880 4552 352640 4696
rect 880 4416 353451 4552
rect 289 3880 353451 4416
rect 880 3744 353451 3880
rect 880 3600 352640 3744
rect 289 3464 352640 3600
rect 289 3200 353451 3464
rect 880 2920 353451 3200
rect 289 2656 353451 2920
rect 289 2520 352640 2656
rect 880 2376 352640 2520
rect 880 2240 353451 2376
rect 289 1840 353451 2240
rect 880 1568 353451 1840
rect 880 1560 352640 1568
rect 289 1288 352640 1560
rect 289 1160 353451 1288
rect 880 880 353451 1160
rect 289 616 353451 880
rect 289 480 352640 616
rect 880 336 352640 480
rect 880 307 353451 336
<< metal4 >>
rect 4208 2128 4528 353104
rect 19568 2128 19888 353104
rect 34928 2128 35248 353104
rect 50288 2128 50608 353104
rect 65648 2128 65968 353104
rect 81008 2128 81328 353104
rect 96368 2128 96688 353104
rect 111728 2128 112048 353104
rect 127088 2128 127408 353104
rect 142448 2128 142768 353104
rect 157808 2128 158128 353104
rect 173168 2128 173488 353104
rect 188528 2128 188848 353104
rect 203888 2128 204208 353104
rect 219248 2128 219568 353104
rect 234608 2128 234928 353104
rect 249968 2128 250288 353104
rect 265328 2128 265648 353104
rect 280688 2128 281008 353104
rect 296048 2128 296368 353104
rect 311408 2128 311728 353104
rect 326768 2128 327088 353104
rect 342128 2128 342448 353104
<< obsm4 >>
rect 795 353184 353405 353565
rect 795 2048 4128 353184
rect 4608 2048 19488 353184
rect 19968 2048 34848 353184
rect 35328 2048 50208 353184
rect 50688 2048 65568 353184
rect 66048 2048 80928 353184
rect 81408 2048 96288 353184
rect 96768 2048 111648 353184
rect 112128 2048 127008 353184
rect 127488 2048 142368 353184
rect 142848 2048 157728 353184
rect 158208 2048 173088 353184
rect 173568 2048 188448 353184
rect 188928 2048 203808 353184
rect 204288 2048 219168 353184
rect 219648 2048 234528 353184
rect 235008 2048 249888 353184
rect 250368 2048 265248 353184
rect 265728 2048 280608 353184
rect 281088 2048 295968 353184
rect 296448 2048 311328 353184
rect 311808 2048 326688 353184
rect 327168 2048 342048 353184
rect 342528 2048 353405 353184
rect 795 1939 353405 2048
<< labels >>
rlabel metal3 s 0 153008 800 153128 6 data_arrays_0_0_ext_ram_addr1[0]
port 1 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 data_arrays_0_0_ext_ram_addr1[1]
port 2 nsew signal output
rlabel metal3 s 0 154504 800 154624 6 data_arrays_0_0_ext_ram_addr1[2]
port 3 nsew signal output
rlabel metal3 s 0 155184 800 155304 6 data_arrays_0_0_ext_ram_addr1[3]
port 4 nsew signal output
rlabel metal3 s 0 155864 800 155984 6 data_arrays_0_0_ext_ram_addr1[4]
port 5 nsew signal output
rlabel metal3 s 0 156544 800 156664 6 data_arrays_0_0_ext_ram_addr1[5]
port 6 nsew signal output
rlabel metal3 s 0 157224 800 157344 6 data_arrays_0_0_ext_ram_addr1[6]
port 7 nsew signal output
rlabel metal3 s 0 157904 800 158024 6 data_arrays_0_0_ext_ram_addr1[7]
port 8 nsew signal output
rlabel metal3 s 0 158720 800 158840 6 data_arrays_0_0_ext_ram_addr1[8]
port 9 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 data_arrays_0_0_ext_ram_addr[0]
port 10 nsew signal output
rlabel metal3 s 0 90992 800 91112 6 data_arrays_0_0_ext_ram_addr[1]
port 11 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 data_arrays_0_0_ext_ram_addr[2]
port 12 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 data_arrays_0_0_ext_ram_addr[3]
port 13 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 data_arrays_0_0_ext_ram_addr[4]
port 14 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 data_arrays_0_0_ext_ram_addr[5]
port 15 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 data_arrays_0_0_ext_ram_addr[6]
port 16 nsew signal output
rlabel metal3 s 0 95344 800 95464 6 data_arrays_0_0_ext_ram_addr[7]
port 17 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 data_arrays_0_0_ext_ram_addr[8]
port 18 nsew signal output
rlabel metal3 s 0 96704 800 96824 6 data_arrays_0_0_ext_ram_clk
port 19 nsew signal output
rlabel metal3 s 0 147432 800 147552 6 data_arrays_0_0_ext_ram_csb1[0]
port 20 nsew signal output
rlabel metal3 s 0 148112 800 148232 6 data_arrays_0_0_ext_ram_csb1[1]
port 21 nsew signal output
rlabel metal3 s 0 148792 800 148912 6 data_arrays_0_0_ext_ram_csb1[2]
port 22 nsew signal output
rlabel metal3 s 0 149472 800 149592 6 data_arrays_0_0_ext_ram_csb1[3]
port 23 nsew signal output
rlabel metal3 s 0 150152 800 150272 6 data_arrays_0_0_ext_ram_csb1[4]
port 24 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 data_arrays_0_0_ext_ram_csb1[5]
port 25 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 data_arrays_0_0_ext_ram_csb1[6]
port 26 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 data_arrays_0_0_ext_ram_csb1[7]
port 27 nsew signal output
rlabel metal3 s 0 143896 800 144016 6 data_arrays_0_0_ext_ram_csb[0]
port 28 nsew signal output
rlabel metal3 s 0 144576 800 144696 6 data_arrays_0_0_ext_ram_csb[1]
port 29 nsew signal output
rlabel metal3 s 0 145256 800 145376 6 data_arrays_0_0_ext_ram_csb[2]
port 30 nsew signal output
rlabel metal3 s 0 145936 800 146056 6 data_arrays_0_0_ext_ram_csb[3]
port 31 nsew signal output
rlabel metal3 s 0 280 800 400 6 data_arrays_0_0_ext_ram_rdata0[0]
port 32 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 data_arrays_0_0_ext_ram_rdata0[10]
port 33 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 data_arrays_0_0_ext_ram_rdata0[11]
port 34 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 data_arrays_0_0_ext_ram_rdata0[12]
port 35 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 data_arrays_0_0_ext_ram_rdata0[13]
port 36 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 data_arrays_0_0_ext_ram_rdata0[14]
port 37 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 data_arrays_0_0_ext_ram_rdata0[15]
port 38 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 data_arrays_0_0_ext_ram_rdata0[16]
port 39 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 data_arrays_0_0_ext_ram_rdata0[17]
port 40 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 data_arrays_0_0_ext_ram_rdata0[18]
port 41 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 data_arrays_0_0_ext_ram_rdata0[19]
port 42 nsew signal input
rlabel metal3 s 0 960 800 1080 6 data_arrays_0_0_ext_ram_rdata0[1]
port 43 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 data_arrays_0_0_ext_ram_rdata0[20]
port 44 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 data_arrays_0_0_ext_ram_rdata0[21]
port 45 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 data_arrays_0_0_ext_ram_rdata0[22]
port 46 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 data_arrays_0_0_ext_ram_rdata0[23]
port 47 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 data_arrays_0_0_ext_ram_rdata0[24]
port 48 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 data_arrays_0_0_ext_ram_rdata0[25]
port 49 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 data_arrays_0_0_ext_ram_rdata0[26]
port 50 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 data_arrays_0_0_ext_ram_rdata0[27]
port 51 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 data_arrays_0_0_ext_ram_rdata0[28]
port 52 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 data_arrays_0_0_ext_ram_rdata0[29]
port 53 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 data_arrays_0_0_ext_ram_rdata0[2]
port 54 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 data_arrays_0_0_ext_ram_rdata0[30]
port 55 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 data_arrays_0_0_ext_ram_rdata0[31]
port 56 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 data_arrays_0_0_ext_ram_rdata0[32]
port 57 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 data_arrays_0_0_ext_ram_rdata0[33]
port 58 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 data_arrays_0_0_ext_ram_rdata0[34]
port 59 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 data_arrays_0_0_ext_ram_rdata0[35]
port 60 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 data_arrays_0_0_ext_ram_rdata0[36]
port 61 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 data_arrays_0_0_ext_ram_rdata0[37]
port 62 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 data_arrays_0_0_ext_ram_rdata0[38]
port 63 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 data_arrays_0_0_ext_ram_rdata0[39]
port 64 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 data_arrays_0_0_ext_ram_rdata0[3]
port 65 nsew signal input
rlabel metal3 s 0 28432 800 28552 6 data_arrays_0_0_ext_ram_rdata0[40]
port 66 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 data_arrays_0_0_ext_ram_rdata0[41]
port 67 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 data_arrays_0_0_ext_ram_rdata0[42]
port 68 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 data_arrays_0_0_ext_ram_rdata0[43]
port 69 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 data_arrays_0_0_ext_ram_rdata0[44]
port 70 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 data_arrays_0_0_ext_ram_rdata0[45]
port 71 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 data_arrays_0_0_ext_ram_rdata0[46]
port 72 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 data_arrays_0_0_ext_ram_rdata0[47]
port 73 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 data_arrays_0_0_ext_ram_rdata0[48]
port 74 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 data_arrays_0_0_ext_ram_rdata0[49]
port 75 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 data_arrays_0_0_ext_ram_rdata0[4]
port 76 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 data_arrays_0_0_ext_ram_rdata0[50]
port 77 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 data_arrays_0_0_ext_ram_rdata0[51]
port 78 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 data_arrays_0_0_ext_ram_rdata0[52]
port 79 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 data_arrays_0_0_ext_ram_rdata0[53]
port 80 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 data_arrays_0_0_ext_ram_rdata0[54]
port 81 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 data_arrays_0_0_ext_ram_rdata0[55]
port 82 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 data_arrays_0_0_ext_ram_rdata0[56]
port 83 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 data_arrays_0_0_ext_ram_rdata0[57]
port 84 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 data_arrays_0_0_ext_ram_rdata0[58]
port 85 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 data_arrays_0_0_ext_ram_rdata0[59]
port 86 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 data_arrays_0_0_ext_ram_rdata0[5]
port 87 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 data_arrays_0_0_ext_ram_rdata0[60]
port 88 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 data_arrays_0_0_ext_ram_rdata0[61]
port 89 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 data_arrays_0_0_ext_ram_rdata0[62]
port 90 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 data_arrays_0_0_ext_ram_rdata0[63]
port 91 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 data_arrays_0_0_ext_ram_rdata0[6]
port 92 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 data_arrays_0_0_ext_ram_rdata0[7]
port 93 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 data_arrays_0_0_ext_ram_rdata0[8]
port 94 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 data_arrays_0_0_ext_ram_rdata0[9]
port 95 nsew signal input
rlabel metal3 s 0 45296 800 45416 6 data_arrays_0_0_ext_ram_rdata1[0]
port 96 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 data_arrays_0_0_ext_ram_rdata1[10]
port 97 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 data_arrays_0_0_ext_ram_rdata1[11]
port 98 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 data_arrays_0_0_ext_ram_rdata1[12]
port 99 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 data_arrays_0_0_ext_ram_rdata1[13]
port 100 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 data_arrays_0_0_ext_ram_rdata1[14]
port 101 nsew signal input
rlabel metal3 s 0 55904 800 56024 6 data_arrays_0_0_ext_ram_rdata1[15]
port 102 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 data_arrays_0_0_ext_ram_rdata1[16]
port 103 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 data_arrays_0_0_ext_ram_rdata1[17]
port 104 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 data_arrays_0_0_ext_ram_rdata1[18]
port 105 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 data_arrays_0_0_ext_ram_rdata1[19]
port 106 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 data_arrays_0_0_ext_ram_rdata1[1]
port 107 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 data_arrays_0_0_ext_ram_rdata1[20]
port 108 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 data_arrays_0_0_ext_ram_rdata1[21]
port 109 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 data_arrays_0_0_ext_ram_rdata1[22]
port 110 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 data_arrays_0_0_ext_ram_rdata1[23]
port 111 nsew signal input
rlabel metal3 s 0 62160 800 62280 6 data_arrays_0_0_ext_ram_rdata1[24]
port 112 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 data_arrays_0_0_ext_ram_rdata1[25]
port 113 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 data_arrays_0_0_ext_ram_rdata1[26]
port 114 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 data_arrays_0_0_ext_ram_rdata1[27]
port 115 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 data_arrays_0_0_ext_ram_rdata1[28]
port 116 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 data_arrays_0_0_ext_ram_rdata1[29]
port 117 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 data_arrays_0_0_ext_ram_rdata1[2]
port 118 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 data_arrays_0_0_ext_ram_rdata1[30]
port 119 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 data_arrays_0_0_ext_ram_rdata1[31]
port 120 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 data_arrays_0_0_ext_ram_rdata1[32]
port 121 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 data_arrays_0_0_ext_ram_rdata1[33]
port 122 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 data_arrays_0_0_ext_ram_rdata1[34]
port 123 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 data_arrays_0_0_ext_ram_rdata1[35]
port 124 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 data_arrays_0_0_ext_ram_rdata1[36]
port 125 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 data_arrays_0_0_ext_ram_rdata1[37]
port 126 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 data_arrays_0_0_ext_ram_rdata1[38]
port 127 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 data_arrays_0_0_ext_ram_rdata1[39]
port 128 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 data_arrays_0_0_ext_ram_rdata1[3]
port 129 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 data_arrays_0_0_ext_ram_rdata1[40]
port 130 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 data_arrays_0_0_ext_ram_rdata1[41]
port 131 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 data_arrays_0_0_ext_ram_rdata1[42]
port 132 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 data_arrays_0_0_ext_ram_rdata1[43]
port 133 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 data_arrays_0_0_ext_ram_rdata1[44]
port 134 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 data_arrays_0_0_ext_ram_rdata1[45]
port 135 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 data_arrays_0_0_ext_ram_rdata1[46]
port 136 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 data_arrays_0_0_ext_ram_rdata1[47]
port 137 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 data_arrays_0_0_ext_ram_rdata1[48]
port 138 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 data_arrays_0_0_ext_ram_rdata1[49]
port 139 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 data_arrays_0_0_ext_ram_rdata1[4]
port 140 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 data_arrays_0_0_ext_ram_rdata1[50]
port 141 nsew signal input
rlabel metal3 s 0 81200 800 81320 6 data_arrays_0_0_ext_ram_rdata1[51]
port 142 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 data_arrays_0_0_ext_ram_rdata1[52]
port 143 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 data_arrays_0_0_ext_ram_rdata1[53]
port 144 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 data_arrays_0_0_ext_ram_rdata1[54]
port 145 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 data_arrays_0_0_ext_ram_rdata1[55]
port 146 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 data_arrays_0_0_ext_ram_rdata1[56]
port 147 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 data_arrays_0_0_ext_ram_rdata1[57]
port 148 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 data_arrays_0_0_ext_ram_rdata1[58]
port 149 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 data_arrays_0_0_ext_ram_rdata1[59]
port 150 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 data_arrays_0_0_ext_ram_rdata1[5]
port 151 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 data_arrays_0_0_ext_ram_rdata1[60]
port 152 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 data_arrays_0_0_ext_ram_rdata1[61]
port 153 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 data_arrays_0_0_ext_ram_rdata1[62]
port 154 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 data_arrays_0_0_ext_ram_rdata1[63]
port 155 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 data_arrays_0_0_ext_ram_rdata1[6]
port 156 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 data_arrays_0_0_ext_ram_rdata1[7]
port 157 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 data_arrays_0_0_ext_ram_rdata1[8]
port 158 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 data_arrays_0_0_ext_ram_rdata1[9]
port 159 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 data_arrays_0_0_ext_ram_rdata2[0]
port 160 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 data_arrays_0_0_ext_ram_rdata2[10]
port 161 nsew signal input
rlabel metal3 s 0 167152 800 167272 6 data_arrays_0_0_ext_ram_rdata2[11]
port 162 nsew signal input
rlabel metal3 s 0 167832 800 167952 6 data_arrays_0_0_ext_ram_rdata2[12]
port 163 nsew signal input
rlabel metal3 s 0 168512 800 168632 6 data_arrays_0_0_ext_ram_rdata2[13]
port 164 nsew signal input
rlabel metal3 s 0 169192 800 169312 6 data_arrays_0_0_ext_ram_rdata2[14]
port 165 nsew signal input
rlabel metal3 s 0 169872 800 169992 6 data_arrays_0_0_ext_ram_rdata2[15]
port 166 nsew signal input
rlabel metal3 s 0 170688 800 170808 6 data_arrays_0_0_ext_ram_rdata2[16]
port 167 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 data_arrays_0_0_ext_ram_rdata2[17]
port 168 nsew signal input
rlabel metal3 s 0 172048 800 172168 6 data_arrays_0_0_ext_ram_rdata2[18]
port 169 nsew signal input
rlabel metal3 s 0 172728 800 172848 6 data_arrays_0_0_ext_ram_rdata2[19]
port 170 nsew signal input
rlabel metal3 s 0 160080 800 160200 6 data_arrays_0_0_ext_ram_rdata2[1]
port 171 nsew signal input
rlabel metal3 s 0 173408 800 173528 6 data_arrays_0_0_ext_ram_rdata2[20]
port 172 nsew signal input
rlabel metal3 s 0 174224 800 174344 6 data_arrays_0_0_ext_ram_rdata2[21]
port 173 nsew signal input
rlabel metal3 s 0 174904 800 175024 6 data_arrays_0_0_ext_ram_rdata2[22]
port 174 nsew signal input
rlabel metal3 s 0 175584 800 175704 6 data_arrays_0_0_ext_ram_rdata2[23]
port 175 nsew signal input
rlabel metal3 s 0 176264 800 176384 6 data_arrays_0_0_ext_ram_rdata2[24]
port 176 nsew signal input
rlabel metal3 s 0 176944 800 177064 6 data_arrays_0_0_ext_ram_rdata2[25]
port 177 nsew signal input
rlabel metal3 s 0 177624 800 177744 6 data_arrays_0_0_ext_ram_rdata2[26]
port 178 nsew signal input
rlabel metal3 s 0 178440 800 178560 6 data_arrays_0_0_ext_ram_rdata2[27]
port 179 nsew signal input
rlabel metal3 s 0 179120 800 179240 6 data_arrays_0_0_ext_ram_rdata2[28]
port 180 nsew signal input
rlabel metal3 s 0 179800 800 179920 6 data_arrays_0_0_ext_ram_rdata2[29]
port 181 nsew signal input
rlabel metal3 s 0 160760 800 160880 6 data_arrays_0_0_ext_ram_rdata2[2]
port 182 nsew signal input
rlabel metal3 s 0 180480 800 180600 6 data_arrays_0_0_ext_ram_rdata2[30]
port 183 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 data_arrays_0_0_ext_ram_rdata2[31]
port 184 nsew signal input
rlabel metal3 s 0 181840 800 181960 6 data_arrays_0_0_ext_ram_rdata2[32]
port 185 nsew signal input
rlabel metal3 s 0 182656 800 182776 6 data_arrays_0_0_ext_ram_rdata2[33]
port 186 nsew signal input
rlabel metal3 s 0 183336 800 183456 6 data_arrays_0_0_ext_ram_rdata2[34]
port 187 nsew signal input
rlabel metal3 s 0 184016 800 184136 6 data_arrays_0_0_ext_ram_rdata2[35]
port 188 nsew signal input
rlabel metal3 s 0 184696 800 184816 6 data_arrays_0_0_ext_ram_rdata2[36]
port 189 nsew signal input
rlabel metal3 s 0 185376 800 185496 6 data_arrays_0_0_ext_ram_rdata2[37]
port 190 nsew signal input
rlabel metal3 s 0 186192 800 186312 6 data_arrays_0_0_ext_ram_rdata2[38]
port 191 nsew signal input
rlabel metal3 s 0 186872 800 186992 6 data_arrays_0_0_ext_ram_rdata2[39]
port 192 nsew signal input
rlabel metal3 s 0 161440 800 161560 6 data_arrays_0_0_ext_ram_rdata2[3]
port 193 nsew signal input
rlabel metal3 s 0 187552 800 187672 6 data_arrays_0_0_ext_ram_rdata2[40]
port 194 nsew signal input
rlabel metal3 s 0 188232 800 188352 6 data_arrays_0_0_ext_ram_rdata2[41]
port 195 nsew signal input
rlabel metal3 s 0 188912 800 189032 6 data_arrays_0_0_ext_ram_rdata2[42]
port 196 nsew signal input
rlabel metal3 s 0 189592 800 189712 6 data_arrays_0_0_ext_ram_rdata2[43]
port 197 nsew signal input
rlabel metal3 s 0 190408 800 190528 6 data_arrays_0_0_ext_ram_rdata2[44]
port 198 nsew signal input
rlabel metal3 s 0 191088 800 191208 6 data_arrays_0_0_ext_ram_rdata2[45]
port 199 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 data_arrays_0_0_ext_ram_rdata2[46]
port 200 nsew signal input
rlabel metal3 s 0 192448 800 192568 6 data_arrays_0_0_ext_ram_rdata2[47]
port 201 nsew signal input
rlabel metal3 s 0 193128 800 193248 6 data_arrays_0_0_ext_ram_rdata2[48]
port 202 nsew signal input
rlabel metal3 s 0 193944 800 194064 6 data_arrays_0_0_ext_ram_rdata2[49]
port 203 nsew signal input
rlabel metal3 s 0 162120 800 162240 6 data_arrays_0_0_ext_ram_rdata2[4]
port 204 nsew signal input
rlabel metal3 s 0 194624 800 194744 6 data_arrays_0_0_ext_ram_rdata2[50]
port 205 nsew signal input
rlabel metal3 s 0 195304 800 195424 6 data_arrays_0_0_ext_ram_rdata2[51]
port 206 nsew signal input
rlabel metal3 s 0 195984 800 196104 6 data_arrays_0_0_ext_ram_rdata2[52]
port 207 nsew signal input
rlabel metal3 s 0 196664 800 196784 6 data_arrays_0_0_ext_ram_rdata2[53]
port 208 nsew signal input
rlabel metal3 s 0 197344 800 197464 6 data_arrays_0_0_ext_ram_rdata2[54]
port 209 nsew signal input
rlabel metal3 s 0 198160 800 198280 6 data_arrays_0_0_ext_ram_rdata2[55]
port 210 nsew signal input
rlabel metal3 s 0 198840 800 198960 6 data_arrays_0_0_ext_ram_rdata2[56]
port 211 nsew signal input
rlabel metal3 s 0 199520 800 199640 6 data_arrays_0_0_ext_ram_rdata2[57]
port 212 nsew signal input
rlabel metal3 s 0 200200 800 200320 6 data_arrays_0_0_ext_ram_rdata2[58]
port 213 nsew signal input
rlabel metal3 s 0 200880 800 201000 6 data_arrays_0_0_ext_ram_rdata2[59]
port 214 nsew signal input
rlabel metal3 s 0 162936 800 163056 6 data_arrays_0_0_ext_ram_rdata2[5]
port 215 nsew signal input
rlabel metal3 s 0 201560 800 201680 6 data_arrays_0_0_ext_ram_rdata2[60]
port 216 nsew signal input
rlabel metal3 s 0 202376 800 202496 6 data_arrays_0_0_ext_ram_rdata2[61]
port 217 nsew signal input
rlabel metal3 s 0 203056 800 203176 6 data_arrays_0_0_ext_ram_rdata2[62]
port 218 nsew signal input
rlabel metal3 s 0 203736 800 203856 6 data_arrays_0_0_ext_ram_rdata2[63]
port 219 nsew signal input
rlabel metal3 s 0 163616 800 163736 6 data_arrays_0_0_ext_ram_rdata2[6]
port 220 nsew signal input
rlabel metal3 s 0 164296 800 164416 6 data_arrays_0_0_ext_ram_rdata2[7]
port 221 nsew signal input
rlabel metal3 s 0 164976 800 165096 6 data_arrays_0_0_ext_ram_rdata2[8]
port 222 nsew signal input
rlabel metal3 s 0 165656 800 165776 6 data_arrays_0_0_ext_ram_rdata2[9]
port 223 nsew signal input
rlabel metal3 s 0 204416 800 204536 6 data_arrays_0_0_ext_ram_rdata3[0]
port 224 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 data_arrays_0_0_ext_ram_rdata3[10]
port 225 nsew signal input
rlabel metal3 s 0 212168 800 212288 6 data_arrays_0_0_ext_ram_rdata3[11]
port 226 nsew signal input
rlabel metal3 s 0 212848 800 212968 6 data_arrays_0_0_ext_ram_rdata3[12]
port 227 nsew signal input
rlabel metal3 s 0 213664 800 213784 6 data_arrays_0_0_ext_ram_rdata3[13]
port 228 nsew signal input
rlabel metal3 s 0 214344 800 214464 6 data_arrays_0_0_ext_ram_rdata3[14]
port 229 nsew signal input
rlabel metal3 s 0 215024 800 215144 6 data_arrays_0_0_ext_ram_rdata3[15]
port 230 nsew signal input
rlabel metal3 s 0 215704 800 215824 6 data_arrays_0_0_ext_ram_rdata3[16]
port 231 nsew signal input
rlabel metal3 s 0 216384 800 216504 6 data_arrays_0_0_ext_ram_rdata3[17]
port 232 nsew signal input
rlabel metal3 s 0 217064 800 217184 6 data_arrays_0_0_ext_ram_rdata3[18]
port 233 nsew signal input
rlabel metal3 s 0 217880 800 218000 6 data_arrays_0_0_ext_ram_rdata3[19]
port 234 nsew signal input
rlabel metal3 s 0 205096 800 205216 6 data_arrays_0_0_ext_ram_rdata3[1]
port 235 nsew signal input
rlabel metal3 s 0 218560 800 218680 6 data_arrays_0_0_ext_ram_rdata3[20]
port 236 nsew signal input
rlabel metal3 s 0 219240 800 219360 6 data_arrays_0_0_ext_ram_rdata3[21]
port 237 nsew signal input
rlabel metal3 s 0 219920 800 220040 6 data_arrays_0_0_ext_ram_rdata3[22]
port 238 nsew signal input
rlabel metal3 s 0 220600 800 220720 6 data_arrays_0_0_ext_ram_rdata3[23]
port 239 nsew signal input
rlabel metal3 s 0 221280 800 221400 6 data_arrays_0_0_ext_ram_rdata3[24]
port 240 nsew signal input
rlabel metal3 s 0 222096 800 222216 6 data_arrays_0_0_ext_ram_rdata3[25]
port 241 nsew signal input
rlabel metal3 s 0 222776 800 222896 6 data_arrays_0_0_ext_ram_rdata3[26]
port 242 nsew signal input
rlabel metal3 s 0 223456 800 223576 6 data_arrays_0_0_ext_ram_rdata3[27]
port 243 nsew signal input
rlabel metal3 s 0 224136 800 224256 6 data_arrays_0_0_ext_ram_rdata3[28]
port 244 nsew signal input
rlabel metal3 s 0 224816 800 224936 6 data_arrays_0_0_ext_ram_rdata3[29]
port 245 nsew signal input
rlabel metal3 s 0 205912 800 206032 6 data_arrays_0_0_ext_ram_rdata3[2]
port 246 nsew signal input
rlabel metal3 s 0 225632 800 225752 6 data_arrays_0_0_ext_ram_rdata3[30]
port 247 nsew signal input
rlabel metal3 s 0 226312 800 226432 6 data_arrays_0_0_ext_ram_rdata3[31]
port 248 nsew signal input
rlabel metal3 s 0 226992 800 227112 6 data_arrays_0_0_ext_ram_rdata3[32]
port 249 nsew signal input
rlabel metal3 s 0 227672 800 227792 6 data_arrays_0_0_ext_ram_rdata3[33]
port 250 nsew signal input
rlabel metal3 s 0 228352 800 228472 6 data_arrays_0_0_ext_ram_rdata3[34]
port 251 nsew signal input
rlabel metal3 s 0 229032 800 229152 6 data_arrays_0_0_ext_ram_rdata3[35]
port 252 nsew signal input
rlabel metal3 s 0 229848 800 229968 6 data_arrays_0_0_ext_ram_rdata3[36]
port 253 nsew signal input
rlabel metal3 s 0 230528 800 230648 6 data_arrays_0_0_ext_ram_rdata3[37]
port 254 nsew signal input
rlabel metal3 s 0 231208 800 231328 6 data_arrays_0_0_ext_ram_rdata3[38]
port 255 nsew signal input
rlabel metal3 s 0 231888 800 232008 6 data_arrays_0_0_ext_ram_rdata3[39]
port 256 nsew signal input
rlabel metal3 s 0 206592 800 206712 6 data_arrays_0_0_ext_ram_rdata3[3]
port 257 nsew signal input
rlabel metal3 s 0 232568 800 232688 6 data_arrays_0_0_ext_ram_rdata3[40]
port 258 nsew signal input
rlabel metal3 s 0 233248 800 233368 6 data_arrays_0_0_ext_ram_rdata3[41]
port 259 nsew signal input
rlabel metal3 s 0 234064 800 234184 6 data_arrays_0_0_ext_ram_rdata3[42]
port 260 nsew signal input
rlabel metal3 s 0 234744 800 234864 6 data_arrays_0_0_ext_ram_rdata3[43]
port 261 nsew signal input
rlabel metal3 s 0 235424 800 235544 6 data_arrays_0_0_ext_ram_rdata3[44]
port 262 nsew signal input
rlabel metal3 s 0 236104 800 236224 6 data_arrays_0_0_ext_ram_rdata3[45]
port 263 nsew signal input
rlabel metal3 s 0 236784 800 236904 6 data_arrays_0_0_ext_ram_rdata3[46]
port 264 nsew signal input
rlabel metal3 s 0 237600 800 237720 6 data_arrays_0_0_ext_ram_rdata3[47]
port 265 nsew signal input
rlabel metal3 s 0 238280 800 238400 6 data_arrays_0_0_ext_ram_rdata3[48]
port 266 nsew signal input
rlabel metal3 s 0 238960 800 239080 6 data_arrays_0_0_ext_ram_rdata3[49]
port 267 nsew signal input
rlabel metal3 s 0 207272 800 207392 6 data_arrays_0_0_ext_ram_rdata3[4]
port 268 nsew signal input
rlabel metal3 s 0 239640 800 239760 6 data_arrays_0_0_ext_ram_rdata3[50]
port 269 nsew signal input
rlabel metal3 s 0 240320 800 240440 6 data_arrays_0_0_ext_ram_rdata3[51]
port 270 nsew signal input
rlabel metal3 s 0 241000 800 241120 6 data_arrays_0_0_ext_ram_rdata3[52]
port 271 nsew signal input
rlabel metal3 s 0 241816 800 241936 6 data_arrays_0_0_ext_ram_rdata3[53]
port 272 nsew signal input
rlabel metal3 s 0 242496 800 242616 6 data_arrays_0_0_ext_ram_rdata3[54]
port 273 nsew signal input
rlabel metal3 s 0 243176 800 243296 6 data_arrays_0_0_ext_ram_rdata3[55]
port 274 nsew signal input
rlabel metal3 s 0 243856 800 243976 6 data_arrays_0_0_ext_ram_rdata3[56]
port 275 nsew signal input
rlabel metal3 s 0 244536 800 244656 6 data_arrays_0_0_ext_ram_rdata3[57]
port 276 nsew signal input
rlabel metal3 s 0 245352 800 245472 6 data_arrays_0_0_ext_ram_rdata3[58]
port 277 nsew signal input
rlabel metal3 s 0 246032 800 246152 6 data_arrays_0_0_ext_ram_rdata3[59]
port 278 nsew signal input
rlabel metal3 s 0 207952 800 208072 6 data_arrays_0_0_ext_ram_rdata3[5]
port 279 nsew signal input
rlabel metal3 s 0 246712 800 246832 6 data_arrays_0_0_ext_ram_rdata3[60]
port 280 nsew signal input
rlabel metal3 s 0 247392 800 247512 6 data_arrays_0_0_ext_ram_rdata3[61]
port 281 nsew signal input
rlabel metal3 s 0 248072 800 248192 6 data_arrays_0_0_ext_ram_rdata3[62]
port 282 nsew signal input
rlabel metal3 s 0 248752 800 248872 6 data_arrays_0_0_ext_ram_rdata3[63]
port 283 nsew signal input
rlabel metal3 s 0 208632 800 208752 6 data_arrays_0_0_ext_ram_rdata3[6]
port 284 nsew signal input
rlabel metal3 s 0 209312 800 209432 6 data_arrays_0_0_ext_ram_rdata3[7]
port 285 nsew signal input
rlabel metal3 s 0 210128 800 210248 6 data_arrays_0_0_ext_ram_rdata3[8]
port 286 nsew signal input
rlabel metal3 s 0 210808 800 210928 6 data_arrays_0_0_ext_ram_rdata3[9]
port 287 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 data_arrays_0_0_ext_ram_wdata[0]
port 288 nsew signal output
rlabel metal3 s 0 104456 800 104576 6 data_arrays_0_0_ext_ram_wdata[10]
port 289 nsew signal output
rlabel metal3 s 0 105136 800 105256 6 data_arrays_0_0_ext_ram_wdata[11]
port 290 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 data_arrays_0_0_ext_ram_wdata[12]
port 291 nsew signal output
rlabel metal3 s 0 106496 800 106616 6 data_arrays_0_0_ext_ram_wdata[13]
port 292 nsew signal output
rlabel metal3 s 0 107312 800 107432 6 data_arrays_0_0_ext_ram_wdata[14]
port 293 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 data_arrays_0_0_ext_ram_wdata[15]
port 294 nsew signal output
rlabel metal3 s 0 108672 800 108792 6 data_arrays_0_0_ext_ram_wdata[16]
port 295 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 data_arrays_0_0_ext_ram_wdata[17]
port 296 nsew signal output
rlabel metal3 s 0 110032 800 110152 6 data_arrays_0_0_ext_ram_wdata[18]
port 297 nsew signal output
rlabel metal3 s 0 110712 800 110832 6 data_arrays_0_0_ext_ram_wdata[19]
port 298 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 data_arrays_0_0_ext_ram_wdata[1]
port 299 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 data_arrays_0_0_ext_ram_wdata[20]
port 300 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 data_arrays_0_0_ext_ram_wdata[21]
port 301 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 data_arrays_0_0_ext_ram_wdata[22]
port 302 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 data_arrays_0_0_ext_ram_wdata[23]
port 303 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 data_arrays_0_0_ext_ram_wdata[24]
port 304 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 data_arrays_0_0_ext_ram_wdata[25]
port 305 nsew signal output
rlabel metal3 s 0 115744 800 115864 6 data_arrays_0_0_ext_ram_wdata[26]
port 306 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 data_arrays_0_0_ext_ram_wdata[27]
port 307 nsew signal output
rlabel metal3 s 0 117104 800 117224 6 data_arrays_0_0_ext_ram_wdata[28]
port 308 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 data_arrays_0_0_ext_ram_wdata[29]
port 309 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 data_arrays_0_0_ext_ram_wdata[2]
port 310 nsew signal output
rlabel metal3 s 0 118464 800 118584 6 data_arrays_0_0_ext_ram_wdata[30]
port 311 nsew signal output
rlabel metal3 s 0 119280 800 119400 6 data_arrays_0_0_ext_ram_wdata[31]
port 312 nsew signal output
rlabel metal3 s 0 119960 800 120080 6 data_arrays_0_0_ext_ram_wdata[32]
port 313 nsew signal output
rlabel metal3 s 0 120640 800 120760 6 data_arrays_0_0_ext_ram_wdata[33]
port 314 nsew signal output
rlabel metal3 s 0 121320 800 121440 6 data_arrays_0_0_ext_ram_wdata[34]
port 315 nsew signal output
rlabel metal3 s 0 122000 800 122120 6 data_arrays_0_0_ext_ram_wdata[35]
port 316 nsew signal output
rlabel metal3 s 0 122816 800 122936 6 data_arrays_0_0_ext_ram_wdata[36]
port 317 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 data_arrays_0_0_ext_ram_wdata[37]
port 318 nsew signal output
rlabel metal3 s 0 124176 800 124296 6 data_arrays_0_0_ext_ram_wdata[38]
port 319 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 data_arrays_0_0_ext_ram_wdata[39]
port 320 nsew signal output
rlabel metal3 s 0 99560 800 99680 6 data_arrays_0_0_ext_ram_wdata[3]
port 321 nsew signal output
rlabel metal3 s 0 125536 800 125656 6 data_arrays_0_0_ext_ram_wdata[40]
port 322 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 data_arrays_0_0_ext_ram_wdata[41]
port 323 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 data_arrays_0_0_ext_ram_wdata[42]
port 324 nsew signal output
rlabel metal3 s 0 127712 800 127832 6 data_arrays_0_0_ext_ram_wdata[43]
port 325 nsew signal output
rlabel metal3 s 0 128392 800 128512 6 data_arrays_0_0_ext_ram_wdata[44]
port 326 nsew signal output
rlabel metal3 s 0 129072 800 129192 6 data_arrays_0_0_ext_ram_wdata[45]
port 327 nsew signal output
rlabel metal3 s 0 129752 800 129872 6 data_arrays_0_0_ext_ram_wdata[46]
port 328 nsew signal output
rlabel metal3 s 0 130432 800 130552 6 data_arrays_0_0_ext_ram_wdata[47]
port 329 nsew signal output
rlabel metal3 s 0 131248 800 131368 6 data_arrays_0_0_ext_ram_wdata[48]
port 330 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 data_arrays_0_0_ext_ram_wdata[49]
port 331 nsew signal output
rlabel metal3 s 0 100240 800 100360 6 data_arrays_0_0_ext_ram_wdata[4]
port 332 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 data_arrays_0_0_ext_ram_wdata[50]
port 333 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 data_arrays_0_0_ext_ram_wdata[51]
port 334 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 data_arrays_0_0_ext_ram_wdata[52]
port 335 nsew signal output
rlabel metal3 s 0 134784 800 134904 6 data_arrays_0_0_ext_ram_wdata[53]
port 336 nsew signal output
rlabel metal3 s 0 135464 800 135584 6 data_arrays_0_0_ext_ram_wdata[54]
port 337 nsew signal output
rlabel metal3 s 0 136144 800 136264 6 data_arrays_0_0_ext_ram_wdata[55]
port 338 nsew signal output
rlabel metal3 s 0 136824 800 136944 6 data_arrays_0_0_ext_ram_wdata[56]
port 339 nsew signal output
rlabel metal3 s 0 137504 800 137624 6 data_arrays_0_0_ext_ram_wdata[57]
port 340 nsew signal output
rlabel metal3 s 0 138184 800 138304 6 data_arrays_0_0_ext_ram_wdata[58]
port 341 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 data_arrays_0_0_ext_ram_wdata[59]
port 342 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 data_arrays_0_0_ext_ram_wdata[5]
port 343 nsew signal output
rlabel metal3 s 0 139680 800 139800 6 data_arrays_0_0_ext_ram_wdata[60]
port 344 nsew signal output
rlabel metal3 s 0 140360 800 140480 6 data_arrays_0_0_ext_ram_wdata[61]
port 345 nsew signal output
rlabel metal3 s 0 141040 800 141160 6 data_arrays_0_0_ext_ram_wdata[62]
port 346 nsew signal output
rlabel metal3 s 0 141720 800 141840 6 data_arrays_0_0_ext_ram_wdata[63]
port 347 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 data_arrays_0_0_ext_ram_wdata[6]
port 348 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 data_arrays_0_0_ext_ram_wdata[7]
port 349 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 data_arrays_0_0_ext_ram_wdata[8]
port 350 nsew signal output
rlabel metal3 s 0 103776 800 103896 6 data_arrays_0_0_ext_ram_wdata[9]
port 351 nsew signal output
rlabel metal3 s 0 146752 800 146872 6 data_arrays_0_0_ext_ram_web
port 352 nsew signal output
rlabel metal3 s 0 142536 800 142656 6 data_arrays_0_0_ext_ram_wmask[0]
port 353 nsew signal output
rlabel metal3 s 0 143216 800 143336 6 data_arrays_0_0_ext_ram_wmask[1]
port 354 nsew signal output
rlabel metal3 s 352720 207408 353520 207528 6 data_arrays_0_ext_ram_addr1[0]
port 355 nsew signal output
rlabel metal3 s 352720 208496 353520 208616 6 data_arrays_0_ext_ram_addr1[1]
port 356 nsew signal output
rlabel metal3 s 352720 209584 353520 209704 6 data_arrays_0_ext_ram_addr1[2]
port 357 nsew signal output
rlabel metal3 s 352720 210672 353520 210792 6 data_arrays_0_ext_ram_addr1[3]
port 358 nsew signal output
rlabel metal3 s 352720 211760 353520 211880 6 data_arrays_0_ext_ram_addr1[4]
port 359 nsew signal output
rlabel metal3 s 352720 212848 353520 212968 6 data_arrays_0_ext_ram_addr1[5]
port 360 nsew signal output
rlabel metal3 s 352720 213936 353520 214056 6 data_arrays_0_ext_ram_addr1[6]
port 361 nsew signal output
rlabel metal3 s 352720 215024 353520 215144 6 data_arrays_0_ext_ram_addr1[7]
port 362 nsew signal output
rlabel metal3 s 352720 216112 353520 216232 6 data_arrays_0_ext_ram_addr1[8]
port 363 nsew signal output
rlabel metal3 s 352720 139136 353520 139256 6 data_arrays_0_ext_ram_addr[0]
port 364 nsew signal output
rlabel metal3 s 352720 140224 353520 140344 6 data_arrays_0_ext_ram_addr[1]
port 365 nsew signal output
rlabel metal3 s 352720 141312 353520 141432 6 data_arrays_0_ext_ram_addr[2]
port 366 nsew signal output
rlabel metal3 s 352720 142400 353520 142520 6 data_arrays_0_ext_ram_addr[3]
port 367 nsew signal output
rlabel metal3 s 352720 143488 353520 143608 6 data_arrays_0_ext_ram_addr[4]
port 368 nsew signal output
rlabel metal3 s 352720 144576 353520 144696 6 data_arrays_0_ext_ram_addr[5]
port 369 nsew signal output
rlabel metal3 s 352720 145664 353520 145784 6 data_arrays_0_ext_ram_addr[6]
port 370 nsew signal output
rlabel metal3 s 352720 146752 353520 146872 6 data_arrays_0_ext_ram_addr[7]
port 371 nsew signal output
rlabel metal3 s 352720 147840 353520 147960 6 data_arrays_0_ext_ram_addr[8]
port 372 nsew signal output
rlabel metal3 s 352720 148928 353520 149048 6 data_arrays_0_ext_ram_clk
port 373 nsew signal output
rlabel metal3 s 352720 198704 353520 198824 6 data_arrays_0_ext_ram_csb1[0]
port 374 nsew signal output
rlabel metal3 s 352720 199792 353520 199912 6 data_arrays_0_ext_ram_csb1[1]
port 375 nsew signal output
rlabel metal3 s 352720 200880 353520 201000 6 data_arrays_0_ext_ram_csb1[2]
port 376 nsew signal output
rlabel metal3 s 352720 201968 353520 202088 6 data_arrays_0_ext_ram_csb1[3]
port 377 nsew signal output
rlabel metal3 s 352720 203056 353520 203176 6 data_arrays_0_ext_ram_csb1[4]
port 378 nsew signal output
rlabel metal3 s 352720 204144 353520 204264 6 data_arrays_0_ext_ram_csb1[5]
port 379 nsew signal output
rlabel metal3 s 352720 205232 353520 205352 6 data_arrays_0_ext_ram_csb1[6]
port 380 nsew signal output
rlabel metal3 s 352720 206320 353520 206440 6 data_arrays_0_ext_ram_csb1[7]
port 381 nsew signal output
rlabel metal3 s 352720 189048 353520 189168 6 data_arrays_0_ext_ram_csb[0]
port 382 nsew signal output
rlabel metal3 s 352720 190136 353520 190256 6 data_arrays_0_ext_ram_csb[1]
port 383 nsew signal output
rlabel metal3 s 352720 191224 353520 191344 6 data_arrays_0_ext_ram_csb[2]
port 384 nsew signal output
rlabel metal3 s 352720 192312 353520 192432 6 data_arrays_0_ext_ram_csb[3]
port 385 nsew signal output
rlabel metal3 s 352720 193400 353520 193520 6 data_arrays_0_ext_ram_csb[4]
port 386 nsew signal output
rlabel metal3 s 352720 194488 353520 194608 6 data_arrays_0_ext_ram_csb[5]
port 387 nsew signal output
rlabel metal3 s 352720 195576 353520 195696 6 data_arrays_0_ext_ram_csb[6]
port 388 nsew signal output
rlabel metal3 s 352720 196664 353520 196784 6 data_arrays_0_ext_ram_csb[7]
port 389 nsew signal output
rlabel metal3 s 352720 416 353520 536 6 data_arrays_0_ext_ram_rdata0[0]
port 390 nsew signal input
rlabel metal3 s 352720 11160 353520 11280 6 data_arrays_0_ext_ram_rdata0[10]
port 391 nsew signal input
rlabel metal3 s 352720 12248 353520 12368 6 data_arrays_0_ext_ram_rdata0[11]
port 392 nsew signal input
rlabel metal3 s 352720 13336 353520 13456 6 data_arrays_0_ext_ram_rdata0[12]
port 393 nsew signal input
rlabel metal3 s 352720 14424 353520 14544 6 data_arrays_0_ext_ram_rdata0[13]
port 394 nsew signal input
rlabel metal3 s 352720 15512 353520 15632 6 data_arrays_0_ext_ram_rdata0[14]
port 395 nsew signal input
rlabel metal3 s 352720 16600 353520 16720 6 data_arrays_0_ext_ram_rdata0[15]
port 396 nsew signal input
rlabel metal3 s 352720 17688 353520 17808 6 data_arrays_0_ext_ram_rdata0[16]
port 397 nsew signal input
rlabel metal3 s 352720 18776 353520 18896 6 data_arrays_0_ext_ram_rdata0[17]
port 398 nsew signal input
rlabel metal3 s 352720 19864 353520 19984 6 data_arrays_0_ext_ram_rdata0[18]
port 399 nsew signal input
rlabel metal3 s 352720 20952 353520 21072 6 data_arrays_0_ext_ram_rdata0[19]
port 400 nsew signal input
rlabel metal3 s 352720 1368 353520 1488 6 data_arrays_0_ext_ram_rdata0[1]
port 401 nsew signal input
rlabel metal3 s 352720 22040 353520 22160 6 data_arrays_0_ext_ram_rdata0[20]
port 402 nsew signal input
rlabel metal3 s 352720 23128 353520 23248 6 data_arrays_0_ext_ram_rdata0[21]
port 403 nsew signal input
rlabel metal3 s 352720 24216 353520 24336 6 data_arrays_0_ext_ram_rdata0[22]
port 404 nsew signal input
rlabel metal3 s 352720 25304 353520 25424 6 data_arrays_0_ext_ram_rdata0[23]
port 405 nsew signal input
rlabel metal3 s 352720 26392 353520 26512 6 data_arrays_0_ext_ram_rdata0[24]
port 406 nsew signal input
rlabel metal3 s 352720 27480 353520 27600 6 data_arrays_0_ext_ram_rdata0[25]
port 407 nsew signal input
rlabel metal3 s 352720 28568 353520 28688 6 data_arrays_0_ext_ram_rdata0[26]
port 408 nsew signal input
rlabel metal3 s 352720 29656 353520 29776 6 data_arrays_0_ext_ram_rdata0[27]
port 409 nsew signal input
rlabel metal3 s 352720 30744 353520 30864 6 data_arrays_0_ext_ram_rdata0[28]
port 410 nsew signal input
rlabel metal3 s 352720 31832 353520 31952 6 data_arrays_0_ext_ram_rdata0[29]
port 411 nsew signal input
rlabel metal3 s 352720 2456 353520 2576 6 data_arrays_0_ext_ram_rdata0[2]
port 412 nsew signal input
rlabel metal3 s 352720 32920 353520 33040 6 data_arrays_0_ext_ram_rdata0[30]
port 413 nsew signal input
rlabel metal3 s 352720 34008 353520 34128 6 data_arrays_0_ext_ram_rdata0[31]
port 414 nsew signal input
rlabel metal3 s 352720 3544 353520 3664 6 data_arrays_0_ext_ram_rdata0[3]
port 415 nsew signal input
rlabel metal3 s 352720 4632 353520 4752 6 data_arrays_0_ext_ram_rdata0[4]
port 416 nsew signal input
rlabel metal3 s 352720 5720 353520 5840 6 data_arrays_0_ext_ram_rdata0[5]
port 417 nsew signal input
rlabel metal3 s 352720 6808 353520 6928 6 data_arrays_0_ext_ram_rdata0[6]
port 418 nsew signal input
rlabel metal3 s 352720 7896 353520 8016 6 data_arrays_0_ext_ram_rdata0[7]
port 419 nsew signal input
rlabel metal3 s 352720 8984 353520 9104 6 data_arrays_0_ext_ram_rdata0[8]
port 420 nsew signal input
rlabel metal3 s 352720 10072 353520 10192 6 data_arrays_0_ext_ram_rdata0[9]
port 421 nsew signal input
rlabel metal3 s 352720 35096 353520 35216 6 data_arrays_0_ext_ram_rdata1[0]
port 422 nsew signal input
rlabel metal3 s 352720 45840 353520 45960 6 data_arrays_0_ext_ram_rdata1[10]
port 423 nsew signal input
rlabel metal3 s 352720 46928 353520 47048 6 data_arrays_0_ext_ram_rdata1[11]
port 424 nsew signal input
rlabel metal3 s 352720 48016 353520 48136 6 data_arrays_0_ext_ram_rdata1[12]
port 425 nsew signal input
rlabel metal3 s 352720 49104 353520 49224 6 data_arrays_0_ext_ram_rdata1[13]
port 426 nsew signal input
rlabel metal3 s 352720 50192 353520 50312 6 data_arrays_0_ext_ram_rdata1[14]
port 427 nsew signal input
rlabel metal3 s 352720 51280 353520 51400 6 data_arrays_0_ext_ram_rdata1[15]
port 428 nsew signal input
rlabel metal3 s 352720 52368 353520 52488 6 data_arrays_0_ext_ram_rdata1[16]
port 429 nsew signal input
rlabel metal3 s 352720 53456 353520 53576 6 data_arrays_0_ext_ram_rdata1[17]
port 430 nsew signal input
rlabel metal3 s 352720 54544 353520 54664 6 data_arrays_0_ext_ram_rdata1[18]
port 431 nsew signal input
rlabel metal3 s 352720 55632 353520 55752 6 data_arrays_0_ext_ram_rdata1[19]
port 432 nsew signal input
rlabel metal3 s 352720 36184 353520 36304 6 data_arrays_0_ext_ram_rdata1[1]
port 433 nsew signal input
rlabel metal3 s 352720 56720 353520 56840 6 data_arrays_0_ext_ram_rdata1[20]
port 434 nsew signal input
rlabel metal3 s 352720 57808 353520 57928 6 data_arrays_0_ext_ram_rdata1[21]
port 435 nsew signal input
rlabel metal3 s 352720 58896 353520 59016 6 data_arrays_0_ext_ram_rdata1[22]
port 436 nsew signal input
rlabel metal3 s 352720 59984 353520 60104 6 data_arrays_0_ext_ram_rdata1[23]
port 437 nsew signal input
rlabel metal3 s 352720 61072 353520 61192 6 data_arrays_0_ext_ram_rdata1[24]
port 438 nsew signal input
rlabel metal3 s 352720 62160 353520 62280 6 data_arrays_0_ext_ram_rdata1[25]
port 439 nsew signal input
rlabel metal3 s 352720 63248 353520 63368 6 data_arrays_0_ext_ram_rdata1[26]
port 440 nsew signal input
rlabel metal3 s 352720 64336 353520 64456 6 data_arrays_0_ext_ram_rdata1[27]
port 441 nsew signal input
rlabel metal3 s 352720 65424 353520 65544 6 data_arrays_0_ext_ram_rdata1[28]
port 442 nsew signal input
rlabel metal3 s 352720 66512 353520 66632 6 data_arrays_0_ext_ram_rdata1[29]
port 443 nsew signal input
rlabel metal3 s 352720 37272 353520 37392 6 data_arrays_0_ext_ram_rdata1[2]
port 444 nsew signal input
rlabel metal3 s 352720 67600 353520 67720 6 data_arrays_0_ext_ram_rdata1[30]
port 445 nsew signal input
rlabel metal3 s 352720 68688 353520 68808 6 data_arrays_0_ext_ram_rdata1[31]
port 446 nsew signal input
rlabel metal3 s 352720 38360 353520 38480 6 data_arrays_0_ext_ram_rdata1[3]
port 447 nsew signal input
rlabel metal3 s 352720 39448 353520 39568 6 data_arrays_0_ext_ram_rdata1[4]
port 448 nsew signal input
rlabel metal3 s 352720 40400 353520 40520 6 data_arrays_0_ext_ram_rdata1[5]
port 449 nsew signal input
rlabel metal3 s 352720 41488 353520 41608 6 data_arrays_0_ext_ram_rdata1[6]
port 450 nsew signal input
rlabel metal3 s 352720 42576 353520 42696 6 data_arrays_0_ext_ram_rdata1[7]
port 451 nsew signal input
rlabel metal3 s 352720 43664 353520 43784 6 data_arrays_0_ext_ram_rdata1[8]
port 452 nsew signal input
rlabel metal3 s 352720 44752 353520 44872 6 data_arrays_0_ext_ram_rdata1[9]
port 453 nsew signal input
rlabel metal3 s 352720 69776 353520 69896 6 data_arrays_0_ext_ram_rdata2[0]
port 454 nsew signal input
rlabel metal3 s 352720 80520 353520 80640 6 data_arrays_0_ext_ram_rdata2[10]
port 455 nsew signal input
rlabel metal3 s 352720 81608 353520 81728 6 data_arrays_0_ext_ram_rdata2[11]
port 456 nsew signal input
rlabel metal3 s 352720 82696 353520 82816 6 data_arrays_0_ext_ram_rdata2[12]
port 457 nsew signal input
rlabel metal3 s 352720 83784 353520 83904 6 data_arrays_0_ext_ram_rdata2[13]
port 458 nsew signal input
rlabel metal3 s 352720 84872 353520 84992 6 data_arrays_0_ext_ram_rdata2[14]
port 459 nsew signal input
rlabel metal3 s 352720 85960 353520 86080 6 data_arrays_0_ext_ram_rdata2[15]
port 460 nsew signal input
rlabel metal3 s 352720 87048 353520 87168 6 data_arrays_0_ext_ram_rdata2[16]
port 461 nsew signal input
rlabel metal3 s 352720 88136 353520 88256 6 data_arrays_0_ext_ram_rdata2[17]
port 462 nsew signal input
rlabel metal3 s 352720 89224 353520 89344 6 data_arrays_0_ext_ram_rdata2[18]
port 463 nsew signal input
rlabel metal3 s 352720 90312 353520 90432 6 data_arrays_0_ext_ram_rdata2[19]
port 464 nsew signal input
rlabel metal3 s 352720 70864 353520 70984 6 data_arrays_0_ext_ram_rdata2[1]
port 465 nsew signal input
rlabel metal3 s 352720 91400 353520 91520 6 data_arrays_0_ext_ram_rdata2[20]
port 466 nsew signal input
rlabel metal3 s 352720 92488 353520 92608 6 data_arrays_0_ext_ram_rdata2[21]
port 467 nsew signal input
rlabel metal3 s 352720 93576 353520 93696 6 data_arrays_0_ext_ram_rdata2[22]
port 468 nsew signal input
rlabel metal3 s 352720 94664 353520 94784 6 data_arrays_0_ext_ram_rdata2[23]
port 469 nsew signal input
rlabel metal3 s 352720 95752 353520 95872 6 data_arrays_0_ext_ram_rdata2[24]
port 470 nsew signal input
rlabel metal3 s 352720 96840 353520 96960 6 data_arrays_0_ext_ram_rdata2[25]
port 471 nsew signal input
rlabel metal3 s 352720 97928 353520 98048 6 data_arrays_0_ext_ram_rdata2[26]
port 472 nsew signal input
rlabel metal3 s 352720 99016 353520 99136 6 data_arrays_0_ext_ram_rdata2[27]
port 473 nsew signal input
rlabel metal3 s 352720 100104 353520 100224 6 data_arrays_0_ext_ram_rdata2[28]
port 474 nsew signal input
rlabel metal3 s 352720 101192 353520 101312 6 data_arrays_0_ext_ram_rdata2[29]
port 475 nsew signal input
rlabel metal3 s 352720 71952 353520 72072 6 data_arrays_0_ext_ram_rdata2[2]
port 476 nsew signal input
rlabel metal3 s 352720 102280 353520 102400 6 data_arrays_0_ext_ram_rdata2[30]
port 477 nsew signal input
rlabel metal3 s 352720 103368 353520 103488 6 data_arrays_0_ext_ram_rdata2[31]
port 478 nsew signal input
rlabel metal3 s 352720 73040 353520 73160 6 data_arrays_0_ext_ram_rdata2[3]
port 479 nsew signal input
rlabel metal3 s 352720 74128 353520 74248 6 data_arrays_0_ext_ram_rdata2[4]
port 480 nsew signal input
rlabel metal3 s 352720 75216 353520 75336 6 data_arrays_0_ext_ram_rdata2[5]
port 481 nsew signal input
rlabel metal3 s 352720 76304 353520 76424 6 data_arrays_0_ext_ram_rdata2[6]
port 482 nsew signal input
rlabel metal3 s 352720 77392 353520 77512 6 data_arrays_0_ext_ram_rdata2[7]
port 483 nsew signal input
rlabel metal3 s 352720 78480 353520 78600 6 data_arrays_0_ext_ram_rdata2[8]
port 484 nsew signal input
rlabel metal3 s 352720 79432 353520 79552 6 data_arrays_0_ext_ram_rdata2[9]
port 485 nsew signal input
rlabel metal3 s 352720 104456 353520 104576 6 data_arrays_0_ext_ram_rdata3[0]
port 486 nsew signal input
rlabel metal3 s 352720 115336 353520 115456 6 data_arrays_0_ext_ram_rdata3[10]
port 487 nsew signal input
rlabel metal3 s 352720 116424 353520 116544 6 data_arrays_0_ext_ram_rdata3[11]
port 488 nsew signal input
rlabel metal3 s 352720 117512 353520 117632 6 data_arrays_0_ext_ram_rdata3[12]
port 489 nsew signal input
rlabel metal3 s 352720 118600 353520 118720 6 data_arrays_0_ext_ram_rdata3[13]
port 490 nsew signal input
rlabel metal3 s 352720 119552 353520 119672 6 data_arrays_0_ext_ram_rdata3[14]
port 491 nsew signal input
rlabel metal3 s 352720 120640 353520 120760 6 data_arrays_0_ext_ram_rdata3[15]
port 492 nsew signal input
rlabel metal3 s 352720 121728 353520 121848 6 data_arrays_0_ext_ram_rdata3[16]
port 493 nsew signal input
rlabel metal3 s 352720 122816 353520 122936 6 data_arrays_0_ext_ram_rdata3[17]
port 494 nsew signal input
rlabel metal3 s 352720 123904 353520 124024 6 data_arrays_0_ext_ram_rdata3[18]
port 495 nsew signal input
rlabel metal3 s 352720 124992 353520 125112 6 data_arrays_0_ext_ram_rdata3[19]
port 496 nsew signal input
rlabel metal3 s 352720 105544 353520 105664 6 data_arrays_0_ext_ram_rdata3[1]
port 497 nsew signal input
rlabel metal3 s 352720 126080 353520 126200 6 data_arrays_0_ext_ram_rdata3[20]
port 498 nsew signal input
rlabel metal3 s 352720 127168 353520 127288 6 data_arrays_0_ext_ram_rdata3[21]
port 499 nsew signal input
rlabel metal3 s 352720 128256 353520 128376 6 data_arrays_0_ext_ram_rdata3[22]
port 500 nsew signal input
rlabel metal3 s 352720 129344 353520 129464 6 data_arrays_0_ext_ram_rdata3[23]
port 501 nsew signal input
rlabel metal3 s 352720 130432 353520 130552 6 data_arrays_0_ext_ram_rdata3[24]
port 502 nsew signal input
rlabel metal3 s 352720 131520 353520 131640 6 data_arrays_0_ext_ram_rdata3[25]
port 503 nsew signal input
rlabel metal3 s 352720 132608 353520 132728 6 data_arrays_0_ext_ram_rdata3[26]
port 504 nsew signal input
rlabel metal3 s 352720 133696 353520 133816 6 data_arrays_0_ext_ram_rdata3[27]
port 505 nsew signal input
rlabel metal3 s 352720 134784 353520 134904 6 data_arrays_0_ext_ram_rdata3[28]
port 506 nsew signal input
rlabel metal3 s 352720 135872 353520 135992 6 data_arrays_0_ext_ram_rdata3[29]
port 507 nsew signal input
rlabel metal3 s 352720 106632 353520 106752 6 data_arrays_0_ext_ram_rdata3[2]
port 508 nsew signal input
rlabel metal3 s 352720 136960 353520 137080 6 data_arrays_0_ext_ram_rdata3[30]
port 509 nsew signal input
rlabel metal3 s 352720 138048 353520 138168 6 data_arrays_0_ext_ram_rdata3[31]
port 510 nsew signal input
rlabel metal3 s 352720 107720 353520 107840 6 data_arrays_0_ext_ram_rdata3[3]
port 511 nsew signal input
rlabel metal3 s 352720 108808 353520 108928 6 data_arrays_0_ext_ram_rdata3[4]
port 512 nsew signal input
rlabel metal3 s 352720 109896 353520 110016 6 data_arrays_0_ext_ram_rdata3[5]
port 513 nsew signal input
rlabel metal3 s 352720 110984 353520 111104 6 data_arrays_0_ext_ram_rdata3[6]
port 514 nsew signal input
rlabel metal3 s 352720 112072 353520 112192 6 data_arrays_0_ext_ram_rdata3[7]
port 515 nsew signal input
rlabel metal3 s 352720 113160 353520 113280 6 data_arrays_0_ext_ram_rdata3[8]
port 516 nsew signal input
rlabel metal3 s 352720 114248 353520 114368 6 data_arrays_0_ext_ram_rdata3[9]
port 517 nsew signal input
rlabel metal3 s 352720 217200 353520 217320 6 data_arrays_0_ext_ram_rdata4[0]
port 518 nsew signal input
rlabel metal3 s 352720 228080 353520 228200 6 data_arrays_0_ext_ram_rdata4[10]
port 519 nsew signal input
rlabel metal3 s 352720 229168 353520 229288 6 data_arrays_0_ext_ram_rdata4[11]
port 520 nsew signal input
rlabel metal3 s 352720 230256 353520 230376 6 data_arrays_0_ext_ram_rdata4[12]
port 521 nsew signal input
rlabel metal3 s 352720 231344 353520 231464 6 data_arrays_0_ext_ram_rdata4[13]
port 522 nsew signal input
rlabel metal3 s 352720 232432 353520 232552 6 data_arrays_0_ext_ram_rdata4[14]
port 523 nsew signal input
rlabel metal3 s 352720 233520 353520 233640 6 data_arrays_0_ext_ram_rdata4[15]
port 524 nsew signal input
rlabel metal3 s 352720 234608 353520 234728 6 data_arrays_0_ext_ram_rdata4[16]
port 525 nsew signal input
rlabel metal3 s 352720 235696 353520 235816 6 data_arrays_0_ext_ram_rdata4[17]
port 526 nsew signal input
rlabel metal3 s 352720 236784 353520 236904 6 data_arrays_0_ext_ram_rdata4[18]
port 527 nsew signal input
rlabel metal3 s 352720 237736 353520 237856 6 data_arrays_0_ext_ram_rdata4[19]
port 528 nsew signal input
rlabel metal3 s 352720 218288 353520 218408 6 data_arrays_0_ext_ram_rdata4[1]
port 529 nsew signal input
rlabel metal3 s 352720 238824 353520 238944 6 data_arrays_0_ext_ram_rdata4[20]
port 530 nsew signal input
rlabel metal3 s 352720 239912 353520 240032 6 data_arrays_0_ext_ram_rdata4[21]
port 531 nsew signal input
rlabel metal3 s 352720 241000 353520 241120 6 data_arrays_0_ext_ram_rdata4[22]
port 532 nsew signal input
rlabel metal3 s 352720 242088 353520 242208 6 data_arrays_0_ext_ram_rdata4[23]
port 533 nsew signal input
rlabel metal3 s 352720 243176 353520 243296 6 data_arrays_0_ext_ram_rdata4[24]
port 534 nsew signal input
rlabel metal3 s 352720 244264 353520 244384 6 data_arrays_0_ext_ram_rdata4[25]
port 535 nsew signal input
rlabel metal3 s 352720 245352 353520 245472 6 data_arrays_0_ext_ram_rdata4[26]
port 536 nsew signal input
rlabel metal3 s 352720 246440 353520 246560 6 data_arrays_0_ext_ram_rdata4[27]
port 537 nsew signal input
rlabel metal3 s 352720 247528 353520 247648 6 data_arrays_0_ext_ram_rdata4[28]
port 538 nsew signal input
rlabel metal3 s 352720 248616 353520 248736 6 data_arrays_0_ext_ram_rdata4[29]
port 539 nsew signal input
rlabel metal3 s 352720 219376 353520 219496 6 data_arrays_0_ext_ram_rdata4[2]
port 540 nsew signal input
rlabel metal3 s 352720 249704 353520 249824 6 data_arrays_0_ext_ram_rdata4[30]
port 541 nsew signal input
rlabel metal3 s 352720 250792 353520 250912 6 data_arrays_0_ext_ram_rdata4[31]
port 542 nsew signal input
rlabel metal3 s 352720 220464 353520 220584 6 data_arrays_0_ext_ram_rdata4[3]
port 543 nsew signal input
rlabel metal3 s 352720 221552 353520 221672 6 data_arrays_0_ext_ram_rdata4[4]
port 544 nsew signal input
rlabel metal3 s 352720 222640 353520 222760 6 data_arrays_0_ext_ram_rdata4[5]
port 545 nsew signal input
rlabel metal3 s 352720 223728 353520 223848 6 data_arrays_0_ext_ram_rdata4[6]
port 546 nsew signal input
rlabel metal3 s 352720 224816 353520 224936 6 data_arrays_0_ext_ram_rdata4[7]
port 547 nsew signal input
rlabel metal3 s 352720 225904 353520 226024 6 data_arrays_0_ext_ram_rdata4[8]
port 548 nsew signal input
rlabel metal3 s 352720 226992 353520 227112 6 data_arrays_0_ext_ram_rdata4[9]
port 549 nsew signal input
rlabel metal3 s 352720 251880 353520 252000 6 data_arrays_0_ext_ram_rdata5[0]
port 550 nsew signal input
rlabel metal3 s 352720 262760 353520 262880 6 data_arrays_0_ext_ram_rdata5[10]
port 551 nsew signal input
rlabel metal3 s 352720 263848 353520 263968 6 data_arrays_0_ext_ram_rdata5[11]
port 552 nsew signal input
rlabel metal3 s 352720 264936 353520 265056 6 data_arrays_0_ext_ram_rdata5[12]
port 553 nsew signal input
rlabel metal3 s 352720 266024 353520 266144 6 data_arrays_0_ext_ram_rdata5[13]
port 554 nsew signal input
rlabel metal3 s 352720 267112 353520 267232 6 data_arrays_0_ext_ram_rdata5[14]
port 555 nsew signal input
rlabel metal3 s 352720 268200 353520 268320 6 data_arrays_0_ext_ram_rdata5[15]
port 556 nsew signal input
rlabel metal3 s 352720 269288 353520 269408 6 data_arrays_0_ext_ram_rdata5[16]
port 557 nsew signal input
rlabel metal3 s 352720 270376 353520 270496 6 data_arrays_0_ext_ram_rdata5[17]
port 558 nsew signal input
rlabel metal3 s 352720 271464 353520 271584 6 data_arrays_0_ext_ram_rdata5[18]
port 559 nsew signal input
rlabel metal3 s 352720 272552 353520 272672 6 data_arrays_0_ext_ram_rdata5[19]
port 560 nsew signal input
rlabel metal3 s 352720 252968 353520 253088 6 data_arrays_0_ext_ram_rdata5[1]
port 561 nsew signal input
rlabel metal3 s 352720 273640 353520 273760 6 data_arrays_0_ext_ram_rdata5[20]
port 562 nsew signal input
rlabel metal3 s 352720 274728 353520 274848 6 data_arrays_0_ext_ram_rdata5[21]
port 563 nsew signal input
rlabel metal3 s 352720 275816 353520 275936 6 data_arrays_0_ext_ram_rdata5[22]
port 564 nsew signal input
rlabel metal3 s 352720 276904 353520 277024 6 data_arrays_0_ext_ram_rdata5[23]
port 565 nsew signal input
rlabel metal3 s 352720 277856 353520 277976 6 data_arrays_0_ext_ram_rdata5[24]
port 566 nsew signal input
rlabel metal3 s 352720 278944 353520 279064 6 data_arrays_0_ext_ram_rdata5[25]
port 567 nsew signal input
rlabel metal3 s 352720 280032 353520 280152 6 data_arrays_0_ext_ram_rdata5[26]
port 568 nsew signal input
rlabel metal3 s 352720 281120 353520 281240 6 data_arrays_0_ext_ram_rdata5[27]
port 569 nsew signal input
rlabel metal3 s 352720 282208 353520 282328 6 data_arrays_0_ext_ram_rdata5[28]
port 570 nsew signal input
rlabel metal3 s 352720 283296 353520 283416 6 data_arrays_0_ext_ram_rdata5[29]
port 571 nsew signal input
rlabel metal3 s 352720 254056 353520 254176 6 data_arrays_0_ext_ram_rdata5[2]
port 572 nsew signal input
rlabel metal3 s 352720 284384 353520 284504 6 data_arrays_0_ext_ram_rdata5[30]
port 573 nsew signal input
rlabel metal3 s 352720 285472 353520 285592 6 data_arrays_0_ext_ram_rdata5[31]
port 574 nsew signal input
rlabel metal3 s 352720 255144 353520 255264 6 data_arrays_0_ext_ram_rdata5[3]
port 575 nsew signal input
rlabel metal3 s 352720 256232 353520 256352 6 data_arrays_0_ext_ram_rdata5[4]
port 576 nsew signal input
rlabel metal3 s 352720 257320 353520 257440 6 data_arrays_0_ext_ram_rdata5[5]
port 577 nsew signal input
rlabel metal3 s 352720 258408 353520 258528 6 data_arrays_0_ext_ram_rdata5[6]
port 578 nsew signal input
rlabel metal3 s 352720 259496 353520 259616 6 data_arrays_0_ext_ram_rdata5[7]
port 579 nsew signal input
rlabel metal3 s 352720 260584 353520 260704 6 data_arrays_0_ext_ram_rdata5[8]
port 580 nsew signal input
rlabel metal3 s 352720 261672 353520 261792 6 data_arrays_0_ext_ram_rdata5[9]
port 581 nsew signal input
rlabel metal3 s 352720 286560 353520 286680 6 data_arrays_0_ext_ram_rdata6[0]
port 582 nsew signal input
rlabel metal3 s 352720 297440 353520 297560 6 data_arrays_0_ext_ram_rdata6[10]
port 583 nsew signal input
rlabel metal3 s 352720 298528 353520 298648 6 data_arrays_0_ext_ram_rdata6[11]
port 584 nsew signal input
rlabel metal3 s 352720 299616 353520 299736 6 data_arrays_0_ext_ram_rdata6[12]
port 585 nsew signal input
rlabel metal3 s 352720 300704 353520 300824 6 data_arrays_0_ext_ram_rdata6[13]
port 586 nsew signal input
rlabel metal3 s 352720 301792 353520 301912 6 data_arrays_0_ext_ram_rdata6[14]
port 587 nsew signal input
rlabel metal3 s 352720 302880 353520 303000 6 data_arrays_0_ext_ram_rdata6[15]
port 588 nsew signal input
rlabel metal3 s 352720 303968 353520 304088 6 data_arrays_0_ext_ram_rdata6[16]
port 589 nsew signal input
rlabel metal3 s 352720 305056 353520 305176 6 data_arrays_0_ext_ram_rdata6[17]
port 590 nsew signal input
rlabel metal3 s 352720 306144 353520 306264 6 data_arrays_0_ext_ram_rdata6[18]
port 591 nsew signal input
rlabel metal3 s 352720 307232 353520 307352 6 data_arrays_0_ext_ram_rdata6[19]
port 592 nsew signal input
rlabel metal3 s 352720 287648 353520 287768 6 data_arrays_0_ext_ram_rdata6[1]
port 593 nsew signal input
rlabel metal3 s 352720 308320 353520 308440 6 data_arrays_0_ext_ram_rdata6[20]
port 594 nsew signal input
rlabel metal3 s 352720 309408 353520 309528 6 data_arrays_0_ext_ram_rdata6[21]
port 595 nsew signal input
rlabel metal3 s 352720 310496 353520 310616 6 data_arrays_0_ext_ram_rdata6[22]
port 596 nsew signal input
rlabel metal3 s 352720 311584 353520 311704 6 data_arrays_0_ext_ram_rdata6[23]
port 597 nsew signal input
rlabel metal3 s 352720 312672 353520 312792 6 data_arrays_0_ext_ram_rdata6[24]
port 598 nsew signal input
rlabel metal3 s 352720 313760 353520 313880 6 data_arrays_0_ext_ram_rdata6[25]
port 599 nsew signal input
rlabel metal3 s 352720 314848 353520 314968 6 data_arrays_0_ext_ram_rdata6[26]
port 600 nsew signal input
rlabel metal3 s 352720 315936 353520 316056 6 data_arrays_0_ext_ram_rdata6[27]
port 601 nsew signal input
rlabel metal3 s 352720 316888 353520 317008 6 data_arrays_0_ext_ram_rdata6[28]
port 602 nsew signal input
rlabel metal3 s 352720 317976 353520 318096 6 data_arrays_0_ext_ram_rdata6[29]
port 603 nsew signal input
rlabel metal3 s 352720 288736 353520 288856 6 data_arrays_0_ext_ram_rdata6[2]
port 604 nsew signal input
rlabel metal3 s 352720 319064 353520 319184 6 data_arrays_0_ext_ram_rdata6[30]
port 605 nsew signal input
rlabel metal3 s 352720 320152 353520 320272 6 data_arrays_0_ext_ram_rdata6[31]
port 606 nsew signal input
rlabel metal3 s 352720 289824 353520 289944 6 data_arrays_0_ext_ram_rdata6[3]
port 607 nsew signal input
rlabel metal3 s 352720 290912 353520 291032 6 data_arrays_0_ext_ram_rdata6[4]
port 608 nsew signal input
rlabel metal3 s 352720 292000 353520 292120 6 data_arrays_0_ext_ram_rdata6[5]
port 609 nsew signal input
rlabel metal3 s 352720 293088 353520 293208 6 data_arrays_0_ext_ram_rdata6[6]
port 610 nsew signal input
rlabel metal3 s 352720 294176 353520 294296 6 data_arrays_0_ext_ram_rdata6[7]
port 611 nsew signal input
rlabel metal3 s 352720 295264 353520 295384 6 data_arrays_0_ext_ram_rdata6[8]
port 612 nsew signal input
rlabel metal3 s 352720 296352 353520 296472 6 data_arrays_0_ext_ram_rdata6[9]
port 613 nsew signal input
rlabel metal3 s 352720 321240 353520 321360 6 data_arrays_0_ext_ram_rdata7[0]
port 614 nsew signal input
rlabel metal3 s 352720 332120 353520 332240 6 data_arrays_0_ext_ram_rdata7[10]
port 615 nsew signal input
rlabel metal3 s 352720 333208 353520 333328 6 data_arrays_0_ext_ram_rdata7[11]
port 616 nsew signal input
rlabel metal3 s 352720 334296 353520 334416 6 data_arrays_0_ext_ram_rdata7[12]
port 617 nsew signal input
rlabel metal3 s 352720 335384 353520 335504 6 data_arrays_0_ext_ram_rdata7[13]
port 618 nsew signal input
rlabel metal3 s 352720 336472 353520 336592 6 data_arrays_0_ext_ram_rdata7[14]
port 619 nsew signal input
rlabel metal3 s 352720 337560 353520 337680 6 data_arrays_0_ext_ram_rdata7[15]
port 620 nsew signal input
rlabel metal3 s 352720 338648 353520 338768 6 data_arrays_0_ext_ram_rdata7[16]
port 621 nsew signal input
rlabel metal3 s 352720 339736 353520 339856 6 data_arrays_0_ext_ram_rdata7[17]
port 622 nsew signal input
rlabel metal3 s 352720 340824 353520 340944 6 data_arrays_0_ext_ram_rdata7[18]
port 623 nsew signal input
rlabel metal3 s 352720 341912 353520 342032 6 data_arrays_0_ext_ram_rdata7[19]
port 624 nsew signal input
rlabel metal3 s 352720 322328 353520 322448 6 data_arrays_0_ext_ram_rdata7[1]
port 625 nsew signal input
rlabel metal3 s 352720 343000 353520 343120 6 data_arrays_0_ext_ram_rdata7[20]
port 626 nsew signal input
rlabel metal3 s 352720 344088 353520 344208 6 data_arrays_0_ext_ram_rdata7[21]
port 627 nsew signal input
rlabel metal3 s 352720 345176 353520 345296 6 data_arrays_0_ext_ram_rdata7[22]
port 628 nsew signal input
rlabel metal3 s 352720 346264 353520 346384 6 data_arrays_0_ext_ram_rdata7[23]
port 629 nsew signal input
rlabel metal3 s 352720 347352 353520 347472 6 data_arrays_0_ext_ram_rdata7[24]
port 630 nsew signal input
rlabel metal3 s 352720 348440 353520 348560 6 data_arrays_0_ext_ram_rdata7[25]
port 631 nsew signal input
rlabel metal3 s 352720 349528 353520 349648 6 data_arrays_0_ext_ram_rdata7[26]
port 632 nsew signal input
rlabel metal3 s 352720 350616 353520 350736 6 data_arrays_0_ext_ram_rdata7[27]
port 633 nsew signal input
rlabel metal3 s 352720 351704 353520 351824 6 data_arrays_0_ext_ram_rdata7[28]
port 634 nsew signal input
rlabel metal3 s 352720 352792 353520 352912 6 data_arrays_0_ext_ram_rdata7[29]
port 635 nsew signal input
rlabel metal3 s 352720 323416 353520 323536 6 data_arrays_0_ext_ram_rdata7[2]
port 636 nsew signal input
rlabel metal3 s 352720 353880 353520 354000 6 data_arrays_0_ext_ram_rdata7[30]
port 637 nsew signal input
rlabel metal3 s 352720 354968 353520 355088 6 data_arrays_0_ext_ram_rdata7[31]
port 638 nsew signal input
rlabel metal3 s 352720 324504 353520 324624 6 data_arrays_0_ext_ram_rdata7[3]
port 639 nsew signal input
rlabel metal3 s 352720 325592 353520 325712 6 data_arrays_0_ext_ram_rdata7[4]
port 640 nsew signal input
rlabel metal3 s 352720 326680 353520 326800 6 data_arrays_0_ext_ram_rdata7[5]
port 641 nsew signal input
rlabel metal3 s 352720 327768 353520 327888 6 data_arrays_0_ext_ram_rdata7[6]
port 642 nsew signal input
rlabel metal3 s 352720 328856 353520 328976 6 data_arrays_0_ext_ram_rdata7[7]
port 643 nsew signal input
rlabel metal3 s 352720 329944 353520 330064 6 data_arrays_0_ext_ram_rdata7[8]
port 644 nsew signal input
rlabel metal3 s 352720 331032 353520 331152 6 data_arrays_0_ext_ram_rdata7[9]
port 645 nsew signal input
rlabel metal3 s 352720 150016 353520 150136 6 data_arrays_0_ext_ram_wdata[0]
port 646 nsew signal output
rlabel metal3 s 352720 160760 353520 160880 6 data_arrays_0_ext_ram_wdata[10]
port 647 nsew signal output
rlabel metal3 s 352720 161848 353520 161968 6 data_arrays_0_ext_ram_wdata[11]
port 648 nsew signal output
rlabel metal3 s 352720 162936 353520 163056 6 data_arrays_0_ext_ram_wdata[12]
port 649 nsew signal output
rlabel metal3 s 352720 164024 353520 164144 6 data_arrays_0_ext_ram_wdata[13]
port 650 nsew signal output
rlabel metal3 s 352720 165112 353520 165232 6 data_arrays_0_ext_ram_wdata[14]
port 651 nsew signal output
rlabel metal3 s 352720 166200 353520 166320 6 data_arrays_0_ext_ram_wdata[15]
port 652 nsew signal output
rlabel metal3 s 352720 167288 353520 167408 6 data_arrays_0_ext_ram_wdata[16]
port 653 nsew signal output
rlabel metal3 s 352720 168376 353520 168496 6 data_arrays_0_ext_ram_wdata[17]
port 654 nsew signal output
rlabel metal3 s 352720 169464 353520 169584 6 data_arrays_0_ext_ram_wdata[18]
port 655 nsew signal output
rlabel metal3 s 352720 170552 353520 170672 6 data_arrays_0_ext_ram_wdata[19]
port 656 nsew signal output
rlabel metal3 s 352720 151104 353520 151224 6 data_arrays_0_ext_ram_wdata[1]
port 657 nsew signal output
rlabel metal3 s 352720 171640 353520 171760 6 data_arrays_0_ext_ram_wdata[20]
port 658 nsew signal output
rlabel metal3 s 352720 172728 353520 172848 6 data_arrays_0_ext_ram_wdata[21]
port 659 nsew signal output
rlabel metal3 s 352720 173816 353520 173936 6 data_arrays_0_ext_ram_wdata[22]
port 660 nsew signal output
rlabel metal3 s 352720 174904 353520 175024 6 data_arrays_0_ext_ram_wdata[23]
port 661 nsew signal output
rlabel metal3 s 352720 175992 353520 176112 6 data_arrays_0_ext_ram_wdata[24]
port 662 nsew signal output
rlabel metal3 s 352720 177080 353520 177200 6 data_arrays_0_ext_ram_wdata[25]
port 663 nsew signal output
rlabel metal3 s 352720 178168 353520 178288 6 data_arrays_0_ext_ram_wdata[26]
port 664 nsew signal output
rlabel metal3 s 352720 179256 353520 179376 6 data_arrays_0_ext_ram_wdata[27]
port 665 nsew signal output
rlabel metal3 s 352720 180344 353520 180464 6 data_arrays_0_ext_ram_wdata[28]
port 666 nsew signal output
rlabel metal3 s 352720 181432 353520 181552 6 data_arrays_0_ext_ram_wdata[29]
port 667 nsew signal output
rlabel metal3 s 352720 152192 353520 152312 6 data_arrays_0_ext_ram_wdata[2]
port 668 nsew signal output
rlabel metal3 s 352720 182520 353520 182640 6 data_arrays_0_ext_ram_wdata[30]
port 669 nsew signal output
rlabel metal3 s 352720 183608 353520 183728 6 data_arrays_0_ext_ram_wdata[31]
port 670 nsew signal output
rlabel metal3 s 352720 153280 353520 153400 6 data_arrays_0_ext_ram_wdata[3]
port 671 nsew signal output
rlabel metal3 s 352720 154368 353520 154488 6 data_arrays_0_ext_ram_wdata[4]
port 672 nsew signal output
rlabel metal3 s 352720 155456 353520 155576 6 data_arrays_0_ext_ram_wdata[5]
port 673 nsew signal output
rlabel metal3 s 352720 156544 353520 156664 6 data_arrays_0_ext_ram_wdata[6]
port 674 nsew signal output
rlabel metal3 s 352720 157632 353520 157752 6 data_arrays_0_ext_ram_wdata[7]
port 675 nsew signal output
rlabel metal3 s 352720 158584 353520 158704 6 data_arrays_0_ext_ram_wdata[8]
port 676 nsew signal output
rlabel metal3 s 352720 159672 353520 159792 6 data_arrays_0_ext_ram_wdata[9]
port 677 nsew signal output
rlabel metal3 s 352720 197752 353520 197872 6 data_arrays_0_ext_ram_web
port 678 nsew signal output
rlabel metal3 s 352720 184696 353520 184816 6 data_arrays_0_ext_ram_wmask[0]
port 679 nsew signal output
rlabel metal3 s 352720 185784 353520 185904 6 data_arrays_0_ext_ram_wmask[1]
port 680 nsew signal output
rlabel metal3 s 352720 186872 353520 186992 6 data_arrays_0_ext_ram_wmask[2]
port 681 nsew signal output
rlabel metal3 s 352720 187960 353520 188080 6 data_arrays_0_ext_ram_wmask[3]
port 682 nsew signal output
rlabel metal2 s 1490 354864 1546 355664 6 io_in[0]
port 683 nsew signal input
rlabel metal2 s 94502 354864 94558 355664 6 io_in[10]
port 684 nsew signal input
rlabel metal2 s 103794 354864 103850 355664 6 io_in[11]
port 685 nsew signal input
rlabel metal2 s 113086 354864 113142 355664 6 io_in[12]
port 686 nsew signal input
rlabel metal2 s 122378 354864 122434 355664 6 io_in[13]
port 687 nsew signal input
rlabel metal2 s 131670 354864 131726 355664 6 io_in[14]
port 688 nsew signal input
rlabel metal2 s 140962 354864 141018 355664 6 io_in[15]
port 689 nsew signal input
rlabel metal2 s 150346 354864 150402 355664 6 io_in[16]
port 690 nsew signal input
rlabel metal2 s 159638 354864 159694 355664 6 io_in[17]
port 691 nsew signal input
rlabel metal2 s 168930 354864 168986 355664 6 io_in[18]
port 692 nsew signal input
rlabel metal2 s 178222 354864 178278 355664 6 io_in[19]
port 693 nsew signal input
rlabel metal2 s 10782 354864 10838 355664 6 io_in[1]
port 694 nsew signal input
rlabel metal2 s 187514 354864 187570 355664 6 io_in[20]
port 695 nsew signal input
rlabel metal2 s 196806 354864 196862 355664 6 io_in[21]
port 696 nsew signal input
rlabel metal2 s 206098 354864 206154 355664 6 io_in[22]
port 697 nsew signal input
rlabel metal2 s 215482 354864 215538 355664 6 io_in[23]
port 698 nsew signal input
rlabel metal2 s 224774 354864 224830 355664 6 io_in[24]
port 699 nsew signal input
rlabel metal2 s 234066 354864 234122 355664 6 io_in[25]
port 700 nsew signal input
rlabel metal2 s 243358 354864 243414 355664 6 io_in[26]
port 701 nsew signal input
rlabel metal2 s 252650 354864 252706 355664 6 io_in[27]
port 702 nsew signal input
rlabel metal2 s 261942 354864 261998 355664 6 io_in[28]
port 703 nsew signal input
rlabel metal2 s 271234 354864 271290 355664 6 io_in[29]
port 704 nsew signal input
rlabel metal2 s 20074 354864 20130 355664 6 io_in[2]
port 705 nsew signal input
rlabel metal2 s 280526 354864 280582 355664 6 io_in[30]
port 706 nsew signal input
rlabel metal2 s 289910 354864 289966 355664 6 io_in[31]
port 707 nsew signal input
rlabel metal2 s 299202 354864 299258 355664 6 io_in[32]
port 708 nsew signal input
rlabel metal2 s 308494 354864 308550 355664 6 io_in[33]
port 709 nsew signal input
rlabel metal2 s 317786 354864 317842 355664 6 io_in[34]
port 710 nsew signal input
rlabel metal2 s 327078 354864 327134 355664 6 io_in[35]
port 711 nsew signal input
rlabel metal2 s 336370 354864 336426 355664 6 io_in[36]
port 712 nsew signal input
rlabel metal2 s 345662 354864 345718 355664 6 io_in[37]
port 713 nsew signal input
rlabel metal2 s 29366 354864 29422 355664 6 io_in[3]
port 714 nsew signal input
rlabel metal2 s 38658 354864 38714 355664 6 io_in[4]
port 715 nsew signal input
rlabel metal2 s 47950 354864 48006 355664 6 io_in[5]
port 716 nsew signal input
rlabel metal2 s 57242 354864 57298 355664 6 io_in[6]
port 717 nsew signal input
rlabel metal2 s 66534 354864 66590 355664 6 io_in[7]
port 718 nsew signal input
rlabel metal2 s 75918 354864 75974 355664 6 io_in[8]
port 719 nsew signal input
rlabel metal2 s 85210 354864 85266 355664 6 io_in[9]
port 720 nsew signal input
rlabel metal2 s 4526 354864 4582 355664 6 io_oeb[0]
port 721 nsew signal output
rlabel metal2 s 97630 354864 97686 355664 6 io_oeb[10]
port 722 nsew signal output
rlabel metal2 s 106922 354864 106978 355664 6 io_oeb[11]
port 723 nsew signal output
rlabel metal2 s 116214 354864 116270 355664 6 io_oeb[12]
port 724 nsew signal output
rlabel metal2 s 125506 354864 125562 355664 6 io_oeb[13]
port 725 nsew signal output
rlabel metal2 s 134798 354864 134854 355664 6 io_oeb[14]
port 726 nsew signal output
rlabel metal2 s 144090 354864 144146 355664 6 io_oeb[15]
port 727 nsew signal output
rlabel metal2 s 153382 354864 153438 355664 6 io_oeb[16]
port 728 nsew signal output
rlabel metal2 s 162674 354864 162730 355664 6 io_oeb[17]
port 729 nsew signal output
rlabel metal2 s 172058 354864 172114 355664 6 io_oeb[18]
port 730 nsew signal output
rlabel metal2 s 181350 354864 181406 355664 6 io_oeb[19]
port 731 nsew signal output
rlabel metal2 s 13818 354864 13874 355664 6 io_oeb[1]
port 732 nsew signal output
rlabel metal2 s 190642 354864 190698 355664 6 io_oeb[20]
port 733 nsew signal output
rlabel metal2 s 199934 354864 199990 355664 6 io_oeb[21]
port 734 nsew signal output
rlabel metal2 s 209226 354864 209282 355664 6 io_oeb[22]
port 735 nsew signal output
rlabel metal2 s 218518 354864 218574 355664 6 io_oeb[23]
port 736 nsew signal output
rlabel metal2 s 227810 354864 227866 355664 6 io_oeb[24]
port 737 nsew signal output
rlabel metal2 s 237194 354864 237250 355664 6 io_oeb[25]
port 738 nsew signal output
rlabel metal2 s 246486 354864 246542 355664 6 io_oeb[26]
port 739 nsew signal output
rlabel metal2 s 255778 354864 255834 355664 6 io_oeb[27]
port 740 nsew signal output
rlabel metal2 s 265070 354864 265126 355664 6 io_oeb[28]
port 741 nsew signal output
rlabel metal2 s 274362 354864 274418 355664 6 io_oeb[29]
port 742 nsew signal output
rlabel metal2 s 23110 354864 23166 355664 6 io_oeb[2]
port 743 nsew signal output
rlabel metal2 s 283654 354864 283710 355664 6 io_oeb[30]
port 744 nsew signal output
rlabel metal2 s 292946 354864 293002 355664 6 io_oeb[31]
port 745 nsew signal output
rlabel metal2 s 302238 354864 302294 355664 6 io_oeb[32]
port 746 nsew signal output
rlabel metal2 s 311622 354864 311678 355664 6 io_oeb[33]
port 747 nsew signal output
rlabel metal2 s 320914 354864 320970 355664 6 io_oeb[34]
port 748 nsew signal output
rlabel metal2 s 330206 354864 330262 355664 6 io_oeb[35]
port 749 nsew signal output
rlabel metal2 s 339498 354864 339554 355664 6 io_oeb[36]
port 750 nsew signal output
rlabel metal2 s 348790 354864 348846 355664 6 io_oeb[37]
port 751 nsew signal output
rlabel metal2 s 32494 354864 32550 355664 6 io_oeb[3]
port 752 nsew signal output
rlabel metal2 s 41786 354864 41842 355664 6 io_oeb[4]
port 753 nsew signal output
rlabel metal2 s 51078 354864 51134 355664 6 io_oeb[5]
port 754 nsew signal output
rlabel metal2 s 60370 354864 60426 355664 6 io_oeb[6]
port 755 nsew signal output
rlabel metal2 s 69662 354864 69718 355664 6 io_oeb[7]
port 756 nsew signal output
rlabel metal2 s 78954 354864 79010 355664 6 io_oeb[8]
port 757 nsew signal output
rlabel metal2 s 88246 354864 88302 355664 6 io_oeb[9]
port 758 nsew signal output
rlabel metal2 s 7654 354864 7710 355664 6 io_out[0]
port 759 nsew signal output
rlabel metal2 s 100666 354864 100722 355664 6 io_out[10]
port 760 nsew signal output
rlabel metal2 s 109958 354864 110014 355664 6 io_out[11]
port 761 nsew signal output
rlabel metal2 s 119342 354864 119398 355664 6 io_out[12]
port 762 nsew signal output
rlabel metal2 s 128634 354864 128690 355664 6 io_out[13]
port 763 nsew signal output
rlabel metal2 s 137926 354864 137982 355664 6 io_out[14]
port 764 nsew signal output
rlabel metal2 s 147218 354864 147274 355664 6 io_out[15]
port 765 nsew signal output
rlabel metal2 s 156510 354864 156566 355664 6 io_out[16]
port 766 nsew signal output
rlabel metal2 s 165802 354864 165858 355664 6 io_out[17]
port 767 nsew signal output
rlabel metal2 s 175094 354864 175150 355664 6 io_out[18]
port 768 nsew signal output
rlabel metal2 s 184386 354864 184442 355664 6 io_out[19]
port 769 nsew signal output
rlabel metal2 s 16946 354864 17002 355664 6 io_out[1]
port 770 nsew signal output
rlabel metal2 s 193770 354864 193826 355664 6 io_out[20]
port 771 nsew signal output
rlabel metal2 s 203062 354864 203118 355664 6 io_out[21]
port 772 nsew signal output
rlabel metal2 s 212354 354864 212410 355664 6 io_out[22]
port 773 nsew signal output
rlabel metal2 s 221646 354864 221702 355664 6 io_out[23]
port 774 nsew signal output
rlabel metal2 s 230938 354864 230994 355664 6 io_out[24]
port 775 nsew signal output
rlabel metal2 s 240230 354864 240286 355664 6 io_out[25]
port 776 nsew signal output
rlabel metal2 s 249522 354864 249578 355664 6 io_out[26]
port 777 nsew signal output
rlabel metal2 s 258814 354864 258870 355664 6 io_out[27]
port 778 nsew signal output
rlabel metal2 s 268198 354864 268254 355664 6 io_out[28]
port 779 nsew signal output
rlabel metal2 s 277490 354864 277546 355664 6 io_out[29]
port 780 nsew signal output
rlabel metal2 s 26238 354864 26294 355664 6 io_out[2]
port 781 nsew signal output
rlabel metal2 s 286782 354864 286838 355664 6 io_out[30]
port 782 nsew signal output
rlabel metal2 s 296074 354864 296130 355664 6 io_out[31]
port 783 nsew signal output
rlabel metal2 s 305366 354864 305422 355664 6 io_out[32]
port 784 nsew signal output
rlabel metal2 s 314658 354864 314714 355664 6 io_out[33]
port 785 nsew signal output
rlabel metal2 s 323950 354864 324006 355664 6 io_out[34]
port 786 nsew signal output
rlabel metal2 s 333334 354864 333390 355664 6 io_out[35]
port 787 nsew signal output
rlabel metal2 s 342626 354864 342682 355664 6 io_out[36]
port 788 nsew signal output
rlabel metal2 s 351918 354864 351974 355664 6 io_out[37]
port 789 nsew signal output
rlabel metal2 s 35530 354864 35586 355664 6 io_out[3]
port 790 nsew signal output
rlabel metal2 s 44822 354864 44878 355664 6 io_out[4]
port 791 nsew signal output
rlabel metal2 s 54206 354864 54262 355664 6 io_out[5]
port 792 nsew signal output
rlabel metal2 s 63498 354864 63554 355664 6 io_out[6]
port 793 nsew signal output
rlabel metal2 s 72790 354864 72846 355664 6 io_out[7]
port 794 nsew signal output
rlabel metal2 s 82082 354864 82138 355664 6 io_out[8]
port 795 nsew signal output
rlabel metal2 s 91374 354864 91430 355664 6 io_out[9]
port 796 nsew signal output
rlabel metal2 s 351642 0 351698 800 6 irq[0]
port 797 nsew signal output
rlabel metal2 s 352378 0 352434 800 6 irq[1]
port 798 nsew signal output
rlabel metal2 s 353114 0 353170 800 6 irq[2]
port 799 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 la_data_in[0]
port 800 nsew signal input
rlabel metal2 s 291382 0 291438 800 6 la_data_in[100]
port 801 nsew signal input
rlabel metal2 s 293590 0 293646 800 6 la_data_in[101]
port 802 nsew signal input
rlabel metal2 s 295706 0 295762 800 6 la_data_in[102]
port 803 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_data_in[103]
port 804 nsew signal input
rlabel metal2 s 300030 0 300086 800 6 la_data_in[104]
port 805 nsew signal input
rlabel metal2 s 302146 0 302202 800 6 la_data_in[105]
port 806 nsew signal input
rlabel metal2 s 304354 0 304410 800 6 la_data_in[106]
port 807 nsew signal input
rlabel metal2 s 306470 0 306526 800 6 la_data_in[107]
port 808 nsew signal input
rlabel metal2 s 308586 0 308642 800 6 la_data_in[108]
port 809 nsew signal input
rlabel metal2 s 310794 0 310850 800 6 la_data_in[109]
port 810 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[10]
port 811 nsew signal input
rlabel metal2 s 312910 0 312966 800 6 la_data_in[110]
port 812 nsew signal input
rlabel metal2 s 315118 0 315174 800 6 la_data_in[111]
port 813 nsew signal input
rlabel metal2 s 317234 0 317290 800 6 la_data_in[112]
port 814 nsew signal input
rlabel metal2 s 319350 0 319406 800 6 la_data_in[113]
port 815 nsew signal input
rlabel metal2 s 321558 0 321614 800 6 la_data_in[114]
port 816 nsew signal input
rlabel metal2 s 323674 0 323730 800 6 la_data_in[115]
port 817 nsew signal input
rlabel metal2 s 325790 0 325846 800 6 la_data_in[116]
port 818 nsew signal input
rlabel metal2 s 327998 0 328054 800 6 la_data_in[117]
port 819 nsew signal input
rlabel metal2 s 330114 0 330170 800 6 la_data_in[118]
port 820 nsew signal input
rlabel metal2 s 332322 0 332378 800 6 la_data_in[119]
port 821 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[11]
port 822 nsew signal input
rlabel metal2 s 334438 0 334494 800 6 la_data_in[120]
port 823 nsew signal input
rlabel metal2 s 336554 0 336610 800 6 la_data_in[121]
port 824 nsew signal input
rlabel metal2 s 338762 0 338818 800 6 la_data_in[122]
port 825 nsew signal input
rlabel metal2 s 340878 0 340934 800 6 la_data_in[123]
port 826 nsew signal input
rlabel metal2 s 343086 0 343142 800 6 la_data_in[124]
port 827 nsew signal input
rlabel metal2 s 345202 0 345258 800 6 la_data_in[125]
port 828 nsew signal input
rlabel metal2 s 347318 0 347374 800 6 la_data_in[126]
port 829 nsew signal input
rlabel metal2 s 349526 0 349582 800 6 la_data_in[127]
port 830 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[12]
port 831 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[13]
port 832 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_data_in[14]
port 833 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_data_in[15]
port 834 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[16]
port 835 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[17]
port 836 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_data_in[18]
port 837 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[19]
port 838 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[1]
port 839 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[20]
port 840 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[21]
port 841 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_data_in[22]
port 842 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_data_in[23]
port 843 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_data_in[24]
port 844 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[25]
port 845 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[26]
port 846 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[27]
port 847 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[28]
port 848 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_data_in[29]
port 849 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[2]
port 850 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[30]
port 851 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[31]
port 852 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[32]
port 853 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_data_in[33]
port 854 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[34]
port 855 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_data_in[35]
port 856 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_data_in[36]
port 857 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_data_in[37]
port 858 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[38]
port 859 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_data_in[39]
port 860 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[3]
port 861 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_data_in[40]
port 862 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_data_in[41]
port 863 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_data_in[42]
port 864 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[43]
port 865 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[44]
port 866 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 la_data_in[45]
port 867 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_data_in[46]
port 868 nsew signal input
rlabel metal2 s 177394 0 177450 800 6 la_data_in[47]
port 869 nsew signal input
rlabel metal2 s 179510 0 179566 800 6 la_data_in[48]
port 870 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_data_in[49]
port 871 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[4]
port 872 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_data_in[50]
port 873 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_data_in[51]
port 874 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_data_in[52]
port 875 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[53]
port 876 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 la_data_in[54]
port 877 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 la_data_in[55]
port 878 nsew signal input
rlabel metal2 s 196714 0 196770 800 6 la_data_in[56]
port 879 nsew signal input
rlabel metal2 s 198922 0 198978 800 6 la_data_in[57]
port 880 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_data_in[58]
port 881 nsew signal input
rlabel metal2 s 203246 0 203302 800 6 la_data_in[59]
port 882 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[5]
port 883 nsew signal input
rlabel metal2 s 205362 0 205418 800 6 la_data_in[60]
port 884 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_data_in[61]
port 885 nsew signal input
rlabel metal2 s 209686 0 209742 800 6 la_data_in[62]
port 886 nsew signal input
rlabel metal2 s 211802 0 211858 800 6 la_data_in[63]
port 887 nsew signal input
rlabel metal2 s 213918 0 213974 800 6 la_data_in[64]
port 888 nsew signal input
rlabel metal2 s 216126 0 216182 800 6 la_data_in[65]
port 889 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_data_in[66]
port 890 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_data_in[67]
port 891 nsew signal input
rlabel metal2 s 222566 0 222622 800 6 la_data_in[68]
port 892 nsew signal input
rlabel metal2 s 224682 0 224738 800 6 la_data_in[69]
port 893 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[6]
port 894 nsew signal input
rlabel metal2 s 226890 0 226946 800 6 la_data_in[70]
port 895 nsew signal input
rlabel metal2 s 229006 0 229062 800 6 la_data_in[71]
port 896 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 la_data_in[72]
port 897 nsew signal input
rlabel metal2 s 233330 0 233386 800 6 la_data_in[73]
port 898 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_data_in[74]
port 899 nsew signal input
rlabel metal2 s 237654 0 237710 800 6 la_data_in[75]
port 900 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_data_in[76]
port 901 nsew signal input
rlabel metal2 s 241886 0 241942 800 6 la_data_in[77]
port 902 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 la_data_in[78]
port 903 nsew signal input
rlabel metal2 s 246210 0 246266 800 6 la_data_in[79]
port 904 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_data_in[7]
port 905 nsew signal input
rlabel metal2 s 248418 0 248474 800 6 la_data_in[80]
port 906 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_data_in[81]
port 907 nsew signal input
rlabel metal2 s 252650 0 252706 800 6 la_data_in[82]
port 908 nsew signal input
rlabel metal2 s 254858 0 254914 800 6 la_data_in[83]
port 909 nsew signal input
rlabel metal2 s 256974 0 257030 800 6 la_data_in[84]
port 910 nsew signal input
rlabel metal2 s 259182 0 259238 800 6 la_data_in[85]
port 911 nsew signal input
rlabel metal2 s 261298 0 261354 800 6 la_data_in[86]
port 912 nsew signal input
rlabel metal2 s 263414 0 263470 800 6 la_data_in[87]
port 913 nsew signal input
rlabel metal2 s 265622 0 265678 800 6 la_data_in[88]
port 914 nsew signal input
rlabel metal2 s 267738 0 267794 800 6 la_data_in[89]
port 915 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[8]
port 916 nsew signal input
rlabel metal2 s 269854 0 269910 800 6 la_data_in[90]
port 917 nsew signal input
rlabel metal2 s 272062 0 272118 800 6 la_data_in[91]
port 918 nsew signal input
rlabel metal2 s 274178 0 274234 800 6 la_data_in[92]
port 919 nsew signal input
rlabel metal2 s 276386 0 276442 800 6 la_data_in[93]
port 920 nsew signal input
rlabel metal2 s 278502 0 278558 800 6 la_data_in[94]
port 921 nsew signal input
rlabel metal2 s 280618 0 280674 800 6 la_data_in[95]
port 922 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_data_in[96]
port 923 nsew signal input
rlabel metal2 s 284942 0 284998 800 6 la_data_in[97]
port 924 nsew signal input
rlabel metal2 s 287150 0 287206 800 6 la_data_in[98]
port 925 nsew signal input
rlabel metal2 s 289266 0 289322 800 6 la_data_in[99]
port 926 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[9]
port 927 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_data_out[0]
port 928 nsew signal output
rlabel metal2 s 292118 0 292174 800 6 la_data_out[100]
port 929 nsew signal output
rlabel metal2 s 294326 0 294382 800 6 la_data_out[101]
port 930 nsew signal output
rlabel metal2 s 296442 0 296498 800 6 la_data_out[102]
port 931 nsew signal output
rlabel metal2 s 298558 0 298614 800 6 la_data_out[103]
port 932 nsew signal output
rlabel metal2 s 300766 0 300822 800 6 la_data_out[104]
port 933 nsew signal output
rlabel metal2 s 302882 0 302938 800 6 la_data_out[105]
port 934 nsew signal output
rlabel metal2 s 304998 0 305054 800 6 la_data_out[106]
port 935 nsew signal output
rlabel metal2 s 307206 0 307262 800 6 la_data_out[107]
port 936 nsew signal output
rlabel metal2 s 309322 0 309378 800 6 la_data_out[108]
port 937 nsew signal output
rlabel metal2 s 311530 0 311586 800 6 la_data_out[109]
port 938 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[10]
port 939 nsew signal output
rlabel metal2 s 313646 0 313702 800 6 la_data_out[110]
port 940 nsew signal output
rlabel metal2 s 315762 0 315818 800 6 la_data_out[111]
port 941 nsew signal output
rlabel metal2 s 317970 0 318026 800 6 la_data_out[112]
port 942 nsew signal output
rlabel metal2 s 320086 0 320142 800 6 la_data_out[113]
port 943 nsew signal output
rlabel metal2 s 322294 0 322350 800 6 la_data_out[114]
port 944 nsew signal output
rlabel metal2 s 324410 0 324466 800 6 la_data_out[115]
port 945 nsew signal output
rlabel metal2 s 326526 0 326582 800 6 la_data_out[116]
port 946 nsew signal output
rlabel metal2 s 328734 0 328790 800 6 la_data_out[117]
port 947 nsew signal output
rlabel metal2 s 330850 0 330906 800 6 la_data_out[118]
port 948 nsew signal output
rlabel metal2 s 332966 0 333022 800 6 la_data_out[119]
port 949 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[11]
port 950 nsew signal output
rlabel metal2 s 335174 0 335230 800 6 la_data_out[120]
port 951 nsew signal output
rlabel metal2 s 337290 0 337346 800 6 la_data_out[121]
port 952 nsew signal output
rlabel metal2 s 339498 0 339554 800 6 la_data_out[122]
port 953 nsew signal output
rlabel metal2 s 341614 0 341670 800 6 la_data_out[123]
port 954 nsew signal output
rlabel metal2 s 343730 0 343786 800 6 la_data_out[124]
port 955 nsew signal output
rlabel metal2 s 345938 0 345994 800 6 la_data_out[125]
port 956 nsew signal output
rlabel metal2 s 348054 0 348110 800 6 la_data_out[126]
port 957 nsew signal output
rlabel metal2 s 350262 0 350318 800 6 la_data_out[127]
port 958 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[12]
port 959 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 la_data_out[13]
port 960 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[14]
port 961 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[15]
port 962 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[16]
port 963 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 la_data_out[17]
port 964 nsew signal output
rlabel metal2 s 115754 0 115810 800 6 la_data_out[18]
port 965 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[19]
port 966 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[1]
port 967 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 la_data_out[20]
port 968 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 la_data_out[21]
port 969 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 la_data_out[22]
port 970 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[23]
port 971 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[24]
port 972 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[25]
port 973 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[26]
port 974 nsew signal output
rlabel metal2 s 135074 0 135130 800 6 la_data_out[27]
port 975 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[28]
port 976 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[29]
port 977 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[2]
port 978 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[30]
port 979 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 la_data_out[31]
port 980 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[32]
port 981 nsew signal output
rlabel metal2 s 147954 0 148010 800 6 la_data_out[33]
port 982 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[34]
port 983 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[35]
port 984 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[36]
port 985 nsew signal output
rlabel metal2 s 156602 0 156658 800 6 la_data_out[37]
port 986 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 la_data_out[38]
port 987 nsew signal output
rlabel metal2 s 160926 0 160982 800 6 la_data_out[39]
port 988 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[3]
port 989 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 la_data_out[40]
port 990 nsew signal output
rlabel metal2 s 165158 0 165214 800 6 la_data_out[41]
port 991 nsew signal output
rlabel metal2 s 167366 0 167422 800 6 la_data_out[42]
port 992 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[43]
port 993 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 la_data_out[44]
port 994 nsew signal output
rlabel metal2 s 173806 0 173862 800 6 la_data_out[45]
port 995 nsew signal output
rlabel metal2 s 175922 0 175978 800 6 la_data_out[46]
port 996 nsew signal output
rlabel metal2 s 178130 0 178186 800 6 la_data_out[47]
port 997 nsew signal output
rlabel metal2 s 180246 0 180302 800 6 la_data_out[48]
port 998 nsew signal output
rlabel metal2 s 182362 0 182418 800 6 la_data_out[49]
port 999 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[4]
port 1000 nsew signal output
rlabel metal2 s 184570 0 184626 800 6 la_data_out[50]
port 1001 nsew signal output
rlabel metal2 s 186686 0 186742 800 6 la_data_out[51]
port 1002 nsew signal output
rlabel metal2 s 188894 0 188950 800 6 la_data_out[52]
port 1003 nsew signal output
rlabel metal2 s 191010 0 191066 800 6 la_data_out[53]
port 1004 nsew signal output
rlabel metal2 s 193126 0 193182 800 6 la_data_out[54]
port 1005 nsew signal output
rlabel metal2 s 195334 0 195390 800 6 la_data_out[55]
port 1006 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 la_data_out[56]
port 1007 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 la_data_out[57]
port 1008 nsew signal output
rlabel metal2 s 201774 0 201830 800 6 la_data_out[58]
port 1009 nsew signal output
rlabel metal2 s 203890 0 203946 800 6 la_data_out[59]
port 1010 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[5]
port 1011 nsew signal output
rlabel metal2 s 206098 0 206154 800 6 la_data_out[60]
port 1012 nsew signal output
rlabel metal2 s 208214 0 208270 800 6 la_data_out[61]
port 1013 nsew signal output
rlabel metal2 s 210330 0 210386 800 6 la_data_out[62]
port 1014 nsew signal output
rlabel metal2 s 212538 0 212594 800 6 la_data_out[63]
port 1015 nsew signal output
rlabel metal2 s 214654 0 214710 800 6 la_data_out[64]
port 1016 nsew signal output
rlabel metal2 s 216862 0 216918 800 6 la_data_out[65]
port 1017 nsew signal output
rlabel metal2 s 218978 0 219034 800 6 la_data_out[66]
port 1018 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 la_data_out[67]
port 1019 nsew signal output
rlabel metal2 s 223302 0 223358 800 6 la_data_out[68]
port 1020 nsew signal output
rlabel metal2 s 225418 0 225474 800 6 la_data_out[69]
port 1021 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[6]
port 1022 nsew signal output
rlabel metal2 s 227626 0 227682 800 6 la_data_out[70]
port 1023 nsew signal output
rlabel metal2 s 229742 0 229798 800 6 la_data_out[71]
port 1024 nsew signal output
rlabel metal2 s 231858 0 231914 800 6 la_data_out[72]
port 1025 nsew signal output
rlabel metal2 s 234066 0 234122 800 6 la_data_out[73]
port 1026 nsew signal output
rlabel metal2 s 236182 0 236238 800 6 la_data_out[74]
port 1027 nsew signal output
rlabel metal2 s 238298 0 238354 800 6 la_data_out[75]
port 1028 nsew signal output
rlabel metal2 s 240506 0 240562 800 6 la_data_out[76]
port 1029 nsew signal output
rlabel metal2 s 242622 0 242678 800 6 la_data_out[77]
port 1030 nsew signal output
rlabel metal2 s 244830 0 244886 800 6 la_data_out[78]
port 1031 nsew signal output
rlabel metal2 s 246946 0 247002 800 6 la_data_out[79]
port 1032 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[7]
port 1033 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 la_data_out[80]
port 1034 nsew signal output
rlabel metal2 s 251270 0 251326 800 6 la_data_out[81]
port 1035 nsew signal output
rlabel metal2 s 253386 0 253442 800 6 la_data_out[82]
port 1036 nsew signal output
rlabel metal2 s 255594 0 255650 800 6 la_data_out[83]
port 1037 nsew signal output
rlabel metal2 s 257710 0 257766 800 6 la_data_out[84]
port 1038 nsew signal output
rlabel metal2 s 259826 0 259882 800 6 la_data_out[85]
port 1039 nsew signal output
rlabel metal2 s 262034 0 262090 800 6 la_data_out[86]
port 1040 nsew signal output
rlabel metal2 s 264150 0 264206 800 6 la_data_out[87]
port 1041 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[88]
port 1042 nsew signal output
rlabel metal2 s 268474 0 268530 800 6 la_data_out[89]
port 1043 nsew signal output
rlabel metal2 s 94226 0 94282 800 6 la_data_out[8]
port 1044 nsew signal output
rlabel metal2 s 270590 0 270646 800 6 la_data_out[90]
port 1045 nsew signal output
rlabel metal2 s 272798 0 272854 800 6 la_data_out[91]
port 1046 nsew signal output
rlabel metal2 s 274914 0 274970 800 6 la_data_out[92]
port 1047 nsew signal output
rlabel metal2 s 277030 0 277086 800 6 la_data_out[93]
port 1048 nsew signal output
rlabel metal2 s 279238 0 279294 800 6 la_data_out[94]
port 1049 nsew signal output
rlabel metal2 s 281354 0 281410 800 6 la_data_out[95]
port 1050 nsew signal output
rlabel metal2 s 283562 0 283618 800 6 la_data_out[96]
port 1051 nsew signal output
rlabel metal2 s 285678 0 285734 800 6 la_data_out[97]
port 1052 nsew signal output
rlabel metal2 s 287794 0 287850 800 6 la_data_out[98]
port 1053 nsew signal output
rlabel metal2 s 290002 0 290058 800 6 la_data_out[99]
port 1054 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[9]
port 1055 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_oenb[0]
port 1056 nsew signal input
rlabel metal2 s 292854 0 292910 800 6 la_oenb[100]
port 1057 nsew signal input
rlabel metal2 s 294970 0 295026 800 6 la_oenb[101]
port 1058 nsew signal input
rlabel metal2 s 297178 0 297234 800 6 la_oenb[102]
port 1059 nsew signal input
rlabel metal2 s 299294 0 299350 800 6 la_oenb[103]
port 1060 nsew signal input
rlabel metal2 s 301410 0 301466 800 6 la_oenb[104]
port 1061 nsew signal input
rlabel metal2 s 303618 0 303674 800 6 la_oenb[105]
port 1062 nsew signal input
rlabel metal2 s 305734 0 305790 800 6 la_oenb[106]
port 1063 nsew signal input
rlabel metal2 s 307942 0 307998 800 6 la_oenb[107]
port 1064 nsew signal input
rlabel metal2 s 310058 0 310114 800 6 la_oenb[108]
port 1065 nsew signal input
rlabel metal2 s 312174 0 312230 800 6 la_oenb[109]
port 1066 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[10]
port 1067 nsew signal input
rlabel metal2 s 314382 0 314438 800 6 la_oenb[110]
port 1068 nsew signal input
rlabel metal2 s 316498 0 316554 800 6 la_oenb[111]
port 1069 nsew signal input
rlabel metal2 s 318706 0 318762 800 6 la_oenb[112]
port 1070 nsew signal input
rlabel metal2 s 320822 0 320878 800 6 la_oenb[113]
port 1071 nsew signal input
rlabel metal2 s 322938 0 322994 800 6 la_oenb[114]
port 1072 nsew signal input
rlabel metal2 s 325146 0 325202 800 6 la_oenb[115]
port 1073 nsew signal input
rlabel metal2 s 327262 0 327318 800 6 la_oenb[116]
port 1074 nsew signal input
rlabel metal2 s 329378 0 329434 800 6 la_oenb[117]
port 1075 nsew signal input
rlabel metal2 s 331586 0 331642 800 6 la_oenb[118]
port 1076 nsew signal input
rlabel metal2 s 333702 0 333758 800 6 la_oenb[119]
port 1077 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_oenb[11]
port 1078 nsew signal input
rlabel metal2 s 335910 0 335966 800 6 la_oenb[120]
port 1079 nsew signal input
rlabel metal2 s 338026 0 338082 800 6 la_oenb[121]
port 1080 nsew signal input
rlabel metal2 s 340142 0 340198 800 6 la_oenb[122]
port 1081 nsew signal input
rlabel metal2 s 342350 0 342406 800 6 la_oenb[123]
port 1082 nsew signal input
rlabel metal2 s 344466 0 344522 800 6 la_oenb[124]
port 1083 nsew signal input
rlabel metal2 s 346674 0 346730 800 6 la_oenb[125]
port 1084 nsew signal input
rlabel metal2 s 348790 0 348846 800 6 la_oenb[126]
port 1085 nsew signal input
rlabel metal2 s 350906 0 350962 800 6 la_oenb[127]
port 1086 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_oenb[12]
port 1087 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_oenb[13]
port 1088 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_oenb[14]
port 1089 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_oenb[15]
port 1090 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_oenb[16]
port 1091 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_oenb[17]
port 1092 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[18]
port 1093 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_oenb[19]
port 1094 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[1]
port 1095 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[20]
port 1096 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_oenb[21]
port 1097 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_oenb[22]
port 1098 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_oenb[23]
port 1099 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_oenb[24]
port 1100 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[25]
port 1101 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[26]
port 1102 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_oenb[27]
port 1103 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[28]
port 1104 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_oenb[29]
port 1105 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[2]
port 1106 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[30]
port 1107 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_oenb[31]
port 1108 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_oenb[32]
port 1109 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_oenb[33]
port 1110 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_oenb[34]
port 1111 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[35]
port 1112 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oenb[36]
port 1113 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oenb[37]
port 1114 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_oenb[38]
port 1115 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_oenb[39]
port 1116 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[3]
port 1117 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oenb[40]
port 1118 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oenb[41]
port 1119 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_oenb[42]
port 1120 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_oenb[43]
port 1121 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 la_oenb[44]
port 1122 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_oenb[45]
port 1123 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 la_oenb[46]
port 1124 nsew signal input
rlabel metal2 s 178774 0 178830 800 6 la_oenb[47]
port 1125 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_oenb[48]
port 1126 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_oenb[49]
port 1127 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[4]
port 1128 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 la_oenb[50]
port 1129 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_oenb[51]
port 1130 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_oenb[52]
port 1131 nsew signal input
rlabel metal2 s 191746 0 191802 800 6 la_oenb[53]
port 1132 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_oenb[54]
port 1133 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_oenb[55]
port 1134 nsew signal input
rlabel metal2 s 198186 0 198242 800 6 la_oenb[56]
port 1135 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_oenb[57]
port 1136 nsew signal input
rlabel metal2 s 202510 0 202566 800 6 la_oenb[58]
port 1137 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_oenb[59]
port 1138 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[5]
port 1139 nsew signal input
rlabel metal2 s 206742 0 206798 800 6 la_oenb[60]
port 1140 nsew signal input
rlabel metal2 s 208950 0 209006 800 6 la_oenb[61]
port 1141 nsew signal input
rlabel metal2 s 211066 0 211122 800 6 la_oenb[62]
port 1142 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_oenb[63]
port 1143 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_oenb[64]
port 1144 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_oenb[65]
port 1145 nsew signal input
rlabel metal2 s 219714 0 219770 800 6 la_oenb[66]
port 1146 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 la_oenb[67]
port 1147 nsew signal input
rlabel metal2 s 224038 0 224094 800 6 la_oenb[68]
port 1148 nsew signal input
rlabel metal2 s 226154 0 226210 800 6 la_oenb[69]
port 1149 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[6]
port 1150 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_oenb[70]
port 1151 nsew signal input
rlabel metal2 s 230478 0 230534 800 6 la_oenb[71]
port 1152 nsew signal input
rlabel metal2 s 232594 0 232650 800 6 la_oenb[72]
port 1153 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_oenb[73]
port 1154 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 la_oenb[74]
port 1155 nsew signal input
rlabel metal2 s 239034 0 239090 800 6 la_oenb[75]
port 1156 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 la_oenb[76]
port 1157 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_oenb[77]
port 1158 nsew signal input
rlabel metal2 s 245474 0 245530 800 6 la_oenb[78]
port 1159 nsew signal input
rlabel metal2 s 247682 0 247738 800 6 la_oenb[79]
port 1160 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[7]
port 1161 nsew signal input
rlabel metal2 s 249798 0 249854 800 6 la_oenb[80]
port 1162 nsew signal input
rlabel metal2 s 252006 0 252062 800 6 la_oenb[81]
port 1163 nsew signal input
rlabel metal2 s 254122 0 254178 800 6 la_oenb[82]
port 1164 nsew signal input
rlabel metal2 s 256238 0 256294 800 6 la_oenb[83]
port 1165 nsew signal input
rlabel metal2 s 258446 0 258502 800 6 la_oenb[84]
port 1166 nsew signal input
rlabel metal2 s 260562 0 260618 800 6 la_oenb[85]
port 1167 nsew signal input
rlabel metal2 s 262770 0 262826 800 6 la_oenb[86]
port 1168 nsew signal input
rlabel metal2 s 264886 0 264942 800 6 la_oenb[87]
port 1169 nsew signal input
rlabel metal2 s 267002 0 267058 800 6 la_oenb[88]
port 1170 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 la_oenb[89]
port 1171 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[8]
port 1172 nsew signal input
rlabel metal2 s 271326 0 271382 800 6 la_oenb[90]
port 1173 nsew signal input
rlabel metal2 s 273442 0 273498 800 6 la_oenb[91]
port 1174 nsew signal input
rlabel metal2 s 275650 0 275706 800 6 la_oenb[92]
port 1175 nsew signal input
rlabel metal2 s 277766 0 277822 800 6 la_oenb[93]
port 1176 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 la_oenb[94]
port 1177 nsew signal input
rlabel metal2 s 282090 0 282146 800 6 la_oenb[95]
port 1178 nsew signal input
rlabel metal2 s 284206 0 284262 800 6 la_oenb[96]
port 1179 nsew signal input
rlabel metal2 s 286414 0 286470 800 6 la_oenb[97]
port 1180 nsew signal input
rlabel metal2 s 288530 0 288586 800 6 la_oenb[98]
port 1181 nsew signal input
rlabel metal2 s 290738 0 290794 800 6 la_oenb[99]
port 1182 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[9]
port 1183 nsew signal input
rlabel metal3 s 0 327632 800 327752 6 tag_array_ext_ram_addr1[0]
port 1184 nsew signal output
rlabel metal3 s 0 328448 800 328568 6 tag_array_ext_ram_addr1[1]
port 1185 nsew signal output
rlabel metal3 s 0 329128 800 329248 6 tag_array_ext_ram_addr1[2]
port 1186 nsew signal output
rlabel metal3 s 0 329808 800 329928 6 tag_array_ext_ram_addr1[3]
port 1187 nsew signal output
rlabel metal3 s 0 330488 800 330608 6 tag_array_ext_ram_addr1[4]
port 1188 nsew signal output
rlabel metal3 s 0 331168 800 331288 6 tag_array_ext_ram_addr1[5]
port 1189 nsew signal output
rlabel metal3 s 0 331848 800 331968 6 tag_array_ext_ram_addr1[6]
port 1190 nsew signal output
rlabel metal3 s 0 332664 800 332784 6 tag_array_ext_ram_addr1[7]
port 1191 nsew signal output
rlabel metal3 s 0 272008 800 272128 6 tag_array_ext_ram_addr[0]
port 1192 nsew signal output
rlabel metal3 s 0 272688 800 272808 6 tag_array_ext_ram_addr[1]
port 1193 nsew signal output
rlabel metal3 s 0 273504 800 273624 6 tag_array_ext_ram_addr[2]
port 1194 nsew signal output
rlabel metal3 s 0 274184 800 274304 6 tag_array_ext_ram_addr[3]
port 1195 nsew signal output
rlabel metal3 s 0 274864 800 274984 6 tag_array_ext_ram_addr[4]
port 1196 nsew signal output
rlabel metal3 s 0 275544 800 275664 6 tag_array_ext_ram_addr[5]
port 1197 nsew signal output
rlabel metal3 s 0 276224 800 276344 6 tag_array_ext_ram_addr[6]
port 1198 nsew signal output
rlabel metal3 s 0 277040 800 277160 6 tag_array_ext_ram_addr[7]
port 1199 nsew signal output
rlabel metal3 s 0 277720 800 277840 6 tag_array_ext_ram_clk
port 1200 nsew signal output
rlabel metal3 s 0 324912 800 325032 6 tag_array_ext_ram_csb
port 1201 nsew signal output
rlabel metal3 s 0 326272 800 326392 6 tag_array_ext_ram_csb1[0]
port 1202 nsew signal output
rlabel metal3 s 0 326952 800 327072 6 tag_array_ext_ram_csb1[1]
port 1203 nsew signal output
rlabel metal3 s 0 249568 800 249688 6 tag_array_ext_ram_rdata0[0]
port 1204 nsew signal input
rlabel metal3 s 0 256504 800 256624 6 tag_array_ext_ram_rdata0[10]
port 1205 nsew signal input
rlabel metal3 s 0 257320 800 257440 6 tag_array_ext_ram_rdata0[11]
port 1206 nsew signal input
rlabel metal3 s 0 258000 800 258120 6 tag_array_ext_ram_rdata0[12]
port 1207 nsew signal input
rlabel metal3 s 0 258680 800 258800 6 tag_array_ext_ram_rdata0[13]
port 1208 nsew signal input
rlabel metal3 s 0 259360 800 259480 6 tag_array_ext_ram_rdata0[14]
port 1209 nsew signal input
rlabel metal3 s 0 260040 800 260160 6 tag_array_ext_ram_rdata0[15]
port 1210 nsew signal input
rlabel metal3 s 0 260720 800 260840 6 tag_array_ext_ram_rdata0[16]
port 1211 nsew signal input
rlabel metal3 s 0 261536 800 261656 6 tag_array_ext_ram_rdata0[17]
port 1212 nsew signal input
rlabel metal3 s 0 262216 800 262336 6 tag_array_ext_ram_rdata0[18]
port 1213 nsew signal input
rlabel metal3 s 0 262896 800 263016 6 tag_array_ext_ram_rdata0[19]
port 1214 nsew signal input
rlabel metal3 s 0 250248 800 250368 6 tag_array_ext_ram_rdata0[1]
port 1215 nsew signal input
rlabel metal3 s 0 263576 800 263696 6 tag_array_ext_ram_rdata0[20]
port 1216 nsew signal input
rlabel metal3 s 0 264256 800 264376 6 tag_array_ext_ram_rdata0[21]
port 1217 nsew signal input
rlabel metal3 s 0 265072 800 265192 6 tag_array_ext_ram_rdata0[22]
port 1218 nsew signal input
rlabel metal3 s 0 265752 800 265872 6 tag_array_ext_ram_rdata0[23]
port 1219 nsew signal input
rlabel metal3 s 0 266432 800 266552 6 tag_array_ext_ram_rdata0[24]
port 1220 nsew signal input
rlabel metal3 s 0 267112 800 267232 6 tag_array_ext_ram_rdata0[25]
port 1221 nsew signal input
rlabel metal3 s 0 267792 800 267912 6 tag_array_ext_ram_rdata0[26]
port 1222 nsew signal input
rlabel metal3 s 0 268472 800 268592 6 tag_array_ext_ram_rdata0[27]
port 1223 nsew signal input
rlabel metal3 s 0 269288 800 269408 6 tag_array_ext_ram_rdata0[28]
port 1224 nsew signal input
rlabel metal3 s 0 269968 800 270088 6 tag_array_ext_ram_rdata0[29]
port 1225 nsew signal input
rlabel metal3 s 0 250928 800 251048 6 tag_array_ext_ram_rdata0[2]
port 1226 nsew signal input
rlabel metal3 s 0 270648 800 270768 6 tag_array_ext_ram_rdata0[30]
port 1227 nsew signal input
rlabel metal3 s 0 271328 800 271448 6 tag_array_ext_ram_rdata0[31]
port 1228 nsew signal input
rlabel metal3 s 0 251608 800 251728 6 tag_array_ext_ram_rdata0[3]
port 1229 nsew signal input
rlabel metal3 s 0 252288 800 252408 6 tag_array_ext_ram_rdata0[4]
port 1230 nsew signal input
rlabel metal3 s 0 252968 800 253088 6 tag_array_ext_ram_rdata0[5]
port 1231 nsew signal input
rlabel metal3 s 0 253784 800 253904 6 tag_array_ext_ram_rdata0[6]
port 1232 nsew signal input
rlabel metal3 s 0 254464 800 254584 6 tag_array_ext_ram_rdata0[7]
port 1233 nsew signal input
rlabel metal3 s 0 255144 800 255264 6 tag_array_ext_ram_rdata0[8]
port 1234 nsew signal input
rlabel metal3 s 0 255824 800 255944 6 tag_array_ext_ram_rdata0[9]
port 1235 nsew signal input
rlabel metal3 s 0 333344 800 333464 6 tag_array_ext_ram_rdata1[0]
port 1236 nsew signal input
rlabel metal3 s 0 340416 800 340536 6 tag_array_ext_ram_rdata1[10]
port 1237 nsew signal input
rlabel metal3 s 0 341096 800 341216 6 tag_array_ext_ram_rdata1[11]
port 1238 nsew signal input
rlabel metal3 s 0 341776 800 341896 6 tag_array_ext_ram_rdata1[12]
port 1239 nsew signal input
rlabel metal3 s 0 342456 800 342576 6 tag_array_ext_ram_rdata1[13]
port 1240 nsew signal input
rlabel metal3 s 0 343136 800 343256 6 tag_array_ext_ram_rdata1[14]
port 1241 nsew signal input
rlabel metal3 s 0 343816 800 343936 6 tag_array_ext_ram_rdata1[15]
port 1242 nsew signal input
rlabel metal3 s 0 344632 800 344752 6 tag_array_ext_ram_rdata1[16]
port 1243 nsew signal input
rlabel metal3 s 0 345312 800 345432 6 tag_array_ext_ram_rdata1[17]
port 1244 nsew signal input
rlabel metal3 s 0 345992 800 346112 6 tag_array_ext_ram_rdata1[18]
port 1245 nsew signal input
rlabel metal3 s 0 346672 800 346792 6 tag_array_ext_ram_rdata1[19]
port 1246 nsew signal input
rlabel metal3 s 0 334024 800 334144 6 tag_array_ext_ram_rdata1[1]
port 1247 nsew signal input
rlabel metal3 s 0 347352 800 347472 6 tag_array_ext_ram_rdata1[20]
port 1248 nsew signal input
rlabel metal3 s 0 348168 800 348288 6 tag_array_ext_ram_rdata1[21]
port 1249 nsew signal input
rlabel metal3 s 0 348848 800 348968 6 tag_array_ext_ram_rdata1[22]
port 1250 nsew signal input
rlabel metal3 s 0 349528 800 349648 6 tag_array_ext_ram_rdata1[23]
port 1251 nsew signal input
rlabel metal3 s 0 350208 800 350328 6 tag_array_ext_ram_rdata1[24]
port 1252 nsew signal input
rlabel metal3 s 0 350888 800 351008 6 tag_array_ext_ram_rdata1[25]
port 1253 nsew signal input
rlabel metal3 s 0 351568 800 351688 6 tag_array_ext_ram_rdata1[26]
port 1254 nsew signal input
rlabel metal3 s 0 352384 800 352504 6 tag_array_ext_ram_rdata1[27]
port 1255 nsew signal input
rlabel metal3 s 0 353064 800 353184 6 tag_array_ext_ram_rdata1[28]
port 1256 nsew signal input
rlabel metal3 s 0 353744 800 353864 6 tag_array_ext_ram_rdata1[29]
port 1257 nsew signal input
rlabel metal3 s 0 334704 800 334824 6 tag_array_ext_ram_rdata1[2]
port 1258 nsew signal input
rlabel metal3 s 0 354424 800 354544 6 tag_array_ext_ram_rdata1[30]
port 1259 nsew signal input
rlabel metal3 s 0 355104 800 355224 6 tag_array_ext_ram_rdata1[31]
port 1260 nsew signal input
rlabel metal3 s 0 335384 800 335504 6 tag_array_ext_ram_rdata1[3]
port 1261 nsew signal input
rlabel metal3 s 0 336200 800 336320 6 tag_array_ext_ram_rdata1[4]
port 1262 nsew signal input
rlabel metal3 s 0 336880 800 337000 6 tag_array_ext_ram_rdata1[5]
port 1263 nsew signal input
rlabel metal3 s 0 337560 800 337680 6 tag_array_ext_ram_rdata1[6]
port 1264 nsew signal input
rlabel metal3 s 0 338240 800 338360 6 tag_array_ext_ram_rdata1[7]
port 1265 nsew signal input
rlabel metal3 s 0 338920 800 339040 6 tag_array_ext_ram_rdata1[8]
port 1266 nsew signal input
rlabel metal3 s 0 339600 800 339720 6 tag_array_ext_ram_rdata1[9]
port 1267 nsew signal input
rlabel metal3 s 0 278400 800 278520 6 tag_array_ext_ram_wdata[0]
port 1268 nsew signal output
rlabel metal3 s 0 285472 800 285592 6 tag_array_ext_ram_wdata[10]
port 1269 nsew signal output
rlabel metal3 s 0 286152 800 286272 6 tag_array_ext_ram_wdata[11]
port 1270 nsew signal output
rlabel metal3 s 0 286832 800 286952 6 tag_array_ext_ram_wdata[12]
port 1271 nsew signal output
rlabel metal3 s 0 287512 800 287632 6 tag_array_ext_ram_wdata[13]
port 1272 nsew signal output
rlabel metal3 s 0 288192 800 288312 6 tag_array_ext_ram_wdata[14]
port 1273 nsew signal output
rlabel metal3 s 0 289008 800 289128 6 tag_array_ext_ram_wdata[15]
port 1274 nsew signal output
rlabel metal3 s 0 289688 800 289808 6 tag_array_ext_ram_wdata[16]
port 1275 nsew signal output
rlabel metal3 s 0 290368 800 290488 6 tag_array_ext_ram_wdata[17]
port 1276 nsew signal output
rlabel metal3 s 0 291048 800 291168 6 tag_array_ext_ram_wdata[18]
port 1277 nsew signal output
rlabel metal3 s 0 291728 800 291848 6 tag_array_ext_ram_wdata[19]
port 1278 nsew signal output
rlabel metal3 s 0 279080 800 279200 6 tag_array_ext_ram_wdata[1]
port 1279 nsew signal output
rlabel metal3 s 0 292408 800 292528 6 tag_array_ext_ram_wdata[20]
port 1280 nsew signal output
rlabel metal3 s 0 293224 800 293344 6 tag_array_ext_ram_wdata[21]
port 1281 nsew signal output
rlabel metal3 s 0 293904 800 294024 6 tag_array_ext_ram_wdata[22]
port 1282 nsew signal output
rlabel metal3 s 0 294584 800 294704 6 tag_array_ext_ram_wdata[23]
port 1283 nsew signal output
rlabel metal3 s 0 295264 800 295384 6 tag_array_ext_ram_wdata[24]
port 1284 nsew signal output
rlabel metal3 s 0 295944 800 296064 6 tag_array_ext_ram_wdata[25]
port 1285 nsew signal output
rlabel metal3 s 0 296760 800 296880 6 tag_array_ext_ram_wdata[26]
port 1286 nsew signal output
rlabel metal3 s 0 297440 800 297560 6 tag_array_ext_ram_wdata[27]
port 1287 nsew signal output
rlabel metal3 s 0 298120 800 298240 6 tag_array_ext_ram_wdata[28]
port 1288 nsew signal output
rlabel metal3 s 0 298800 800 298920 6 tag_array_ext_ram_wdata[29]
port 1289 nsew signal output
rlabel metal3 s 0 279760 800 279880 6 tag_array_ext_ram_wdata[2]
port 1290 nsew signal output
rlabel metal3 s 0 299480 800 299600 6 tag_array_ext_ram_wdata[30]
port 1291 nsew signal output
rlabel metal3 s 0 300160 800 300280 6 tag_array_ext_ram_wdata[31]
port 1292 nsew signal output
rlabel metal3 s 0 300976 800 301096 6 tag_array_ext_ram_wdata[32]
port 1293 nsew signal output
rlabel metal3 s 0 301656 800 301776 6 tag_array_ext_ram_wdata[33]
port 1294 nsew signal output
rlabel metal3 s 0 302336 800 302456 6 tag_array_ext_ram_wdata[34]
port 1295 nsew signal output
rlabel metal3 s 0 303016 800 303136 6 tag_array_ext_ram_wdata[35]
port 1296 nsew signal output
rlabel metal3 s 0 303696 800 303816 6 tag_array_ext_ram_wdata[36]
port 1297 nsew signal output
rlabel metal3 s 0 304376 800 304496 6 tag_array_ext_ram_wdata[37]
port 1298 nsew signal output
rlabel metal3 s 0 305192 800 305312 6 tag_array_ext_ram_wdata[38]
port 1299 nsew signal output
rlabel metal3 s 0 305872 800 305992 6 tag_array_ext_ram_wdata[39]
port 1300 nsew signal output
rlabel metal3 s 0 280440 800 280560 6 tag_array_ext_ram_wdata[3]
port 1301 nsew signal output
rlabel metal3 s 0 306552 800 306672 6 tag_array_ext_ram_wdata[40]
port 1302 nsew signal output
rlabel metal3 s 0 307232 800 307352 6 tag_array_ext_ram_wdata[41]
port 1303 nsew signal output
rlabel metal3 s 0 307912 800 308032 6 tag_array_ext_ram_wdata[42]
port 1304 nsew signal output
rlabel metal3 s 0 308728 800 308848 6 tag_array_ext_ram_wdata[43]
port 1305 nsew signal output
rlabel metal3 s 0 309408 800 309528 6 tag_array_ext_ram_wdata[44]
port 1306 nsew signal output
rlabel metal3 s 0 310088 800 310208 6 tag_array_ext_ram_wdata[45]
port 1307 nsew signal output
rlabel metal3 s 0 310768 800 310888 6 tag_array_ext_ram_wdata[46]
port 1308 nsew signal output
rlabel metal3 s 0 311448 800 311568 6 tag_array_ext_ram_wdata[47]
port 1309 nsew signal output
rlabel metal3 s 0 312128 800 312248 6 tag_array_ext_ram_wdata[48]
port 1310 nsew signal output
rlabel metal3 s 0 312944 800 313064 6 tag_array_ext_ram_wdata[49]
port 1311 nsew signal output
rlabel metal3 s 0 281256 800 281376 6 tag_array_ext_ram_wdata[4]
port 1312 nsew signal output
rlabel metal3 s 0 313624 800 313744 6 tag_array_ext_ram_wdata[50]
port 1313 nsew signal output
rlabel metal3 s 0 314304 800 314424 6 tag_array_ext_ram_wdata[51]
port 1314 nsew signal output
rlabel metal3 s 0 314984 800 315104 6 tag_array_ext_ram_wdata[52]
port 1315 nsew signal output
rlabel metal3 s 0 315664 800 315784 6 tag_array_ext_ram_wdata[53]
port 1316 nsew signal output
rlabel metal3 s 0 316480 800 316600 6 tag_array_ext_ram_wdata[54]
port 1317 nsew signal output
rlabel metal3 s 0 317160 800 317280 6 tag_array_ext_ram_wdata[55]
port 1318 nsew signal output
rlabel metal3 s 0 317840 800 317960 6 tag_array_ext_ram_wdata[56]
port 1319 nsew signal output
rlabel metal3 s 0 318520 800 318640 6 tag_array_ext_ram_wdata[57]
port 1320 nsew signal output
rlabel metal3 s 0 319200 800 319320 6 tag_array_ext_ram_wdata[58]
port 1321 nsew signal output
rlabel metal3 s 0 319880 800 320000 6 tag_array_ext_ram_wdata[59]
port 1322 nsew signal output
rlabel metal3 s 0 281936 800 282056 6 tag_array_ext_ram_wdata[5]
port 1323 nsew signal output
rlabel metal3 s 0 320696 800 320816 6 tag_array_ext_ram_wdata[60]
port 1324 nsew signal output
rlabel metal3 s 0 321376 800 321496 6 tag_array_ext_ram_wdata[61]
port 1325 nsew signal output
rlabel metal3 s 0 322056 800 322176 6 tag_array_ext_ram_wdata[62]
port 1326 nsew signal output
rlabel metal3 s 0 322736 800 322856 6 tag_array_ext_ram_wdata[63]
port 1327 nsew signal output
rlabel metal3 s 0 282616 800 282736 6 tag_array_ext_ram_wdata[6]
port 1328 nsew signal output
rlabel metal3 s 0 283296 800 283416 6 tag_array_ext_ram_wdata[7]
port 1329 nsew signal output
rlabel metal3 s 0 283976 800 284096 6 tag_array_ext_ram_wdata[8]
port 1330 nsew signal output
rlabel metal3 s 0 284792 800 284912 6 tag_array_ext_ram_wdata[9]
port 1331 nsew signal output
rlabel metal3 s 0 325592 800 325712 6 tag_array_ext_ram_web
port 1332 nsew signal output
rlabel metal3 s 0 323416 800 323536 6 tag_array_ext_ram_wmask[0]
port 1333 nsew signal output
rlabel metal3 s 0 324096 800 324216 6 tag_array_ext_ram_wmask[1]
port 1334 nsew signal output
rlabel metal4 s 4208 2128 4528 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 34928 2128 35248 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 65648 2128 65968 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 96368 2128 96688 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 127088 2128 127408 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 157808 2128 158128 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 188528 2128 188848 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 219248 2128 219568 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 249968 2128 250288 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 280688 2128 281008 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 311408 2128 311728 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 342128 2128 342448 353104 6 vccd1
port 1335 nsew power input
rlabel metal4 s 19568 2128 19888 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 50288 2128 50608 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 81008 2128 81328 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 111728 2128 112048 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 142448 2128 142768 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 173168 2128 173488 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 203888 2128 204208 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 234608 2128 234928 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 265328 2128 265648 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 296048 2128 296368 353104 6 vssd1
port 1336 nsew ground input
rlabel metal4 s 326768 2128 327088 353104 6 vssd1
port 1336 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 1337 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 1338 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_ack_o
port 1339 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[0]
port 1340 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[10]
port 1341 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[11]
port 1342 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[12]
port 1343 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_adr_i[13]
port 1344 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_adr_i[14]
port 1345 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_adr_i[15]
port 1346 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_adr_i[16]
port 1347 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 wbs_adr_i[17]
port 1348 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_adr_i[18]
port 1349 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[19]
port 1350 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[1]
port 1351 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[20]
port 1352 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 wbs_adr_i[21]
port 1353 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 wbs_adr_i[22]
port 1354 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_adr_i[23]
port 1355 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 wbs_adr_i[24]
port 1356 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[25]
port 1357 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 wbs_adr_i[26]
port 1358 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 wbs_adr_i[27]
port 1359 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 wbs_adr_i[28]
port 1360 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 wbs_adr_i[29]
port 1361 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[2]
port 1362 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 wbs_adr_i[30]
port 1363 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_adr_i[31]
port 1364 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_adr_i[3]
port 1365 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[4]
port 1366 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_adr_i[5]
port 1367 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[6]
port 1368 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[7]
port 1369 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[8]
port 1370 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[9]
port 1371 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_cyc_i
port 1372 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_i[0]
port 1373 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_i[10]
port 1374 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[11]
port 1375 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[12]
port 1376 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[13]
port 1377 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[14]
port 1378 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_i[15]
port 1379 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[16]
port 1380 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_i[17]
port 1381 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_i[18]
port 1382 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 wbs_dat_i[19]
port 1383 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[1]
port 1384 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[20]
port 1385 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 wbs_dat_i[21]
port 1386 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_i[22]
port 1387 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_i[23]
port 1388 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_i[24]
port 1389 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_i[25]
port 1390 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_i[26]
port 1391 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wbs_dat_i[27]
port 1392 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_i[28]
port 1393 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 wbs_dat_i[29]
port 1394 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[2]
port 1395 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 wbs_dat_i[30]
port 1396 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 wbs_dat_i[31]
port 1397 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[3]
port 1398 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[4]
port 1399 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[5]
port 1400 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[6]
port 1401 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[7]
port 1402 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[8]
port 1403 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[9]
port 1404 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_o[0]
port 1405 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[10]
port 1406 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_o[11]
port 1407 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_o[12]
port 1408 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[13]
port 1409 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_o[14]
port 1410 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[15]
port 1411 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_o[16]
port 1412 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_o[17]
port 1413 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[18]
port 1414 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_o[19]
port 1415 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[1]
port 1416 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_o[20]
port 1417 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_o[21]
port 1418 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 wbs_dat_o[22]
port 1419 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_o[23]
port 1420 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[24]
port 1421 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 wbs_dat_o[25]
port 1422 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_o[26]
port 1423 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 wbs_dat_o[27]
port 1424 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 wbs_dat_o[28]
port 1425 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 wbs_dat_o[29]
port 1426 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[2]
port 1427 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 wbs_dat_o[30]
port 1428 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_o[31]
port 1429 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[3]
port 1430 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[4]
port 1431 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[5]
port 1432 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_o[6]
port 1433 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[7]
port 1434 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[8]
port 1435 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_o[9]
port 1436 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_sel_i[0]
port 1437 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_sel_i[1]
port 1438 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_sel_i[2]
port 1439 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_sel_i[3]
port 1440 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_stb_i
port 1441 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_we_i
port 1442 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 353520 355664
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 307625600
string GDS_FILE /home/shc/Development/efabless/marmot_asic/openlane/marmot/runs/marmot/results/finishing/Marmot.magic.gds
string GDS_START 2027154
<< end >>

