VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Marmot
  CLASS BLOCK ;
  FOREIGN Marmot ;
  ORIGIN 0.000 0.000 ;
  SIZE 1785.560 BY 1796.280 ;
  PIN data_arrays_0_0_ext_ram_addr00[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END data_arrays_0_0_ext_ram_addr00[0]
  PIN data_arrays_0_0_ext_ram_addr00[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END data_arrays_0_0_ext_ram_addr00[1]
  PIN data_arrays_0_0_ext_ram_addr00[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END data_arrays_0_0_ext_ram_addr00[2]
  PIN data_arrays_0_0_ext_ram_addr00[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END data_arrays_0_0_ext_ram_addr00[3]
  PIN data_arrays_0_0_ext_ram_addr00[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END data_arrays_0_0_ext_ram_addr00[4]
  PIN data_arrays_0_0_ext_ram_addr00[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END data_arrays_0_0_ext_ram_addr00[5]
  PIN data_arrays_0_0_ext_ram_addr00[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END data_arrays_0_0_ext_ram_addr00[6]
  PIN data_arrays_0_0_ext_ram_addr00[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END data_arrays_0_0_ext_ram_addr00[7]
  PIN data_arrays_0_0_ext_ram_addr00[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END data_arrays_0_0_ext_ram_addr00[8]
  PIN data_arrays_0_0_ext_ram_addr01[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1283.200 4.000 1283.800 ;
    END
  END data_arrays_0_0_ext_ram_addr01[0]
  PIN data_arrays_0_0_ext_ram_addr01[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1289.320 4.000 1289.920 ;
    END
  END data_arrays_0_0_ext_ram_addr01[1]
  PIN data_arrays_0_0_ext_ram_addr01[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1294.760 4.000 1295.360 ;
    END
  END data_arrays_0_0_ext_ram_addr01[2]
  PIN data_arrays_0_0_ext_ram_addr01[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.880 4.000 1301.480 ;
    END
  END data_arrays_0_0_ext_ram_addr01[3]
  PIN data_arrays_0_0_ext_ram_addr01[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1307.000 4.000 1307.600 ;
    END
  END data_arrays_0_0_ext_ram_addr01[4]
  PIN data_arrays_0_0_ext_ram_addr01[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1313.120 4.000 1313.720 ;
    END
  END data_arrays_0_0_ext_ram_addr01[5]
  PIN data_arrays_0_0_ext_ram_addr01[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1318.560 4.000 1319.160 ;
    END
  END data_arrays_0_0_ext_ram_addr01[6]
  PIN data_arrays_0_0_ext_ram_addr01[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1324.680 4.000 1325.280 ;
    END
  END data_arrays_0_0_ext_ram_addr01[7]
  PIN data_arrays_0_0_ext_ram_addr01[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1330.800 4.000 1331.400 ;
    END
  END data_arrays_0_0_ext_ram_addr01[8]
  PIN data_arrays_0_0_ext_ram_addr02[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 1792.280 311.330 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr02[0]
  PIN data_arrays_0_0_ext_ram_addr02[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 1792.280 314.550 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr02[1]
  PIN data_arrays_0_0_ext_ram_addr02[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 1792.280 317.770 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr02[2]
  PIN data_arrays_0_0_ext_ram_addr02[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 1792.280 320.990 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr02[3]
  PIN data_arrays_0_0_ext_ram_addr02[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 1792.280 324.210 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr02[4]
  PIN data_arrays_0_0_ext_ram_addr02[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 1792.280 327.890 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr02[5]
  PIN data_arrays_0_0_ext_ram_addr02[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 1792.280 331.110 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr02[6]
  PIN data_arrays_0_0_ext_ram_addr02[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 1792.280 334.330 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr02[7]
  PIN data_arrays_0_0_ext_ram_addr02[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 1792.280 337.550 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr02[8]
  PIN data_arrays_0_0_ext_ram_addr03[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.130 1792.280 1506.410 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr03[0]
  PIN data_arrays_0_0_ext_ram_addr03[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.350 1792.280 1509.630 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr03[1]
  PIN data_arrays_0_0_ext_ram_addr03[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.570 1792.280 1512.850 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr03[2]
  PIN data_arrays_0_0_ext_ram_addr03[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.790 1792.280 1516.070 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr03[3]
  PIN data_arrays_0_0_ext_ram_addr03[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.010 1792.280 1519.290 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr03[4]
  PIN data_arrays_0_0_ext_ram_addr03[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.230 1792.280 1522.510 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr03[5]
  PIN data_arrays_0_0_ext_ram_addr03[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.450 1792.280 1525.730 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr03[6]
  PIN data_arrays_0_0_ext_ram_addr03[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.670 1792.280 1528.950 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr03[7]
  PIN data_arrays_0_0_ext_ram_addr03[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.890 1792.280 1532.170 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr03[8]
  PIN data_arrays_0_0_ext_ram_addr10[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END data_arrays_0_0_ext_ram_addr10[0]
  PIN data_arrays_0_0_ext_ram_addr10[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.160 4.000 856.760 ;
    END
  END data_arrays_0_0_ext_ram_addr10[1]
  PIN data_arrays_0_0_ext_ram_addr10[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END data_arrays_0_0_ext_ram_addr10[2]
  PIN data_arrays_0_0_ext_ram_addr10[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 868.400 4.000 869.000 ;
    END
  END data_arrays_0_0_ext_ram_addr10[3]
  PIN data_arrays_0_0_ext_ram_addr10[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END data_arrays_0_0_ext_ram_addr10[4]
  PIN data_arrays_0_0_ext_ram_addr10[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.960 4.000 880.560 ;
    END
  END data_arrays_0_0_ext_ram_addr10[5]
  PIN data_arrays_0_0_ext_ram_addr10[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END data_arrays_0_0_ext_ram_addr10[6]
  PIN data_arrays_0_0_ext_ram_addr10[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 891.520 4.000 892.120 ;
    END
  END data_arrays_0_0_ext_ram_addr10[7]
  PIN data_arrays_0_0_ext_ram_addr10[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END data_arrays_0_0_ext_ram_addr10[8]
  PIN data_arrays_0_0_ext_ram_addr11[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1745.600 4.000 1746.200 ;
    END
  END data_arrays_0_0_ext_ram_addr11[0]
  PIN data_arrays_0_0_ext_ram_addr11[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.720 4.000 1752.320 ;
    END
  END data_arrays_0_0_ext_ram_addr11[1]
  PIN data_arrays_0_0_ext_ram_addr11[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.160 4.000 1757.760 ;
    END
  END data_arrays_0_0_ext_ram_addr11[2]
  PIN data_arrays_0_0_ext_ram_addr11[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1763.280 4.000 1763.880 ;
    END
  END data_arrays_0_0_ext_ram_addr11[3]
  PIN data_arrays_0_0_ext_ram_addr11[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1769.400 4.000 1770.000 ;
    END
  END data_arrays_0_0_ext_ram_addr11[4]
  PIN data_arrays_0_0_ext_ram_addr11[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1775.520 4.000 1776.120 ;
    END
  END data_arrays_0_0_ext_ram_addr11[5]
  PIN data_arrays_0_0_ext_ram_addr11[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1780.960 4.000 1781.560 ;
    END
  END data_arrays_0_0_ext_ram_addr11[6]
  PIN data_arrays_0_0_ext_ram_addr11[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1787.080 4.000 1787.680 ;
    END
  END data_arrays_0_0_ext_ram_addr11[7]
  PIN data_arrays_0_0_ext_ram_addr11[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1793.200 4.000 1793.800 ;
    END
  END data_arrays_0_0_ext_ram_addr11[8]
  PIN data_arrays_0_0_ext_ram_addr12[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 1792.280 563.410 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr12[0]
  PIN data_arrays_0_0_ext_ram_addr12[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 1792.280 566.630 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr12[1]
  PIN data_arrays_0_0_ext_ram_addr12[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 1792.280 569.850 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr12[2]
  PIN data_arrays_0_0_ext_ram_addr12[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 1792.280 573.070 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr12[3]
  PIN data_arrays_0_0_ext_ram_addr12[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 1792.280 576.290 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr12[4]
  PIN data_arrays_0_0_ext_ram_addr12[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 1792.280 579.510 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr12[5]
  PIN data_arrays_0_0_ext_ram_addr12[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 1792.280 582.730 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr12[6]
  PIN data_arrays_0_0_ext_ram_addr12[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 1792.280 585.950 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr12[7]
  PIN data_arrays_0_0_ext_ram_addr12[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 1792.280 589.170 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr12[8]
  PIN data_arrays_0_0_ext_ram_addr13[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.750 1792.280 1758.030 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr13[0]
  PIN data_arrays_0_0_ext_ram_addr13[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.970 1792.280 1761.250 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr13[1]
  PIN data_arrays_0_0_ext_ram_addr13[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.190 1792.280 1764.470 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr13[2]
  PIN data_arrays_0_0_ext_ram_addr13[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.410 1792.280 1767.690 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr13[3]
  PIN data_arrays_0_0_ext_ram_addr13[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.630 1792.280 1770.910 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr13[4]
  PIN data_arrays_0_0_ext_ram_addr13[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.850 1792.280 1774.130 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr13[5]
  PIN data_arrays_0_0_ext_ram_addr13[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.070 1792.280 1777.350 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr13[6]
  PIN data_arrays_0_0_ext_ram_addr13[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.290 1792.280 1780.570 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr13[7]
  PIN data_arrays_0_0_ext_ram_addr13[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.510 1792.280 1783.790 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_addr13[8]
  PIN data_arrays_0_0_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END data_arrays_0_0_ext_ram_clk
  PIN data_arrays_0_0_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 4.000 845.200 ;
    END
  END data_arrays_0_0_ext_ram_csb1[0]
  PIN data_arrays_0_0_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1739.480 4.000 1740.080 ;
    END
  END data_arrays_0_0_ext_ram_csb1[1]
  PIN data_arrays_0_0_ext_ram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 1792.280 560.190 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_csb1[2]
  PIN data_arrays_0_0_ext_ram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.530 1792.280 1754.810 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_csb1[3]
  PIN data_arrays_0_0_ext_ram_csb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END data_arrays_0_0_ext_ram_csb[0]
  PIN data_arrays_0_0_ext_ram_csb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.920 4.000 1728.520 ;
    END
  END data_arrays_0_0_ext_ram_csb[1]
  PIN data_arrays_0_0_ext_ram_csb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 1792.280 553.750 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_csb[2]
  PIN data_arrays_0_0_ext_ram_csb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.090 1792.280 1748.370 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_csb[3]
  PIN data_arrays_0_0_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[0]
  PIN data_arrays_0_0_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[10]
  PIN data_arrays_0_0_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[11]
  PIN data_arrays_0_0_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[12]
  PIN data_arrays_0_0_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[13]
  PIN data_arrays_0_0_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[14]
  PIN data_arrays_0_0_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[15]
  PIN data_arrays_0_0_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[16]
  PIN data_arrays_0_0_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[17]
  PIN data_arrays_0_0_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[18]
  PIN data_arrays_0_0_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[19]
  PIN data_arrays_0_0_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[1]
  PIN data_arrays_0_0_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[20]
  PIN data_arrays_0_0_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[21]
  PIN data_arrays_0_0_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[22]
  PIN data_arrays_0_0_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[23]
  PIN data_arrays_0_0_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[24]
  PIN data_arrays_0_0_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[25]
  PIN data_arrays_0_0_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[26]
  PIN data_arrays_0_0_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[27]
  PIN data_arrays_0_0_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[28]
  PIN data_arrays_0_0_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[29]
  PIN data_arrays_0_0_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[2]
  PIN data_arrays_0_0_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[30]
  PIN data_arrays_0_0_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[31]
  PIN data_arrays_0_0_ext_ram_rdata0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[32]
  PIN data_arrays_0_0_ext_ram_rdata0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[33]
  PIN data_arrays_0_0_ext_ram_rdata0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[34]
  PIN data_arrays_0_0_ext_ram_rdata0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[35]
  PIN data_arrays_0_0_ext_ram_rdata0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[36]
  PIN data_arrays_0_0_ext_ram_rdata0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[37]
  PIN data_arrays_0_0_ext_ram_rdata0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[38]
  PIN data_arrays_0_0_ext_ram_rdata0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[39]
  PIN data_arrays_0_0_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[3]
  PIN data_arrays_0_0_ext_ram_rdata0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[40]
  PIN data_arrays_0_0_ext_ram_rdata0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[41]
  PIN data_arrays_0_0_ext_ram_rdata0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[42]
  PIN data_arrays_0_0_ext_ram_rdata0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[43]
  PIN data_arrays_0_0_ext_ram_rdata0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[44]
  PIN data_arrays_0_0_ext_ram_rdata0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[45]
  PIN data_arrays_0_0_ext_ram_rdata0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[46]
  PIN data_arrays_0_0_ext_ram_rdata0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[47]
  PIN data_arrays_0_0_ext_ram_rdata0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[48]
  PIN data_arrays_0_0_ext_ram_rdata0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[49]
  PIN data_arrays_0_0_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[4]
  PIN data_arrays_0_0_ext_ram_rdata0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[50]
  PIN data_arrays_0_0_ext_ram_rdata0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[51]
  PIN data_arrays_0_0_ext_ram_rdata0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[52]
  PIN data_arrays_0_0_ext_ram_rdata0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[53]
  PIN data_arrays_0_0_ext_ram_rdata0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[54]
  PIN data_arrays_0_0_ext_ram_rdata0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[55]
  PIN data_arrays_0_0_ext_ram_rdata0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[56]
  PIN data_arrays_0_0_ext_ram_rdata0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[57]
  PIN data_arrays_0_0_ext_ram_rdata0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[58]
  PIN data_arrays_0_0_ext_ram_rdata0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[59]
  PIN data_arrays_0_0_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[5]
  PIN data_arrays_0_0_ext_ram_rdata0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[60]
  PIN data_arrays_0_0_ext_ram_rdata0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[61]
  PIN data_arrays_0_0_ext_ram_rdata0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[62]
  PIN data_arrays_0_0_ext_ram_rdata0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[63]
  PIN data_arrays_0_0_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[6]
  PIN data_arrays_0_0_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[7]
  PIN data_arrays_0_0_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[8]
  PIN data_arrays_0_0_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[9]
  PIN data_arrays_0_0_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.760 4.000 904.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[0]
  PIN data_arrays_0_0_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.920 4.000 963.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[10]
  PIN data_arrays_0_0_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[11]
  PIN data_arrays_0_0_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 4.000 975.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[12]
  PIN data_arrays_0_0_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[13]
  PIN data_arrays_0_0_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.720 4.000 987.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[14]
  PIN data_arrays_0_0_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[15]
  PIN data_arrays_0_0_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 998.280 4.000 998.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[16]
  PIN data_arrays_0_0_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1004.400 4.000 1005.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[17]
  PIN data_arrays_0_0_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1010.520 4.000 1011.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[18]
  PIN data_arrays_0_0_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[19]
  PIN data_arrays_0_0_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[1]
  PIN data_arrays_0_0_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1022.080 4.000 1022.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[20]
  PIN data_arrays_0_0_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1028.200 4.000 1028.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[21]
  PIN data_arrays_0_0_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1034.320 4.000 1034.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[22]
  PIN data_arrays_0_0_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1039.760 4.000 1040.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[23]
  PIN data_arrays_0_0_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.880 4.000 1046.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[24]
  PIN data_arrays_0_0_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1052.000 4.000 1052.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[25]
  PIN data_arrays_0_0_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1058.120 4.000 1058.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[26]
  PIN data_arrays_0_0_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1063.560 4.000 1064.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[27]
  PIN data_arrays_0_0_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1069.680 4.000 1070.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[28]
  PIN data_arrays_0_0_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.800 4.000 1076.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[29]
  PIN data_arrays_0_0_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 915.320 4.000 915.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[2]
  PIN data_arrays_0_0_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[30]
  PIN data_arrays_0_0_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1087.360 4.000 1087.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[31]
  PIN data_arrays_0_0_ext_ram_rdata1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1093.480 4.000 1094.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[32]
  PIN data_arrays_0_0_ext_ram_rdata1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[33]
  PIN data_arrays_0_0_ext_ram_rdata1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[34]
  PIN data_arrays_0_0_ext_ram_rdata1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.160 4.000 1111.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[35]
  PIN data_arrays_0_0_ext_ram_rdata1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.280 4.000 1117.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[36]
  PIN data_arrays_0_0_ext_ram_rdata1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.720 4.000 1123.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[37]
  PIN data_arrays_0_0_ext_ram_rdata1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[38]
  PIN data_arrays_0_0_ext_ram_rdata1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1134.960 4.000 1135.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[39]
  PIN data_arrays_0_0_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[3]
  PIN data_arrays_0_0_ext_ram_rdata1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.080 4.000 1141.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[40]
  PIN data_arrays_0_0_ext_ram_rdata1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1146.520 4.000 1147.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[41]
  PIN data_arrays_0_0_ext_ram_rdata1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[42]
  PIN data_arrays_0_0_ext_ram_rdata1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1158.760 4.000 1159.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[43]
  PIN data_arrays_0_0_ext_ram_rdata1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1164.880 4.000 1165.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[44]
  PIN data_arrays_0_0_ext_ram_rdata1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1170.320 4.000 1170.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[45]
  PIN data_arrays_0_0_ext_ram_rdata1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[46]
  PIN data_arrays_0_0_ext_ram_rdata1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1182.560 4.000 1183.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[47]
  PIN data_arrays_0_0_ext_ram_rdata1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1188.000 4.000 1188.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[48]
  PIN data_arrays_0_0_ext_ram_rdata1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.120 4.000 1194.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[49]
  PIN data_arrays_0_0_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 927.560 4.000 928.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[4]
  PIN data_arrays_0_0_ext_ram_rdata1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 4.000 1200.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[50]
  PIN data_arrays_0_0_ext_ram_rdata1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1206.360 4.000 1206.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[51]
  PIN data_arrays_0_0_ext_ram_rdata1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1211.800 4.000 1212.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[52]
  PIN data_arrays_0_0_ext_ram_rdata1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.920 4.000 1218.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[53]
  PIN data_arrays_0_0_ext_ram_rdata1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.040 4.000 1224.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[54]
  PIN data_arrays_0_0_ext_ram_rdata1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1229.480 4.000 1230.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[55]
  PIN data_arrays_0_0_ext_ram_rdata1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1235.600 4.000 1236.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[56]
  PIN data_arrays_0_0_ext_ram_rdata1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.720 4.000 1242.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[57]
  PIN data_arrays_0_0_ext_ram_rdata1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[58]
  PIN data_arrays_0_0_ext_ram_rdata1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1253.280 4.000 1253.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[59]
  PIN data_arrays_0_0_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.000 4.000 933.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[5]
  PIN data_arrays_0_0_ext_ram_rdata1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1259.400 4.000 1260.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[60]
  PIN data_arrays_0_0_ext_ram_rdata1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1265.520 4.000 1266.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[61]
  PIN data_arrays_0_0_ext_ram_rdata1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.960 4.000 1271.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[62]
  PIN data_arrays_0_0_ext_ram_rdata1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1277.080 4.000 1277.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[63]
  PIN data_arrays_0_0_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[6]
  PIN data_arrays_0_0_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[7]
  PIN data_arrays_0_0_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 951.360 4.000 951.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[8]
  PIN data_arrays_0_0_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 956.800 4.000 957.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[9]
  PIN data_arrays_0_0_ext_ram_rdata2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 1792.280 104.790 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[0]
  PIN data_arrays_0_0_ext_ram_rdata2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 1792.280 136.990 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[10]
  PIN data_arrays_0_0_ext_ram_rdata2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 1792.280 140.210 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[11]
  PIN data_arrays_0_0_ext_ram_rdata2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 1792.280 143.430 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[12]
  PIN data_arrays_0_0_ext_ram_rdata2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 1792.280 146.650 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[13]
  PIN data_arrays_0_0_ext_ram_rdata2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 1792.280 149.870 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[14]
  PIN data_arrays_0_0_ext_ram_rdata2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 1792.280 153.090 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[15]
  PIN data_arrays_0_0_ext_ram_rdata2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 1792.280 156.310 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[16]
  PIN data_arrays_0_0_ext_ram_rdata2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 1792.280 159.530 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[17]
  PIN data_arrays_0_0_ext_ram_rdata2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 1792.280 162.750 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[18]
  PIN data_arrays_0_0_ext_ram_rdata2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 1792.280 166.430 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[19]
  PIN data_arrays_0_0_ext_ram_rdata2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 1792.280 108.010 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[1]
  PIN data_arrays_0_0_ext_ram_rdata2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 1792.280 169.650 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[20]
  PIN data_arrays_0_0_ext_ram_rdata2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 1792.280 172.870 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[21]
  PIN data_arrays_0_0_ext_ram_rdata2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 1792.280 176.090 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[22]
  PIN data_arrays_0_0_ext_ram_rdata2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 1792.280 179.310 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[23]
  PIN data_arrays_0_0_ext_ram_rdata2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 1792.280 182.530 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[24]
  PIN data_arrays_0_0_ext_ram_rdata2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 1792.280 185.750 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[25]
  PIN data_arrays_0_0_ext_ram_rdata2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 1792.280 188.970 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[26]
  PIN data_arrays_0_0_ext_ram_rdata2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 1792.280 192.190 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[27]
  PIN data_arrays_0_0_ext_ram_rdata2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 1792.280 195.410 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[28]
  PIN data_arrays_0_0_ext_ram_rdata2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 1792.280 198.630 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[29]
  PIN data_arrays_0_0_ext_ram_rdata2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 1792.280 111.230 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[2]
  PIN data_arrays_0_0_ext_ram_rdata2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 1792.280 201.850 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[30]
  PIN data_arrays_0_0_ext_ram_rdata2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 1792.280 205.070 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[31]
  PIN data_arrays_0_0_ext_ram_rdata2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 1792.280 208.290 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[32]
  PIN data_arrays_0_0_ext_ram_rdata2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 1792.280 211.510 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[33]
  PIN data_arrays_0_0_ext_ram_rdata2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 1792.280 214.730 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[34]
  PIN data_arrays_0_0_ext_ram_rdata2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 1792.280 217.950 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[35]
  PIN data_arrays_0_0_ext_ram_rdata2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 1792.280 221.170 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[36]
  PIN data_arrays_0_0_ext_ram_rdata2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 1792.280 224.390 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[37]
  PIN data_arrays_0_0_ext_ram_rdata2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 1792.280 227.610 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[38]
  PIN data_arrays_0_0_ext_ram_rdata2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 1792.280 230.830 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[39]
  PIN data_arrays_0_0_ext_ram_rdata2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 1792.280 114.450 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[3]
  PIN data_arrays_0_0_ext_ram_rdata2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 1792.280 234.050 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[40]
  PIN data_arrays_0_0_ext_ram_rdata2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 1792.280 237.270 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[41]
  PIN data_arrays_0_0_ext_ram_rdata2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 1792.280 240.490 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[42]
  PIN data_arrays_0_0_ext_ram_rdata2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 1792.280 243.710 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[43]
  PIN data_arrays_0_0_ext_ram_rdata2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 1792.280 246.930 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[44]
  PIN data_arrays_0_0_ext_ram_rdata2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 1792.280 250.150 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[45]
  PIN data_arrays_0_0_ext_ram_rdata2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 1792.280 253.370 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[46]
  PIN data_arrays_0_0_ext_ram_rdata2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 1792.280 256.590 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[47]
  PIN data_arrays_0_0_ext_ram_rdata2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 1792.280 259.810 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[48]
  PIN data_arrays_0_0_ext_ram_rdata2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 1792.280 263.030 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[49]
  PIN data_arrays_0_0_ext_ram_rdata2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 1792.280 117.670 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[4]
  PIN data_arrays_0_0_ext_ram_rdata2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 1792.280 266.250 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[50]
  PIN data_arrays_0_0_ext_ram_rdata2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 1792.280 269.470 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[51]
  PIN data_arrays_0_0_ext_ram_rdata2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 1792.280 272.690 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[52]
  PIN data_arrays_0_0_ext_ram_rdata2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 1792.280 275.910 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[53]
  PIN data_arrays_0_0_ext_ram_rdata2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 1792.280 279.130 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[54]
  PIN data_arrays_0_0_ext_ram_rdata2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 1792.280 282.350 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[55]
  PIN data_arrays_0_0_ext_ram_rdata2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 1792.280 285.570 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[56]
  PIN data_arrays_0_0_ext_ram_rdata2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 1792.280 288.790 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[57]
  PIN data_arrays_0_0_ext_ram_rdata2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 1792.280 292.010 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[58]
  PIN data_arrays_0_0_ext_ram_rdata2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 1792.280 295.230 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[59]
  PIN data_arrays_0_0_ext_ram_rdata2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 1792.280 120.890 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[5]
  PIN data_arrays_0_0_ext_ram_rdata2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 1792.280 298.450 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[60]
  PIN data_arrays_0_0_ext_ram_rdata2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 1792.280 301.670 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[61]
  PIN data_arrays_0_0_ext_ram_rdata2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 1792.280 304.890 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[62]
  PIN data_arrays_0_0_ext_ram_rdata2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 1792.280 308.110 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[63]
  PIN data_arrays_0_0_ext_ram_rdata2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 1792.280 124.110 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[6]
  PIN data_arrays_0_0_ext_ram_rdata2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 1792.280 127.330 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[7]
  PIN data_arrays_0_0_ext_ram_rdata2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 1792.280 130.550 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[8]
  PIN data_arrays_0_0_ext_ram_rdata2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 1792.280 133.770 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[9]
  PIN data_arrays_0_0_ext_ram_rdata3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 1792.280 1299.410 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[0]
  PIN data_arrays_0_0_ext_ram_rdata3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.790 1792.280 1332.070 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[10]
  PIN data_arrays_0_0_ext_ram_rdata3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.010 1792.280 1335.290 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[11]
  PIN data_arrays_0_0_ext_ram_rdata3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.230 1792.280 1338.510 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[12]
  PIN data_arrays_0_0_ext_ram_rdata3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.450 1792.280 1341.730 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[13]
  PIN data_arrays_0_0_ext_ram_rdata3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.670 1792.280 1344.950 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[14]
  PIN data_arrays_0_0_ext_ram_rdata3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.890 1792.280 1348.170 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[15]
  PIN data_arrays_0_0_ext_ram_rdata3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.110 1792.280 1351.390 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[16]
  PIN data_arrays_0_0_ext_ram_rdata3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.330 1792.280 1354.610 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[17]
  PIN data_arrays_0_0_ext_ram_rdata3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.550 1792.280 1357.830 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[18]
  PIN data_arrays_0_0_ext_ram_rdata3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 1792.280 1361.050 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[19]
  PIN data_arrays_0_0_ext_ram_rdata3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.810 1792.280 1303.090 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[1]
  PIN data_arrays_0_0_ext_ram_rdata3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 1792.280 1364.270 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[20]
  PIN data_arrays_0_0_ext_ram_rdata3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.210 1792.280 1367.490 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[21]
  PIN data_arrays_0_0_ext_ram_rdata3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 1792.280 1370.710 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[22]
  PIN data_arrays_0_0_ext_ram_rdata3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.650 1792.280 1373.930 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[23]
  PIN data_arrays_0_0_ext_ram_rdata3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.870 1792.280 1377.150 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[24]
  PIN data_arrays_0_0_ext_ram_rdata3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 1792.280 1380.370 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[25]
  PIN data_arrays_0_0_ext_ram_rdata3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.310 1792.280 1383.590 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[26]
  PIN data_arrays_0_0_ext_ram_rdata3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.530 1792.280 1386.810 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[27]
  PIN data_arrays_0_0_ext_ram_rdata3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.750 1792.280 1390.030 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[28]
  PIN data_arrays_0_0_ext_ram_rdata3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.970 1792.280 1393.250 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[29]
  PIN data_arrays_0_0_ext_ram_rdata3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.030 1792.280 1306.310 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[2]
  PIN data_arrays_0_0_ext_ram_rdata3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.190 1792.280 1396.470 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[30]
  PIN data_arrays_0_0_ext_ram_rdata3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.410 1792.280 1399.690 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[31]
  PIN data_arrays_0_0_ext_ram_rdata3[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.630 1792.280 1402.910 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[32]
  PIN data_arrays_0_0_ext_ram_rdata3[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 1792.280 1406.130 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[33]
  PIN data_arrays_0_0_ext_ram_rdata3[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.070 1792.280 1409.350 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[34]
  PIN data_arrays_0_0_ext_ram_rdata3[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.290 1792.280 1412.570 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[35]
  PIN data_arrays_0_0_ext_ram_rdata3[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.510 1792.280 1415.790 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[36]
  PIN data_arrays_0_0_ext_ram_rdata3[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 1792.280 1419.010 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[37]
  PIN data_arrays_0_0_ext_ram_rdata3[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.950 1792.280 1422.230 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[38]
  PIN data_arrays_0_0_ext_ram_rdata3[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.170 1792.280 1425.450 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[39]
  PIN data_arrays_0_0_ext_ram_rdata3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.250 1792.280 1309.530 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[3]
  PIN data_arrays_0_0_ext_ram_rdata3[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.390 1792.280 1428.670 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[40]
  PIN data_arrays_0_0_ext_ram_rdata3[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.610 1792.280 1431.890 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[41]
  PIN data_arrays_0_0_ext_ram_rdata3[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.830 1792.280 1435.110 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[42]
  PIN data_arrays_0_0_ext_ram_rdata3[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.050 1792.280 1438.330 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[43]
  PIN data_arrays_0_0_ext_ram_rdata3[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.270 1792.280 1441.550 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[44]
  PIN data_arrays_0_0_ext_ram_rdata3[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.490 1792.280 1444.770 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[45]
  PIN data_arrays_0_0_ext_ram_rdata3[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.710 1792.280 1447.990 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[46]
  PIN data_arrays_0_0_ext_ram_rdata3[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.930 1792.280 1451.210 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[47]
  PIN data_arrays_0_0_ext_ram_rdata3[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.150 1792.280 1454.430 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[48]
  PIN data_arrays_0_0_ext_ram_rdata3[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.370 1792.280 1457.650 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[49]
  PIN data_arrays_0_0_ext_ram_rdata3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.470 1792.280 1312.750 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[4]
  PIN data_arrays_0_0_ext_ram_rdata3[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.590 1792.280 1460.870 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[50]
  PIN data_arrays_0_0_ext_ram_rdata3[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 1792.280 1464.550 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[51]
  PIN data_arrays_0_0_ext_ram_rdata3[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.490 1792.280 1467.770 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[52]
  PIN data_arrays_0_0_ext_ram_rdata3[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.710 1792.280 1470.990 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[53]
  PIN data_arrays_0_0_ext_ram_rdata3[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 1792.280 1474.210 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[54]
  PIN data_arrays_0_0_ext_ram_rdata3[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.150 1792.280 1477.430 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[55]
  PIN data_arrays_0_0_ext_ram_rdata3[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.370 1792.280 1480.650 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[56]
  PIN data_arrays_0_0_ext_ram_rdata3[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.590 1792.280 1483.870 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[57]
  PIN data_arrays_0_0_ext_ram_rdata3[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.810 1792.280 1487.090 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[58]
  PIN data_arrays_0_0_ext_ram_rdata3[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.030 1792.280 1490.310 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[59]
  PIN data_arrays_0_0_ext_ram_rdata3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.690 1792.280 1315.970 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[5]
  PIN data_arrays_0_0_ext_ram_rdata3[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.250 1792.280 1493.530 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[60]
  PIN data_arrays_0_0_ext_ram_rdata3[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.470 1792.280 1496.750 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[61]
  PIN data_arrays_0_0_ext_ram_rdata3[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 1792.280 1499.970 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[62]
  PIN data_arrays_0_0_ext_ram_rdata3[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.910 1792.280 1503.190 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[63]
  PIN data_arrays_0_0_ext_ram_rdata3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.910 1792.280 1319.190 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[6]
  PIN data_arrays_0_0_ext_ram_rdata3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.130 1792.280 1322.410 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[7]
  PIN data_arrays_0_0_ext_ram_rdata3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.350 1792.280 1325.630 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[8]
  PIN data_arrays_0_0_ext_ram_rdata3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.570 1792.280 1328.850 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[9]
  PIN data_arrays_0_0_ext_ram_wdata0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[0]
  PIN data_arrays_0_0_ext_ram_wdata0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[10]
  PIN data_arrays_0_0_ext_ram_wdata0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[11]
  PIN data_arrays_0_0_ext_ram_wdata0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.080 4.000 512.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[12]
  PIN data_arrays_0_0_ext_ram_wdata0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[13]
  PIN data_arrays_0_0_ext_ram_wdata0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[14]
  PIN data_arrays_0_0_ext_ram_wdata0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[15]
  PIN data_arrays_0_0_ext_ram_wdata0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[16]
  PIN data_arrays_0_0_ext_ram_wdata0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[17]
  PIN data_arrays_0_0_ext_ram_wdata0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[18]
  PIN data_arrays_0_0_ext_ram_wdata0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[19]
  PIN data_arrays_0_0_ext_ram_wdata0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.800 4.000 447.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[1]
  PIN data_arrays_0_0_ext_ram_wdata0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[20]
  PIN data_arrays_0_0_ext_ram_wdata0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[21]
  PIN data_arrays_0_0_ext_ram_wdata0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[22]
  PIN data_arrays_0_0_ext_ram_wdata0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 577.360 4.000 577.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[23]
  PIN data_arrays_0_0_ext_ram_wdata0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[24]
  PIN data_arrays_0_0_ext_ram_wdata0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[25]
  PIN data_arrays_0_0_ext_ram_wdata0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[26]
  PIN data_arrays_0_0_ext_ram_wdata0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[27]
  PIN data_arrays_0_0_ext_ram_wdata0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[28]
  PIN data_arrays_0_0_ext_ram_wdata0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[29]
  PIN data_arrays_0_0_ext_ram_wdata0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[2]
  PIN data_arrays_0_0_ext_ram_wdata0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[30]
  PIN data_arrays_0_0_ext_ram_wdata0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.960 4.000 625.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[31]
  PIN data_arrays_0_0_ext_ram_wdata0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[32]
  PIN data_arrays_0_0_ext_ram_wdata0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[33]
  PIN data_arrays_0_0_ext_ram_wdata0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[34]
  PIN data_arrays_0_0_ext_ram_wdata0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[35]
  PIN data_arrays_0_0_ext_ram_wdata0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.880 4.000 655.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[36]
  PIN data_arrays_0_0_ext_ram_wdata0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[37]
  PIN data_arrays_0_0_ext_ram_wdata0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[38]
  PIN data_arrays_0_0_ext_ram_wdata0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 672.560 4.000 673.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[39]
  PIN data_arrays_0_0_ext_ram_wdata0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[3]
  PIN data_arrays_0_0_ext_ram_wdata0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[40]
  PIN data_arrays_0_0_ext_ram_wdata0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[41]
  PIN data_arrays_0_0_ext_ram_wdata0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[42]
  PIN data_arrays_0_0_ext_ram_wdata0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[43]
  PIN data_arrays_0_0_ext_ram_wdata0[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[44]
  PIN data_arrays_0_0_ext_ram_wdata0[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.920 4.000 708.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[45]
  PIN data_arrays_0_0_ext_ram_wdata0[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[46]
  PIN data_arrays_0_0_ext_ram_wdata0[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[47]
  PIN data_arrays_0_0_ext_ram_wdata0[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[48]
  PIN data_arrays_0_0_ext_ram_wdata0[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[49]
  PIN data_arrays_0_0_ext_ram_wdata0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[4]
  PIN data_arrays_0_0_ext_ram_wdata0[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[50]
  PIN data_arrays_0_0_ext_ram_wdata0[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[51]
  PIN data_arrays_0_0_ext_ram_wdata0[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[52]
  PIN data_arrays_0_0_ext_ram_wdata0[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[53]
  PIN data_arrays_0_0_ext_ram_wdata0[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[54]
  PIN data_arrays_0_0_ext_ram_wdata0[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 767.080 4.000 767.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[55]
  PIN data_arrays_0_0_ext_ram_wdata0[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[56]
  PIN data_arrays_0_0_ext_ram_wdata0[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[57]
  PIN data_arrays_0_0_ext_ram_wdata0[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[58]
  PIN data_arrays_0_0_ext_ram_wdata0[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.880 4.000 791.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[59]
  PIN data_arrays_0_0_ext_ram_wdata0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[5]
  PIN data_arrays_0_0_ext_ram_wdata0[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[60]
  PIN data_arrays_0_0_ext_ram_wdata0[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.120 4.000 803.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[61]
  PIN data_arrays_0_0_ext_ram_wdata0[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 808.560 4.000 809.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[62]
  PIN data_arrays_0_0_ext_ram_wdata0[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[63]
  PIN data_arrays_0_0_ext_ram_wdata0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[6]
  PIN data_arrays_0_0_ext_ram_wdata0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[7]
  PIN data_arrays_0_0_ext_ram_wdata0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[8]
  PIN data_arrays_0_0_ext_ram_wdata0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 494.400 4.000 495.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata0[9]
  PIN data_arrays_0_0_ext_ram_wdata1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1336.240 4.000 1336.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[0]
  PIN data_arrays_0_0_ext_ram_wdata1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1396.080 4.000 1396.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[10]
  PIN data_arrays_0_0_ext_ram_wdata1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1401.520 4.000 1402.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[11]
  PIN data_arrays_0_0_ext_ram_wdata1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[12]
  PIN data_arrays_0_0_ext_ram_wdata1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1413.760 4.000 1414.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[13]
  PIN data_arrays_0_0_ext_ram_wdata1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1419.200 4.000 1419.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[14]
  PIN data_arrays_0_0_ext_ram_wdata1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1425.320 4.000 1425.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[15]
  PIN data_arrays_0_0_ext_ram_wdata1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[16]
  PIN data_arrays_0_0_ext_ram_wdata1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1437.560 4.000 1438.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[17]
  PIN data_arrays_0_0_ext_ram_wdata1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1443.000 4.000 1443.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[18]
  PIN data_arrays_0_0_ext_ram_wdata1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1449.120 4.000 1449.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[19]
  PIN data_arrays_0_0_ext_ram_wdata1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1342.360 4.000 1342.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[1]
  PIN data_arrays_0_0_ext_ram_wdata1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[20]
  PIN data_arrays_0_0_ext_ram_wdata1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1460.680 4.000 1461.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[21]
  PIN data_arrays_0_0_ext_ram_wdata1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1466.800 4.000 1467.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[22]
  PIN data_arrays_0_0_ext_ram_wdata1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.920 4.000 1473.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[23]
  PIN data_arrays_0_0_ext_ram_wdata1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.040 4.000 1479.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[24]
  PIN data_arrays_0_0_ext_ram_wdata1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1484.480 4.000 1485.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[25]
  PIN data_arrays_0_0_ext_ram_wdata1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1490.600 4.000 1491.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[26]
  PIN data_arrays_0_0_ext_ram_wdata1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1496.720 4.000 1497.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[27]
  PIN data_arrays_0_0_ext_ram_wdata1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1502.840 4.000 1503.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[28]
  PIN data_arrays_0_0_ext_ram_wdata1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1508.280 4.000 1508.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[29]
  PIN data_arrays_0_0_ext_ram_wdata1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1348.480 4.000 1349.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[2]
  PIN data_arrays_0_0_ext_ram_wdata1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1514.400 4.000 1515.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[30]
  PIN data_arrays_0_0_ext_ram_wdata1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1520.520 4.000 1521.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[31]
  PIN data_arrays_0_0_ext_ram_wdata1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1525.960 4.000 1526.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[32]
  PIN data_arrays_0_0_ext_ram_wdata1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1532.080 4.000 1532.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[33]
  PIN data_arrays_0_0_ext_ram_wdata1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1538.200 4.000 1538.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[34]
  PIN data_arrays_0_0_ext_ram_wdata1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1544.320 4.000 1544.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[35]
  PIN data_arrays_0_0_ext_ram_wdata1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1549.760 4.000 1550.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[36]
  PIN data_arrays_0_0_ext_ram_wdata1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1555.880 4.000 1556.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[37]
  PIN data_arrays_0_0_ext_ram_wdata1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1562.000 4.000 1562.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[38]
  PIN data_arrays_0_0_ext_ram_wdata1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1567.440 4.000 1568.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[39]
  PIN data_arrays_0_0_ext_ram_wdata1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1354.600 4.000 1355.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[3]
  PIN data_arrays_0_0_ext_ram_wdata1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1573.560 4.000 1574.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[40]
  PIN data_arrays_0_0_ext_ram_wdata1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1579.680 4.000 1580.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[41]
  PIN data_arrays_0_0_ext_ram_wdata1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1585.800 4.000 1586.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[42]
  PIN data_arrays_0_0_ext_ram_wdata1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1591.240 4.000 1591.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[43]
  PIN data_arrays_0_0_ext_ram_wdata1[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1597.360 4.000 1597.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[44]
  PIN data_arrays_0_0_ext_ram_wdata1[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1603.480 4.000 1604.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[45]
  PIN data_arrays_0_0_ext_ram_wdata1[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1608.920 4.000 1609.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[46]
  PIN data_arrays_0_0_ext_ram_wdata1[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1615.040 4.000 1615.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[47]
  PIN data_arrays_0_0_ext_ram_wdata1[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1621.160 4.000 1621.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[48]
  PIN data_arrays_0_0_ext_ram_wdata1[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1627.280 4.000 1627.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[49]
  PIN data_arrays_0_0_ext_ram_wdata1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[4]
  PIN data_arrays_0_0_ext_ram_wdata1[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1632.720 4.000 1633.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[50]
  PIN data_arrays_0_0_ext_ram_wdata1[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.840 4.000 1639.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[51]
  PIN data_arrays_0_0_ext_ram_wdata1[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1644.960 4.000 1645.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[52]
  PIN data_arrays_0_0_ext_ram_wdata1[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1651.080 4.000 1651.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[53]
  PIN data_arrays_0_0_ext_ram_wdata1[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1656.520 4.000 1657.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[54]
  PIN data_arrays_0_0_ext_ram_wdata1[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1662.640 4.000 1663.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[55]
  PIN data_arrays_0_0_ext_ram_wdata1[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1668.760 4.000 1669.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[56]
  PIN data_arrays_0_0_ext_ram_wdata1[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1674.200 4.000 1674.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[57]
  PIN data_arrays_0_0_ext_ram_wdata1[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1680.320 4.000 1680.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[58]
  PIN data_arrays_0_0_ext_ram_wdata1[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1686.440 4.000 1687.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[59]
  PIN data_arrays_0_0_ext_ram_wdata1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.160 4.000 1366.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[5]
  PIN data_arrays_0_0_ext_ram_wdata1[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1692.560 4.000 1693.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[60]
  PIN data_arrays_0_0_ext_ram_wdata1[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1698.000 4.000 1698.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[61]
  PIN data_arrays_0_0_ext_ram_wdata1[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1704.120 4.000 1704.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[62]
  PIN data_arrays_0_0_ext_ram_wdata1[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[63]
  PIN data_arrays_0_0_ext_ram_wdata1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1372.280 4.000 1372.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[6]
  PIN data_arrays_0_0_ext_ram_wdata1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.720 4.000 1378.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[7]
  PIN data_arrays_0_0_ext_ram_wdata1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[8]
  PIN data_arrays_0_0_ext_ram_wdata1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1389.960 4.000 1390.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata1[9]
  PIN data_arrays_0_0_ext_ram_wdata2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 1792.280 340.770 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[0]
  PIN data_arrays_0_0_ext_ram_wdata2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 1792.280 372.970 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[10]
  PIN data_arrays_0_0_ext_ram_wdata2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 1792.280 376.190 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[11]
  PIN data_arrays_0_0_ext_ram_wdata2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 1792.280 379.410 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[12]
  PIN data_arrays_0_0_ext_ram_wdata2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 1792.280 382.630 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[13]
  PIN data_arrays_0_0_ext_ram_wdata2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 1792.280 385.850 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[14]
  PIN data_arrays_0_0_ext_ram_wdata2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 1792.280 389.070 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[15]
  PIN data_arrays_0_0_ext_ram_wdata2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 1792.280 392.290 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[16]
  PIN data_arrays_0_0_ext_ram_wdata2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 1792.280 395.510 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[17]
  PIN data_arrays_0_0_ext_ram_wdata2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 1792.280 398.730 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[18]
  PIN data_arrays_0_0_ext_ram_wdata2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 1792.280 401.950 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[19]
  PIN data_arrays_0_0_ext_ram_wdata2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 1792.280 343.990 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[1]
  PIN data_arrays_0_0_ext_ram_wdata2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 1792.280 405.170 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[20]
  PIN data_arrays_0_0_ext_ram_wdata2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 1792.280 408.390 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[21]
  PIN data_arrays_0_0_ext_ram_wdata2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 1792.280 411.610 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[22]
  PIN data_arrays_0_0_ext_ram_wdata2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 1792.280 414.830 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[23]
  PIN data_arrays_0_0_ext_ram_wdata2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 1792.280 418.050 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[24]
  PIN data_arrays_0_0_ext_ram_wdata2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 1792.280 421.270 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[25]
  PIN data_arrays_0_0_ext_ram_wdata2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 1792.280 424.490 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[26]
  PIN data_arrays_0_0_ext_ram_wdata2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 1792.280 427.710 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[27]
  PIN data_arrays_0_0_ext_ram_wdata2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 1792.280 430.930 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[28]
  PIN data_arrays_0_0_ext_ram_wdata2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 1792.280 434.150 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[29]
  PIN data_arrays_0_0_ext_ram_wdata2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 1792.280 347.210 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[2]
  PIN data_arrays_0_0_ext_ram_wdata2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 1792.280 437.370 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[30]
  PIN data_arrays_0_0_ext_ram_wdata2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 1792.280 440.590 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[31]
  PIN data_arrays_0_0_ext_ram_wdata2[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 1792.280 443.810 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[32]
  PIN data_arrays_0_0_ext_ram_wdata2[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 1792.280 447.030 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[33]
  PIN data_arrays_0_0_ext_ram_wdata2[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 1792.280 450.250 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[34]
  PIN data_arrays_0_0_ext_ram_wdata2[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 1792.280 453.470 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[35]
  PIN data_arrays_0_0_ext_ram_wdata2[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 1792.280 456.690 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[36]
  PIN data_arrays_0_0_ext_ram_wdata2[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 1792.280 459.910 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[37]
  PIN data_arrays_0_0_ext_ram_wdata2[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 1792.280 463.130 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[38]
  PIN data_arrays_0_0_ext_ram_wdata2[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 1792.280 466.350 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[39]
  PIN data_arrays_0_0_ext_ram_wdata2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 1792.280 350.430 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[3]
  PIN data_arrays_0_0_ext_ram_wdata2[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 1792.280 469.570 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[40]
  PIN data_arrays_0_0_ext_ram_wdata2[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 1792.280 472.790 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[41]
  PIN data_arrays_0_0_ext_ram_wdata2[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 1792.280 476.010 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[42]
  PIN data_arrays_0_0_ext_ram_wdata2[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 1792.280 479.230 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[43]
  PIN data_arrays_0_0_ext_ram_wdata2[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 1792.280 482.450 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[44]
  PIN data_arrays_0_0_ext_ram_wdata2[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 1792.280 485.670 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[45]
  PIN data_arrays_0_0_ext_ram_wdata2[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 1792.280 489.350 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[46]
  PIN data_arrays_0_0_ext_ram_wdata2[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 1792.280 492.570 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[47]
  PIN data_arrays_0_0_ext_ram_wdata2[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 1792.280 495.790 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[48]
  PIN data_arrays_0_0_ext_ram_wdata2[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 1792.280 499.010 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[49]
  PIN data_arrays_0_0_ext_ram_wdata2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 1792.280 353.650 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[4]
  PIN data_arrays_0_0_ext_ram_wdata2[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 1792.280 502.230 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[50]
  PIN data_arrays_0_0_ext_ram_wdata2[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 1792.280 505.450 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[51]
  PIN data_arrays_0_0_ext_ram_wdata2[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 1792.280 508.670 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[52]
  PIN data_arrays_0_0_ext_ram_wdata2[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 1792.280 511.890 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[53]
  PIN data_arrays_0_0_ext_ram_wdata2[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 1792.280 515.110 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[54]
  PIN data_arrays_0_0_ext_ram_wdata2[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 1792.280 518.330 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[55]
  PIN data_arrays_0_0_ext_ram_wdata2[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 1792.280 521.550 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[56]
  PIN data_arrays_0_0_ext_ram_wdata2[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 1792.280 524.770 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[57]
  PIN data_arrays_0_0_ext_ram_wdata2[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 1792.280 527.990 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[58]
  PIN data_arrays_0_0_ext_ram_wdata2[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 1792.280 531.210 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[59]
  PIN data_arrays_0_0_ext_ram_wdata2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 1792.280 356.870 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[5]
  PIN data_arrays_0_0_ext_ram_wdata2[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 1792.280 534.430 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[60]
  PIN data_arrays_0_0_ext_ram_wdata2[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 1792.280 537.650 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[61]
  PIN data_arrays_0_0_ext_ram_wdata2[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 1792.280 540.870 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[62]
  PIN data_arrays_0_0_ext_ram_wdata2[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 1792.280 544.090 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[63]
  PIN data_arrays_0_0_ext_ram_wdata2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 1792.280 360.090 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[6]
  PIN data_arrays_0_0_ext_ram_wdata2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 1792.280 363.310 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[7]
  PIN data_arrays_0_0_ext_ram_wdata2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 1792.280 366.530 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[8]
  PIN data_arrays_0_0_ext_ram_wdata2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 1792.280 369.750 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata2[9]
  PIN data_arrays_0_0_ext_ram_wdata3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.110 1792.280 1535.390 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[0]
  PIN data_arrays_0_0_ext_ram_wdata3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.310 1792.280 1567.590 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[10]
  PIN data_arrays_0_0_ext_ram_wdata3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.530 1792.280 1570.810 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[11]
  PIN data_arrays_0_0_ext_ram_wdata3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.750 1792.280 1574.030 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[12]
  PIN data_arrays_0_0_ext_ram_wdata3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.970 1792.280 1577.250 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[13]
  PIN data_arrays_0_0_ext_ram_wdata3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.190 1792.280 1580.470 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[14]
  PIN data_arrays_0_0_ext_ram_wdata3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.410 1792.280 1583.690 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[15]
  PIN data_arrays_0_0_ext_ram_wdata3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.630 1792.280 1586.910 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[16]
  PIN data_arrays_0_0_ext_ram_wdata3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.850 1792.280 1590.130 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[17]
  PIN data_arrays_0_0_ext_ram_wdata3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.070 1792.280 1593.350 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[18]
  PIN data_arrays_0_0_ext_ram_wdata3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.290 1792.280 1596.570 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[19]
  PIN data_arrays_0_0_ext_ram_wdata3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.330 1792.280 1538.610 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[1]
  PIN data_arrays_0_0_ext_ram_wdata3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.510 1792.280 1599.790 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[20]
  PIN data_arrays_0_0_ext_ram_wdata3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.730 1792.280 1603.010 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[21]
  PIN data_arrays_0_0_ext_ram_wdata3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.950 1792.280 1606.230 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[22]
  PIN data_arrays_0_0_ext_ram_wdata3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.170 1792.280 1609.450 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[23]
  PIN data_arrays_0_0_ext_ram_wdata3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.390 1792.280 1612.670 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[24]
  PIN data_arrays_0_0_ext_ram_wdata3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.610 1792.280 1615.890 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[25]
  PIN data_arrays_0_0_ext_ram_wdata3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.830 1792.280 1619.110 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[26]
  PIN data_arrays_0_0_ext_ram_wdata3[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.050 1792.280 1622.330 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[27]
  PIN data_arrays_0_0_ext_ram_wdata3[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 1792.280 1626.010 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[28]
  PIN data_arrays_0_0_ext_ram_wdata3[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.950 1792.280 1629.230 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[29]
  PIN data_arrays_0_0_ext_ram_wdata3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.550 1792.280 1541.830 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[2]
  PIN data_arrays_0_0_ext_ram_wdata3[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.170 1792.280 1632.450 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[30]
  PIN data_arrays_0_0_ext_ram_wdata3[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.390 1792.280 1635.670 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[31]
  PIN data_arrays_0_0_ext_ram_wdata3[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.610 1792.280 1638.890 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[32]
  PIN data_arrays_0_0_ext_ram_wdata3[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.830 1792.280 1642.110 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[33]
  PIN data_arrays_0_0_ext_ram_wdata3[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.050 1792.280 1645.330 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[34]
  PIN data_arrays_0_0_ext_ram_wdata3[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.270 1792.280 1648.550 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[35]
  PIN data_arrays_0_0_ext_ram_wdata3[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.490 1792.280 1651.770 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[36]
  PIN data_arrays_0_0_ext_ram_wdata3[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.710 1792.280 1654.990 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[37]
  PIN data_arrays_0_0_ext_ram_wdata3[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.930 1792.280 1658.210 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[38]
  PIN data_arrays_0_0_ext_ram_wdata3[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.150 1792.280 1661.430 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[39]
  PIN data_arrays_0_0_ext_ram_wdata3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.770 1792.280 1545.050 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[3]
  PIN data_arrays_0_0_ext_ram_wdata3[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.370 1792.280 1664.650 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[40]
  PIN data_arrays_0_0_ext_ram_wdata3[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 1792.280 1667.870 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[41]
  PIN data_arrays_0_0_ext_ram_wdata3[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.810 1792.280 1671.090 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[42]
  PIN data_arrays_0_0_ext_ram_wdata3[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.030 1792.280 1674.310 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[43]
  PIN data_arrays_0_0_ext_ram_wdata3[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.250 1792.280 1677.530 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[44]
  PIN data_arrays_0_0_ext_ram_wdata3[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.470 1792.280 1680.750 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[45]
  PIN data_arrays_0_0_ext_ram_wdata3[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.690 1792.280 1683.970 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[46]
  PIN data_arrays_0_0_ext_ram_wdata3[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.910 1792.280 1687.190 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[47]
  PIN data_arrays_0_0_ext_ram_wdata3[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.130 1792.280 1690.410 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[48]
  PIN data_arrays_0_0_ext_ram_wdata3[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.350 1792.280 1693.630 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[49]
  PIN data_arrays_0_0_ext_ram_wdata3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.990 1792.280 1548.270 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[4]
  PIN data_arrays_0_0_ext_ram_wdata3[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.570 1792.280 1696.850 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[50]
  PIN data_arrays_0_0_ext_ram_wdata3[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.790 1792.280 1700.070 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[51]
  PIN data_arrays_0_0_ext_ram_wdata3[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.010 1792.280 1703.290 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[52]
  PIN data_arrays_0_0_ext_ram_wdata3[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.230 1792.280 1706.510 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[53]
  PIN data_arrays_0_0_ext_ram_wdata3[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.450 1792.280 1709.730 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[54]
  PIN data_arrays_0_0_ext_ram_wdata3[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.670 1792.280 1712.950 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[55]
  PIN data_arrays_0_0_ext_ram_wdata3[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.890 1792.280 1716.170 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[56]
  PIN data_arrays_0_0_ext_ram_wdata3[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.110 1792.280 1719.390 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[57]
  PIN data_arrays_0_0_ext_ram_wdata3[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.330 1792.280 1722.610 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[58]
  PIN data_arrays_0_0_ext_ram_wdata3[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.550 1792.280 1725.830 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[59]
  PIN data_arrays_0_0_ext_ram_wdata3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.210 1792.280 1551.490 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[5]
  PIN data_arrays_0_0_ext_ram_wdata3[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.770 1792.280 1729.050 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[60]
  PIN data_arrays_0_0_ext_ram_wdata3[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.990 1792.280 1732.270 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[61]
  PIN data_arrays_0_0_ext_ram_wdata3[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.210 1792.280 1735.490 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[62]
  PIN data_arrays_0_0_ext_ram_wdata3[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.430 1792.280 1738.710 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[63]
  PIN data_arrays_0_0_ext_ram_wdata3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.430 1792.280 1554.710 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[6]
  PIN data_arrays_0_0_ext_ram_wdata3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.650 1792.280 1557.930 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[7]
  PIN data_arrays_0_0_ext_ram_wdata3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.870 1792.280 1561.150 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[8]
  PIN data_arrays_0_0_ext_ram_wdata3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.090 1792.280 1564.370 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata3[9]
  PIN data_arrays_0_0_ext_ram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 838.480 4.000 839.080 ;
    END
  END data_arrays_0_0_ext_ram_web0
  PIN data_arrays_0_0_ext_ram_web1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1734.040 4.000 1734.640 ;
    END
  END data_arrays_0_0_ext_ram_web1
  PIN data_arrays_0_0_ext_ram_web2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 1792.280 556.970 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_web2
  PIN data_arrays_0_0_ext_ram_web3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.310 1792.280 1751.590 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_web3
  PIN data_arrays_0_0_ext_ram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.800 4.000 821.400 ;
    END
  END data_arrays_0_0_ext_ram_wmask0[0]
  PIN data_arrays_0_0_ext_ram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.920 4.000 827.520 ;
    END
  END data_arrays_0_0_ext_ram_wmask0[1]
  PIN data_arrays_0_0_ext_ram_wmask1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.680 4.000 1716.280 ;
    END
  END data_arrays_0_0_ext_ram_wmask1[0]
  PIN data_arrays_0_0_ext_ram_wmask1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1721.800 4.000 1722.400 ;
    END
  END data_arrays_0_0_ext_ram_wmask1[1]
  PIN data_arrays_0_0_ext_ram_wmask2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 1792.280 547.310 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wmask2[0]
  PIN data_arrays_0_0_ext_ram_wmask2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 1792.280 550.530 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wmask2[1]
  PIN data_arrays_0_0_ext_ram_wmask3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.650 1792.280 1741.930 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wmask3[0]
  PIN data_arrays_0_0_ext_ram_wmask3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.870 1792.280 1745.150 1796.280 ;
    END
  END data_arrays_0_0_ext_ram_wmask3[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 19.760 1785.560 20.360 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1217.240 1785.560 1217.840 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1336.920 1785.560 1337.520 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1456.600 1785.560 1457.200 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1576.280 1785.560 1576.880 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1695.960 1785.560 1696.560 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.470 1792.280 1289.750 1796.280 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.810 1792.280 1280.090 1796.280 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1270.150 1792.280 1270.430 1796.280 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.490 1792.280 1260.770 1796.280 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.830 1792.280 1251.110 1796.280 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 139.440 1785.560 140.040 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.170 1792.280 1241.450 1796.280 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.510 1792.280 1231.790 1796.280 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.850 1792.280 1222.130 1796.280 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.190 1792.280 1212.470 1796.280 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.530 1792.280 1202.810 1796.280 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.870 1792.280 1193.150 1796.280 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 1792.280 1183.490 1796.280 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.550 1792.280 1173.830 1796.280 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 1792.280 1164.170 1796.280 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.230 1792.280 1154.510 1796.280 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 259.120 1785.560 259.720 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.570 1792.280 1144.850 1796.280 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 1792.280 1134.730 1796.280 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 1792.280 1125.070 1796.280 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 1792.280 1115.410 1796.280 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.470 1792.280 1105.750 1796.280 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 1792.280 1096.090 1796.280 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 1792.280 1086.430 1796.280 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 1792.280 1076.770 1796.280 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 378.800 1785.560 379.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 498.480 1785.560 499.080 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 618.160 1785.560 618.760 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 737.840 1785.560 738.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 857.520 1785.560 858.120 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 977.880 1785.560 978.480 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1097.560 1785.560 1098.160 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 59.200 1785.560 59.800 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1257.360 1785.560 1257.960 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1377.040 1785.560 1377.640 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1496.720 1785.560 1497.320 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1616.400 1785.560 1617.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1736.080 1785.560 1736.680 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.690 1792.280 1292.970 1796.280 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.030 1792.280 1283.310 1796.280 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.370 1792.280 1273.650 1796.280 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.710 1792.280 1263.990 1796.280 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.050 1792.280 1254.330 1796.280 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 178.880 1785.560 179.480 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.390 1792.280 1244.670 1796.280 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.730 1792.280 1235.010 1796.280 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.070 1792.280 1225.350 1796.280 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.410 1792.280 1215.690 1796.280 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.750 1792.280 1206.030 1796.280 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.090 1792.280 1196.370 1796.280 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.430 1792.280 1186.710 1796.280 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 1792.280 1177.050 1796.280 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.110 1792.280 1167.390 1796.280 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 1792.280 1157.730 1796.280 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 298.560 1785.560 299.160 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 1792.280 1148.070 1796.280 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 1792.280 1138.410 1796.280 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 1792.280 1128.290 1796.280 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.350 1792.280 1118.630 1796.280 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.690 1792.280 1108.970 1796.280 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 1792.280 1099.310 1796.280 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 1792.280 1089.650 1796.280 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 1792.280 1079.990 1796.280 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 418.920 1785.560 419.520 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 538.600 1785.560 539.200 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 658.280 1785.560 658.880 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 777.960 1785.560 778.560 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 897.640 1785.560 898.240 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1017.320 1785.560 1017.920 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1137.000 1785.560 1137.600 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 99.320 1785.560 99.920 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1296.800 1785.560 1297.400 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1416.480 1785.560 1417.080 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1536.840 1785.560 1537.440 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1656.520 1785.560 1657.120 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1776.200 1785.560 1776.800 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.910 1792.280 1296.190 1796.280 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.250 1792.280 1286.530 1796.280 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.590 1792.280 1276.870 1796.280 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 1792.280 1267.210 1796.280 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 1792.280 1257.550 1796.280 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 219.000 1785.560 219.600 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 1792.280 1247.890 1796.280 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.950 1792.280 1238.230 1796.280 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.290 1792.280 1228.570 1796.280 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.630 1792.280 1218.910 1796.280 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 1792.280 1209.250 1796.280 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.310 1792.280 1199.590 1796.280 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.650 1792.280 1189.930 1796.280 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.990 1792.280 1180.270 1796.280 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.330 1792.280 1170.610 1796.280 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 1792.280 1160.950 1796.280 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 338.680 1785.560 339.280 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.010 1792.280 1151.290 1796.280 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 1792.280 1141.630 1796.280 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.230 1792.280 1131.510 1796.280 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.570 1792.280 1121.850 1796.280 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 1792.280 1112.190 1796.280 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 1792.280 1102.530 1796.280 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 1792.280 1092.870 1796.280 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 1792.280 1083.210 1796.280 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 458.360 1785.560 458.960 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 578.040 1785.560 578.640 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 698.400 1785.560 699.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 818.080 1785.560 818.680 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 937.760 1785.560 938.360 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1057.440 1785.560 1058.040 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1781.560 1177.120 1785.560 1177.720 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.150 0.000 1776.430 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.830 0.000 1780.110 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.510 0.000 1783.790 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.670 0.000 1482.950 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.710 0.000 1493.990 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.290 0.000 1504.570 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.330 0.000 1515.610 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 0.000 1526.650 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.950 0.000 1537.230 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.990 0.000 1548.270 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 0.000 1558.850 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.610 0.000 1569.890 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 0.000 1580.930 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.230 0.000 1591.510 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.270 0.000 1602.550 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.310 0.000 1613.590 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.890 0.000 1624.170 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.930 0.000 1635.210 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 0.000 1645.790 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.550 0.000 1656.830 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 0.000 1667.870 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.170 0.000 1678.450 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.210 0.000 1689.490 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 0.000 1700.530 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.830 0.000 1711.110 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.870 0.000 1722.150 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 0.000 1732.730 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.490 0.000 1743.770 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.530 0.000 1754.810 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.110 0.000 1765.390 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 0.000 624.590 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 0.000 722.110 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 0.000 765.810 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 0.000 798.470 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 0.000 809.050 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.430 0.000 841.710 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 0.000 852.750 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 0.000 874.370 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 0.000 885.410 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 0.000 907.030 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.370 0.000 928.650 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 0.000 939.690 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.450 0.000 950.730 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 0.000 961.310 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 0.000 993.970 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.310 0.000 1015.590 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 0.000 1026.630 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 0.000 1048.250 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 0.000 1059.290 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 0.000 1080.910 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 0.000 1091.950 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 0.000 1113.570 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 0.000 1124.610 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 0.000 1135.190 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 0.000 1146.230 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.530 0.000 1156.810 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.570 0.000 1167.850 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.190 0.000 1189.470 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.230 0.000 1200.510 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.850 0.000 1222.130 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.890 0.000 1233.170 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.470 0.000 1243.750 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.510 0.000 1254.790 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.130 0.000 1276.410 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.170 0.000 1287.450 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.790 0.000 1309.070 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.830 0.000 1320.110 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 0.000 1330.690 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.450 0.000 1341.730 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.070 0.000 1363.350 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.110 0.000 1374.390 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 0.000 1384.970 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.730 0.000 1396.010 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.770 0.000 1407.050 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 0.000 1417.630 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.390 0.000 1428.670 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.010 0.000 1450.290 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.050 0.000 1461.330 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 0.000 1475.590 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.350 0.000 1486.630 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 0.000 1497.670 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.970 0.000 1508.250 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.010 0.000 1519.290 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 0.000 1529.870 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.630 0.000 1540.910 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.670 0.000 1551.950 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.250 0.000 1562.530 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.290 0.000 1573.570 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 0.000 1584.610 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.910 0.000 1595.190 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.950 0.000 1606.230 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 0.000 1616.810 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.570 0.000 1627.850 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.610 0.000 1638.890 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.190 0.000 1649.470 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.230 0.000 1660.510 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 0.000 1671.550 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.850 0.000 1682.130 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.890 0.000 1693.170 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 0.000 1703.750 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.510 0.000 1714.790 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.550 0.000 1725.830 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.130 0.000 1736.410 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 0.000 1747.450 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.790 0.000 1769.070 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 0.000 725.790 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 0.000 791.110 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 0.000 845.390 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 0.000 856.430 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 0.000 878.050 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 0.000 921.750 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 0.000 943.370 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 0.000 953.950 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 0.000 964.990 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 0.000 986.610 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.370 0.000 997.650 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 0.000 1008.690 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 0.000 1019.270 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.030 0.000 1030.310 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 0.000 1040.890 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 0.000 1051.930 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 0.000 1073.550 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 0.000 1084.590 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 0.000 1095.630 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.930 0.000 1106.210 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.970 0.000 1117.250 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.550 0.000 1127.830 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.590 0.000 1138.870 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.210 0.000 1160.490 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.250 0.000 1171.530 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.290 0.000 1182.570 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.870 0.000 1193.150 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.910 0.000 1204.190 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 0.000 1214.770 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.530 0.000 1225.810 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.190 0.000 1258.470 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.810 0.000 1280.090 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.850 0.000 1291.130 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 0.000 1301.710 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.470 0.000 1312.750 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.090 0.000 1334.370 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.130 0.000 1345.410 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.750 0.000 1367.030 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.790 0.000 1378.070 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.370 0.000 1388.650 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.410 0.000 1399.690 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 0.000 1421.310 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.070 0.000 1432.350 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 0.000 1442.930 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 0.000 1453.970 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.730 0.000 1465.010 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.990 0.000 1479.270 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.030 0.000 1490.310 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 0.000 1500.890 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.650 0.000 1511.930 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.690 0.000 1522.970 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.270 0.000 1533.550 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.310 0.000 1544.590 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 0.000 1555.630 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.930 0.000 1566.210 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.970 0.000 1577.250 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.550 0.000 1587.830 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.590 0.000 1598.870 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.630 0.000 1609.910 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.210 0.000 1620.490 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.250 0.000 1631.530 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 0.000 1642.570 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.870 0.000 1653.150 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.910 0.000 1664.190 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 0.000 1674.770 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.530 0.000 1685.810 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.570 0.000 1696.850 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1707.150 0.000 1707.430 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 0.000 1718.470 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 0.000 1729.510 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.810 0.000 1740.090 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.850 0.000 1751.130 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 0.000 1761.710 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.470 0.000 1772.750 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 0.000 642.530 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 0.000 696.810 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 0.000 740.510 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 0.000 751.090 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 0.000 762.130 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 0.000 794.790 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 0.000 816.410 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 0.000 827.450 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 0.000 838.030 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.070 0.000 903.350 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.110 0.000 914.390 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 0.000 924.970 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 0.000 936.010 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 0.000 957.630 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 0.000 968.670 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 0.000 979.710 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 0.000 990.290 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.050 0.000 1001.330 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.630 0.000 1011.910 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.670 0.000 1022.950 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 0.000 1044.570 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.330 0.000 1055.610 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 0.000 1066.650 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 0.000 1077.230 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.990 0.000 1088.270 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.230 0.000 1131.510 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.270 0.000 1142.550 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.310 0.000 1153.590 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 0.000 1164.170 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.930 0.000 1175.210 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.510 0.000 1185.790 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.550 0.000 1196.830 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.210 0.000 1229.490 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.830 0.000 1251.110 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.870 0.000 1262.150 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 0.000 1272.730 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.490 0.000 1283.770 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.110 0.000 1305.390 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 0.000 1316.430 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.770 0.000 1338.050 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.810 0.000 1349.090 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.390 0.000 1359.670 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 0.000 1370.710 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 0.000 1381.750 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.050 0.000 1392.330 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 0.000 1403.370 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.710 0.000 1424.990 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.750 0.000 1436.030 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 0.000 1446.610 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.370 0.000 1457.650 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END la_oenb[9]
  PIN ram_clk_delay_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 1792.280 1.750 1796.280 ;
    END
  END ram_clk_delay_sel[0]
  PIN ram_clk_delay_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 1792.280 33.950 1796.280 ;
    END
  END ram_clk_delay_sel[10]
  PIN ram_clk_delay_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 1792.280 37.170 1796.280 ;
    END
  END ram_clk_delay_sel[11]
  PIN ram_clk_delay_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 1792.280 40.390 1796.280 ;
    END
  END ram_clk_delay_sel[12]
  PIN ram_clk_delay_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 1792.280 43.610 1796.280 ;
    END
  END ram_clk_delay_sel[13]
  PIN ram_clk_delay_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 1792.280 46.830 1796.280 ;
    END
  END ram_clk_delay_sel[14]
  PIN ram_clk_delay_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 1792.280 50.050 1796.280 ;
    END
  END ram_clk_delay_sel[15]
  PIN ram_clk_delay_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 1792.280 53.270 1796.280 ;
    END
  END ram_clk_delay_sel[16]
  PIN ram_clk_delay_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 1792.280 56.490 1796.280 ;
    END
  END ram_clk_delay_sel[17]
  PIN ram_clk_delay_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 1792.280 59.710 1796.280 ;
    END
  END ram_clk_delay_sel[18]
  PIN ram_clk_delay_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 1792.280 62.930 1796.280 ;
    END
  END ram_clk_delay_sel[19]
  PIN ram_clk_delay_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 1792.280 4.970 1796.280 ;
    END
  END ram_clk_delay_sel[1]
  PIN ram_clk_delay_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 1792.280 66.150 1796.280 ;
    END
  END ram_clk_delay_sel[20]
  PIN ram_clk_delay_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 1792.280 69.370 1796.280 ;
    END
  END ram_clk_delay_sel[21]
  PIN ram_clk_delay_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 1792.280 72.590 1796.280 ;
    END
  END ram_clk_delay_sel[22]
  PIN ram_clk_delay_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 1792.280 75.810 1796.280 ;
    END
  END ram_clk_delay_sel[23]
  PIN ram_clk_delay_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 1792.280 79.030 1796.280 ;
    END
  END ram_clk_delay_sel[24]
  PIN ram_clk_delay_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 1792.280 82.250 1796.280 ;
    END
  END ram_clk_delay_sel[25]
  PIN ram_clk_delay_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 1792.280 85.470 1796.280 ;
    END
  END ram_clk_delay_sel[26]
  PIN ram_clk_delay_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 1792.280 88.690 1796.280 ;
    END
  END ram_clk_delay_sel[27]
  PIN ram_clk_delay_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 1792.280 91.910 1796.280 ;
    END
  END ram_clk_delay_sel[28]
  PIN ram_clk_delay_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 1792.280 95.130 1796.280 ;
    END
  END ram_clk_delay_sel[29]
  PIN ram_clk_delay_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 1792.280 8.190 1796.280 ;
    END
  END ram_clk_delay_sel[2]
  PIN ram_clk_delay_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 1792.280 98.350 1796.280 ;
    END
  END ram_clk_delay_sel[30]
  PIN ram_clk_delay_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 1792.280 101.570 1796.280 ;
    END
  END ram_clk_delay_sel[31]
  PIN ram_clk_delay_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 1792.280 11.410 1796.280 ;
    END
  END ram_clk_delay_sel[3]
  PIN ram_clk_delay_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 1792.280 14.630 1796.280 ;
    END
  END ram_clk_delay_sel[4]
  PIN ram_clk_delay_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 1792.280 17.850 1796.280 ;
    END
  END ram_clk_delay_sel[5]
  PIN ram_clk_delay_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 1792.280 21.070 1796.280 ;
    END
  END ram_clk_delay_sel[6]
  PIN ram_clk_delay_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 1792.280 24.290 1796.280 ;
    END
  END ram_clk_delay_sel[7]
  PIN ram_clk_delay_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 1792.280 27.510 1796.280 ;
    END
  END ram_clk_delay_sel[8]
  PIN ram_clk_delay_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 1792.280 30.730 1796.280 ;
    END
  END ram_clk_delay_sel[9]
  PIN tag_array_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 1792.280 947.510 1796.280 ;
    END
  END tag_array_ext_ram_addr1[0]
  PIN tag_array_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.450 1792.280 950.730 1796.280 ;
    END
  END tag_array_ext_ram_addr1[1]
  PIN tag_array_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 1792.280 953.950 1796.280 ;
    END
  END tag_array_ext_ram_addr1[2]
  PIN tag_array_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.890 1792.280 957.170 1796.280 ;
    END
  END tag_array_ext_ram_addr1[3]
  PIN tag_array_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 1792.280 960.390 1796.280 ;
    END
  END tag_array_ext_ram_addr1[4]
  PIN tag_array_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 1792.280 963.610 1796.280 ;
    END
  END tag_array_ext_ram_addr1[5]
  PIN tag_array_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 1792.280 966.830 1796.280 ;
    END
  END tag_array_ext_ram_addr1[6]
  PIN tag_array_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 1792.280 970.050 1796.280 ;
    END
  END tag_array_ext_ram_addr1[7]
  PIN tag_array_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 1792.280 695.890 1796.280 ;
    END
  END tag_array_ext_ram_addr[0]
  PIN tag_array_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 1792.280 699.110 1796.280 ;
    END
  END tag_array_ext_ram_addr[1]
  PIN tag_array_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 1792.280 702.330 1796.280 ;
    END
  END tag_array_ext_ram_addr[2]
  PIN tag_array_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 1792.280 705.550 1796.280 ;
    END
  END tag_array_ext_ram_addr[3]
  PIN tag_array_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 1792.280 708.770 1796.280 ;
    END
  END tag_array_ext_ram_addr[4]
  PIN tag_array_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 1792.280 711.990 1796.280 ;
    END
  END tag_array_ext_ram_addr[5]
  PIN tag_array_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 1792.280 715.210 1796.280 ;
    END
  END tag_array_ext_ram_addr[6]
  PIN tag_array_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 1792.280 718.430 1796.280 ;
    END
  END tag_array_ext_ram_addr[7]
  PIN tag_array_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1792.280 721.650 1796.280 ;
    END
  END tag_array_ext_ram_clk
  PIN tag_array_ext_ram_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 1792.280 937.850 1796.280 ;
    END
  END tag_array_ext_ram_csb
  PIN tag_array_ext_ram_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 1792.280 944.290 1796.280 ;
    END
  END tag_array_ext_ram_csb1
  PIN tag_array_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 1792.280 592.390 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[0]
  PIN tag_array_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 1792.280 624.590 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[10]
  PIN tag_array_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 1792.280 627.810 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[11]
  PIN tag_array_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 1792.280 631.030 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[12]
  PIN tag_array_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 1792.280 634.250 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[13]
  PIN tag_array_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 1792.280 637.470 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[14]
  PIN tag_array_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 1792.280 640.690 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[15]
  PIN tag_array_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 1792.280 643.910 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[16]
  PIN tag_array_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 1792.280 647.130 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[17]
  PIN tag_array_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 1792.280 650.350 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[18]
  PIN tag_array_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1792.280 654.030 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[19]
  PIN tag_array_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 1792.280 595.610 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[1]
  PIN tag_array_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 1792.280 657.250 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[20]
  PIN tag_array_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 1792.280 660.470 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[21]
  PIN tag_array_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 1792.280 663.690 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[22]
  PIN tag_array_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 1792.280 666.910 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[23]
  PIN tag_array_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 1792.280 670.130 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[24]
  PIN tag_array_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 1792.280 673.350 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[25]
  PIN tag_array_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 1792.280 676.570 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[26]
  PIN tag_array_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 1792.280 679.790 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[27]
  PIN tag_array_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 1792.280 683.010 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[28]
  PIN tag_array_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 1792.280 686.230 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[29]
  PIN tag_array_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 1792.280 598.830 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[2]
  PIN tag_array_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1792.280 689.450 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[30]
  PIN tag_array_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 1792.280 692.670 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[31]
  PIN tag_array_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 1792.280 602.050 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[3]
  PIN tag_array_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 1792.280 605.270 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[4]
  PIN tag_array_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 1792.280 608.490 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[5]
  PIN tag_array_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 1792.280 611.710 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[6]
  PIN tag_array_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 1792.280 614.930 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[7]
  PIN tag_array_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 1792.280 618.150 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[8]
  PIN tag_array_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 1792.280 621.370 1796.280 ;
    END
  END tag_array_ext_ram_rdata0[9]
  PIN tag_array_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.990 1792.280 973.270 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[0]
  PIN tag_array_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.650 1792.280 1005.930 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[10]
  PIN tag_array_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.870 1792.280 1009.150 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[11]
  PIN tag_array_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.090 1792.280 1012.370 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[12]
  PIN tag_array_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.310 1792.280 1015.590 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[13]
  PIN tag_array_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.530 1792.280 1018.810 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[14]
  PIN tag_array_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.750 1792.280 1022.030 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[15]
  PIN tag_array_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 1792.280 1025.250 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[16]
  PIN tag_array_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.190 1792.280 1028.470 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[17]
  PIN tag_array_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.410 1792.280 1031.690 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[18]
  PIN tag_array_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.630 1792.280 1034.910 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[19]
  PIN tag_array_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 1792.280 976.950 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[1]
  PIN tag_array_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 1792.280 1038.130 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[20]
  PIN tag_array_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.070 1792.280 1041.350 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[21]
  PIN tag_array_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 1792.280 1044.570 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[22]
  PIN tag_array_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 1792.280 1047.790 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[23]
  PIN tag_array_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 1792.280 1051.010 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[24]
  PIN tag_array_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 1792.280 1054.230 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[25]
  PIN tag_array_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.170 1792.280 1057.450 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[26]
  PIN tag_array_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.390 1792.280 1060.670 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[27]
  PIN tag_array_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.610 1792.280 1063.890 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[28]
  PIN tag_array_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.830 1792.280 1067.110 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[29]
  PIN tag_array_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 1792.280 980.170 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[2]
  PIN tag_array_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 1792.280 1070.330 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[30]
  PIN tag_array_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 1792.280 1073.550 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[31]
  PIN tag_array_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 1792.280 983.390 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[3]
  PIN tag_array_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 1792.280 986.610 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[4]
  PIN tag_array_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 1792.280 989.830 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[5]
  PIN tag_array_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.770 1792.280 993.050 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[6]
  PIN tag_array_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 1792.280 996.270 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[7]
  PIN tag_array_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 1792.280 999.490 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[8]
  PIN tag_array_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 1792.280 1002.710 1796.280 ;
    END
  END tag_array_ext_ram_rdata1[9]
  PIN tag_array_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 1792.280 724.870 1796.280 ;
    END
  END tag_array_ext_ram_wdata[0]
  PIN tag_array_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 1792.280 757.070 1796.280 ;
    END
  END tag_array_ext_ram_wdata[10]
  PIN tag_array_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 1792.280 760.290 1796.280 ;
    END
  END tag_array_ext_ram_wdata[11]
  PIN tag_array_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1792.280 763.510 1796.280 ;
    END
  END tag_array_ext_ram_wdata[12]
  PIN tag_array_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 1792.280 766.730 1796.280 ;
    END
  END tag_array_ext_ram_wdata[13]
  PIN tag_array_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 1792.280 769.950 1796.280 ;
    END
  END tag_array_ext_ram_wdata[14]
  PIN tag_array_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 1792.280 773.170 1796.280 ;
    END
  END tag_array_ext_ram_wdata[15]
  PIN tag_array_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 1792.280 776.390 1796.280 ;
    END
  END tag_array_ext_ram_wdata[16]
  PIN tag_array_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1792.280 779.610 1796.280 ;
    END
  END tag_array_ext_ram_wdata[17]
  PIN tag_array_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 1792.280 782.830 1796.280 ;
    END
  END tag_array_ext_ram_wdata[18]
  PIN tag_array_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 1792.280 786.050 1796.280 ;
    END
  END tag_array_ext_ram_wdata[19]
  PIN tag_array_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 1792.280 728.090 1796.280 ;
    END
  END tag_array_ext_ram_wdata[1]
  PIN tag_array_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 1792.280 789.270 1796.280 ;
    END
  END tag_array_ext_ram_wdata[20]
  PIN tag_array_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 1792.280 792.490 1796.280 ;
    END
  END tag_array_ext_ram_wdata[21]
  PIN tag_array_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 1792.280 795.710 1796.280 ;
    END
  END tag_array_ext_ram_wdata[22]
  PIN tag_array_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 1792.280 798.930 1796.280 ;
    END
  END tag_array_ext_ram_wdata[23]
  PIN tag_array_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 1792.280 802.150 1796.280 ;
    END
  END tag_array_ext_ram_wdata[24]
  PIN tag_array_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 1792.280 805.370 1796.280 ;
    END
  END tag_array_ext_ram_wdata[25]
  PIN tag_array_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 1792.280 808.590 1796.280 ;
    END
  END tag_array_ext_ram_wdata[26]
  PIN tag_array_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 1792.280 811.810 1796.280 ;
    END
  END tag_array_ext_ram_wdata[27]
  PIN tag_array_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 1792.280 815.490 1796.280 ;
    END
  END tag_array_ext_ram_wdata[28]
  PIN tag_array_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 1792.280 818.710 1796.280 ;
    END
  END tag_array_ext_ram_wdata[29]
  PIN tag_array_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 1792.280 731.310 1796.280 ;
    END
  END tag_array_ext_ram_wdata[2]
  PIN tag_array_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.650 1792.280 821.930 1796.280 ;
    END
  END tag_array_ext_ram_wdata[30]
  PIN tag_array_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 1792.280 825.150 1796.280 ;
    END
  END tag_array_ext_ram_wdata[31]
  PIN tag_array_ext_ram_wdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 1792.280 828.370 1796.280 ;
    END
  END tag_array_ext_ram_wdata[32]
  PIN tag_array_ext_ram_wdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 1792.280 831.590 1796.280 ;
    END
  END tag_array_ext_ram_wdata[33]
  PIN tag_array_ext_ram_wdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 1792.280 834.810 1796.280 ;
    END
  END tag_array_ext_ram_wdata[34]
  PIN tag_array_ext_ram_wdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 1792.280 838.030 1796.280 ;
    END
  END tag_array_ext_ram_wdata[35]
  PIN tag_array_ext_ram_wdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.970 1792.280 841.250 1796.280 ;
    END
  END tag_array_ext_ram_wdata[36]
  PIN tag_array_ext_ram_wdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 1792.280 844.470 1796.280 ;
    END
  END tag_array_ext_ram_wdata[37]
  PIN tag_array_ext_ram_wdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 1792.280 847.690 1796.280 ;
    END
  END tag_array_ext_ram_wdata[38]
  PIN tag_array_ext_ram_wdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 1792.280 850.910 1796.280 ;
    END
  END tag_array_ext_ram_wdata[39]
  PIN tag_array_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 1792.280 734.530 1796.280 ;
    END
  END tag_array_ext_ram_wdata[3]
  PIN tag_array_ext_ram_wdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 1792.280 854.130 1796.280 ;
    END
  END tag_array_ext_ram_wdata[40]
  PIN tag_array_ext_ram_wdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 1792.280 857.350 1796.280 ;
    END
  END tag_array_ext_ram_wdata[41]
  PIN tag_array_ext_ram_wdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 1792.280 860.570 1796.280 ;
    END
  END tag_array_ext_ram_wdata[42]
  PIN tag_array_ext_ram_wdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 1792.280 863.790 1796.280 ;
    END
  END tag_array_ext_ram_wdata[43]
  PIN tag_array_ext_ram_wdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 1792.280 867.010 1796.280 ;
    END
  END tag_array_ext_ram_wdata[44]
  PIN tag_array_ext_ram_wdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 1792.280 870.230 1796.280 ;
    END
  END tag_array_ext_ram_wdata[45]
  PIN tag_array_ext_ram_wdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 1792.280 873.450 1796.280 ;
    END
  END tag_array_ext_ram_wdata[46]
  PIN tag_array_ext_ram_wdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 1792.280 876.670 1796.280 ;
    END
  END tag_array_ext_ram_wdata[47]
  PIN tag_array_ext_ram_wdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 1792.280 879.890 1796.280 ;
    END
  END tag_array_ext_ram_wdata[48]
  PIN tag_array_ext_ram_wdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 1792.280 883.110 1796.280 ;
    END
  END tag_array_ext_ram_wdata[49]
  PIN tag_array_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 1792.280 737.750 1796.280 ;
    END
  END tag_array_ext_ram_wdata[4]
  PIN tag_array_ext_ram_wdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 1792.280 886.330 1796.280 ;
    END
  END tag_array_ext_ram_wdata[50]
  PIN tag_array_ext_ram_wdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 1792.280 889.550 1796.280 ;
    END
  END tag_array_ext_ram_wdata[51]
  PIN tag_array_ext_ram_wdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 1792.280 892.770 1796.280 ;
    END
  END tag_array_ext_ram_wdata[52]
  PIN tag_array_ext_ram_wdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 1792.280 895.990 1796.280 ;
    END
  END tag_array_ext_ram_wdata[53]
  PIN tag_array_ext_ram_wdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 1792.280 899.210 1796.280 ;
    END
  END tag_array_ext_ram_wdata[54]
  PIN tag_array_ext_ram_wdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.150 1792.280 902.430 1796.280 ;
    END
  END tag_array_ext_ram_wdata[55]
  PIN tag_array_ext_ram_wdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 1792.280 905.650 1796.280 ;
    END
  END tag_array_ext_ram_wdata[56]
  PIN tag_array_ext_ram_wdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 1792.280 908.870 1796.280 ;
    END
  END tag_array_ext_ram_wdata[57]
  PIN tag_array_ext_ram_wdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 1792.280 912.090 1796.280 ;
    END
  END tag_array_ext_ram_wdata[58]
  PIN tag_array_ext_ram_wdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 1792.280 915.310 1796.280 ;
    END
  END tag_array_ext_ram_wdata[59]
  PIN tag_array_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 1792.280 740.970 1796.280 ;
    END
  END tag_array_ext_ram_wdata[5]
  PIN tag_array_ext_ram_wdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 1792.280 918.530 1796.280 ;
    END
  END tag_array_ext_ram_wdata[60]
  PIN tag_array_ext_ram_wdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 1792.280 921.750 1796.280 ;
    END
  END tag_array_ext_ram_wdata[61]
  PIN tag_array_ext_ram_wdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 1792.280 924.970 1796.280 ;
    END
  END tag_array_ext_ram_wdata[62]
  PIN tag_array_ext_ram_wdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 1792.280 928.190 1796.280 ;
    END
  END tag_array_ext_ram_wdata[63]
  PIN tag_array_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 1792.280 744.190 1796.280 ;
    END
  END tag_array_ext_ram_wdata[6]
  PIN tag_array_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1792.280 747.410 1796.280 ;
    END
  END tag_array_ext_ram_wdata[7]
  PIN tag_array_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 1792.280 750.630 1796.280 ;
    END
  END tag_array_ext_ram_wdata[8]
  PIN tag_array_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 1792.280 753.850 1796.280 ;
    END
  END tag_array_ext_ram_wdata[9]
  PIN tag_array_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.790 1792.280 941.070 1796.280 ;
    END
  END tag_array_ext_ram_web
  PIN tag_array_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 1792.280 931.410 1796.280 ;
    END
  END tag_array_ext_ram_wmask[0]
  PIN tag_array_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 1792.280 934.630 1796.280 ;
    END
  END tag_array_ext_ram_wmask[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1784.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1784.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1779.740 1784.405 ;
      LAYER met1 ;
        RECT 1.450 2.420 1783.810 1796.180 ;
      LAYER met2 ;
        RECT 0.090 1792.000 1.190 1796.210 ;
        RECT 2.030 1792.000 4.410 1796.210 ;
        RECT 5.250 1792.000 7.630 1796.210 ;
        RECT 8.470 1792.000 10.850 1796.210 ;
        RECT 11.690 1792.000 14.070 1796.210 ;
        RECT 14.910 1792.000 17.290 1796.210 ;
        RECT 18.130 1792.000 20.510 1796.210 ;
        RECT 21.350 1792.000 23.730 1796.210 ;
        RECT 24.570 1792.000 26.950 1796.210 ;
        RECT 27.790 1792.000 30.170 1796.210 ;
        RECT 31.010 1792.000 33.390 1796.210 ;
        RECT 34.230 1792.000 36.610 1796.210 ;
        RECT 37.450 1792.000 39.830 1796.210 ;
        RECT 40.670 1792.000 43.050 1796.210 ;
        RECT 43.890 1792.000 46.270 1796.210 ;
        RECT 47.110 1792.000 49.490 1796.210 ;
        RECT 50.330 1792.000 52.710 1796.210 ;
        RECT 53.550 1792.000 55.930 1796.210 ;
        RECT 56.770 1792.000 59.150 1796.210 ;
        RECT 59.990 1792.000 62.370 1796.210 ;
        RECT 63.210 1792.000 65.590 1796.210 ;
        RECT 66.430 1792.000 68.810 1796.210 ;
        RECT 69.650 1792.000 72.030 1796.210 ;
        RECT 72.870 1792.000 75.250 1796.210 ;
        RECT 76.090 1792.000 78.470 1796.210 ;
        RECT 79.310 1792.000 81.690 1796.210 ;
        RECT 82.530 1792.000 84.910 1796.210 ;
        RECT 85.750 1792.000 88.130 1796.210 ;
        RECT 88.970 1792.000 91.350 1796.210 ;
        RECT 92.190 1792.000 94.570 1796.210 ;
        RECT 95.410 1792.000 97.790 1796.210 ;
        RECT 98.630 1792.000 101.010 1796.210 ;
        RECT 101.850 1792.000 104.230 1796.210 ;
        RECT 105.070 1792.000 107.450 1796.210 ;
        RECT 108.290 1792.000 110.670 1796.210 ;
        RECT 111.510 1792.000 113.890 1796.210 ;
        RECT 114.730 1792.000 117.110 1796.210 ;
        RECT 117.950 1792.000 120.330 1796.210 ;
        RECT 121.170 1792.000 123.550 1796.210 ;
        RECT 124.390 1792.000 126.770 1796.210 ;
        RECT 127.610 1792.000 129.990 1796.210 ;
        RECT 130.830 1792.000 133.210 1796.210 ;
        RECT 134.050 1792.000 136.430 1796.210 ;
        RECT 137.270 1792.000 139.650 1796.210 ;
        RECT 140.490 1792.000 142.870 1796.210 ;
        RECT 143.710 1792.000 146.090 1796.210 ;
        RECT 146.930 1792.000 149.310 1796.210 ;
        RECT 150.150 1792.000 152.530 1796.210 ;
        RECT 153.370 1792.000 155.750 1796.210 ;
        RECT 156.590 1792.000 158.970 1796.210 ;
        RECT 159.810 1792.000 162.190 1796.210 ;
        RECT 163.030 1792.000 165.870 1796.210 ;
        RECT 166.710 1792.000 169.090 1796.210 ;
        RECT 169.930 1792.000 172.310 1796.210 ;
        RECT 173.150 1792.000 175.530 1796.210 ;
        RECT 176.370 1792.000 178.750 1796.210 ;
        RECT 179.590 1792.000 181.970 1796.210 ;
        RECT 182.810 1792.000 185.190 1796.210 ;
        RECT 186.030 1792.000 188.410 1796.210 ;
        RECT 189.250 1792.000 191.630 1796.210 ;
        RECT 192.470 1792.000 194.850 1796.210 ;
        RECT 195.690 1792.000 198.070 1796.210 ;
        RECT 198.910 1792.000 201.290 1796.210 ;
        RECT 202.130 1792.000 204.510 1796.210 ;
        RECT 205.350 1792.000 207.730 1796.210 ;
        RECT 208.570 1792.000 210.950 1796.210 ;
        RECT 211.790 1792.000 214.170 1796.210 ;
        RECT 215.010 1792.000 217.390 1796.210 ;
        RECT 218.230 1792.000 220.610 1796.210 ;
        RECT 221.450 1792.000 223.830 1796.210 ;
        RECT 224.670 1792.000 227.050 1796.210 ;
        RECT 227.890 1792.000 230.270 1796.210 ;
        RECT 231.110 1792.000 233.490 1796.210 ;
        RECT 234.330 1792.000 236.710 1796.210 ;
        RECT 237.550 1792.000 239.930 1796.210 ;
        RECT 240.770 1792.000 243.150 1796.210 ;
        RECT 243.990 1792.000 246.370 1796.210 ;
        RECT 247.210 1792.000 249.590 1796.210 ;
        RECT 250.430 1792.000 252.810 1796.210 ;
        RECT 253.650 1792.000 256.030 1796.210 ;
        RECT 256.870 1792.000 259.250 1796.210 ;
        RECT 260.090 1792.000 262.470 1796.210 ;
        RECT 263.310 1792.000 265.690 1796.210 ;
        RECT 266.530 1792.000 268.910 1796.210 ;
        RECT 269.750 1792.000 272.130 1796.210 ;
        RECT 272.970 1792.000 275.350 1796.210 ;
        RECT 276.190 1792.000 278.570 1796.210 ;
        RECT 279.410 1792.000 281.790 1796.210 ;
        RECT 282.630 1792.000 285.010 1796.210 ;
        RECT 285.850 1792.000 288.230 1796.210 ;
        RECT 289.070 1792.000 291.450 1796.210 ;
        RECT 292.290 1792.000 294.670 1796.210 ;
        RECT 295.510 1792.000 297.890 1796.210 ;
        RECT 298.730 1792.000 301.110 1796.210 ;
        RECT 301.950 1792.000 304.330 1796.210 ;
        RECT 305.170 1792.000 307.550 1796.210 ;
        RECT 308.390 1792.000 310.770 1796.210 ;
        RECT 311.610 1792.000 313.990 1796.210 ;
        RECT 314.830 1792.000 317.210 1796.210 ;
        RECT 318.050 1792.000 320.430 1796.210 ;
        RECT 321.270 1792.000 323.650 1796.210 ;
        RECT 324.490 1792.000 327.330 1796.210 ;
        RECT 328.170 1792.000 330.550 1796.210 ;
        RECT 331.390 1792.000 333.770 1796.210 ;
        RECT 334.610 1792.000 336.990 1796.210 ;
        RECT 337.830 1792.000 340.210 1796.210 ;
        RECT 341.050 1792.000 343.430 1796.210 ;
        RECT 344.270 1792.000 346.650 1796.210 ;
        RECT 347.490 1792.000 349.870 1796.210 ;
        RECT 350.710 1792.000 353.090 1796.210 ;
        RECT 353.930 1792.000 356.310 1796.210 ;
        RECT 357.150 1792.000 359.530 1796.210 ;
        RECT 360.370 1792.000 362.750 1796.210 ;
        RECT 363.590 1792.000 365.970 1796.210 ;
        RECT 366.810 1792.000 369.190 1796.210 ;
        RECT 370.030 1792.000 372.410 1796.210 ;
        RECT 373.250 1792.000 375.630 1796.210 ;
        RECT 376.470 1792.000 378.850 1796.210 ;
        RECT 379.690 1792.000 382.070 1796.210 ;
        RECT 382.910 1792.000 385.290 1796.210 ;
        RECT 386.130 1792.000 388.510 1796.210 ;
        RECT 389.350 1792.000 391.730 1796.210 ;
        RECT 392.570 1792.000 394.950 1796.210 ;
        RECT 395.790 1792.000 398.170 1796.210 ;
        RECT 399.010 1792.000 401.390 1796.210 ;
        RECT 402.230 1792.000 404.610 1796.210 ;
        RECT 405.450 1792.000 407.830 1796.210 ;
        RECT 408.670 1792.000 411.050 1796.210 ;
        RECT 411.890 1792.000 414.270 1796.210 ;
        RECT 415.110 1792.000 417.490 1796.210 ;
        RECT 418.330 1792.000 420.710 1796.210 ;
        RECT 421.550 1792.000 423.930 1796.210 ;
        RECT 424.770 1792.000 427.150 1796.210 ;
        RECT 427.990 1792.000 430.370 1796.210 ;
        RECT 431.210 1792.000 433.590 1796.210 ;
        RECT 434.430 1792.000 436.810 1796.210 ;
        RECT 437.650 1792.000 440.030 1796.210 ;
        RECT 440.870 1792.000 443.250 1796.210 ;
        RECT 444.090 1792.000 446.470 1796.210 ;
        RECT 447.310 1792.000 449.690 1796.210 ;
        RECT 450.530 1792.000 452.910 1796.210 ;
        RECT 453.750 1792.000 456.130 1796.210 ;
        RECT 456.970 1792.000 459.350 1796.210 ;
        RECT 460.190 1792.000 462.570 1796.210 ;
        RECT 463.410 1792.000 465.790 1796.210 ;
        RECT 466.630 1792.000 469.010 1796.210 ;
        RECT 469.850 1792.000 472.230 1796.210 ;
        RECT 473.070 1792.000 475.450 1796.210 ;
        RECT 476.290 1792.000 478.670 1796.210 ;
        RECT 479.510 1792.000 481.890 1796.210 ;
        RECT 482.730 1792.000 485.110 1796.210 ;
        RECT 485.950 1792.000 488.790 1796.210 ;
        RECT 489.630 1792.000 492.010 1796.210 ;
        RECT 492.850 1792.000 495.230 1796.210 ;
        RECT 496.070 1792.000 498.450 1796.210 ;
        RECT 499.290 1792.000 501.670 1796.210 ;
        RECT 502.510 1792.000 504.890 1796.210 ;
        RECT 505.730 1792.000 508.110 1796.210 ;
        RECT 508.950 1792.000 511.330 1796.210 ;
        RECT 512.170 1792.000 514.550 1796.210 ;
        RECT 515.390 1792.000 517.770 1796.210 ;
        RECT 518.610 1792.000 520.990 1796.210 ;
        RECT 521.830 1792.000 524.210 1796.210 ;
        RECT 525.050 1792.000 527.430 1796.210 ;
        RECT 528.270 1792.000 530.650 1796.210 ;
        RECT 531.490 1792.000 533.870 1796.210 ;
        RECT 534.710 1792.000 537.090 1796.210 ;
        RECT 537.930 1792.000 540.310 1796.210 ;
        RECT 541.150 1792.000 543.530 1796.210 ;
        RECT 544.370 1792.000 546.750 1796.210 ;
        RECT 547.590 1792.000 549.970 1796.210 ;
        RECT 550.810 1792.000 553.190 1796.210 ;
        RECT 554.030 1792.000 556.410 1796.210 ;
        RECT 557.250 1792.000 559.630 1796.210 ;
        RECT 560.470 1792.000 562.850 1796.210 ;
        RECT 563.690 1792.000 566.070 1796.210 ;
        RECT 566.910 1792.000 569.290 1796.210 ;
        RECT 570.130 1792.000 572.510 1796.210 ;
        RECT 573.350 1792.000 575.730 1796.210 ;
        RECT 576.570 1792.000 578.950 1796.210 ;
        RECT 579.790 1792.000 582.170 1796.210 ;
        RECT 583.010 1792.000 585.390 1796.210 ;
        RECT 586.230 1792.000 588.610 1796.210 ;
        RECT 589.450 1792.000 591.830 1796.210 ;
        RECT 592.670 1792.000 595.050 1796.210 ;
        RECT 595.890 1792.000 598.270 1796.210 ;
        RECT 599.110 1792.000 601.490 1796.210 ;
        RECT 602.330 1792.000 604.710 1796.210 ;
        RECT 605.550 1792.000 607.930 1796.210 ;
        RECT 608.770 1792.000 611.150 1796.210 ;
        RECT 611.990 1792.000 614.370 1796.210 ;
        RECT 615.210 1792.000 617.590 1796.210 ;
        RECT 618.430 1792.000 620.810 1796.210 ;
        RECT 621.650 1792.000 624.030 1796.210 ;
        RECT 624.870 1792.000 627.250 1796.210 ;
        RECT 628.090 1792.000 630.470 1796.210 ;
        RECT 631.310 1792.000 633.690 1796.210 ;
        RECT 634.530 1792.000 636.910 1796.210 ;
        RECT 637.750 1792.000 640.130 1796.210 ;
        RECT 640.970 1792.000 643.350 1796.210 ;
        RECT 644.190 1792.000 646.570 1796.210 ;
        RECT 647.410 1792.000 649.790 1796.210 ;
        RECT 650.630 1792.000 653.470 1796.210 ;
        RECT 654.310 1792.000 656.690 1796.210 ;
        RECT 657.530 1792.000 659.910 1796.210 ;
        RECT 660.750 1792.000 663.130 1796.210 ;
        RECT 663.970 1792.000 666.350 1796.210 ;
        RECT 667.190 1792.000 669.570 1796.210 ;
        RECT 670.410 1792.000 672.790 1796.210 ;
        RECT 673.630 1792.000 676.010 1796.210 ;
        RECT 676.850 1792.000 679.230 1796.210 ;
        RECT 680.070 1792.000 682.450 1796.210 ;
        RECT 683.290 1792.000 685.670 1796.210 ;
        RECT 686.510 1792.000 688.890 1796.210 ;
        RECT 689.730 1792.000 692.110 1796.210 ;
        RECT 692.950 1792.000 695.330 1796.210 ;
        RECT 696.170 1792.000 698.550 1796.210 ;
        RECT 699.390 1792.000 701.770 1796.210 ;
        RECT 702.610 1792.000 704.990 1796.210 ;
        RECT 705.830 1792.000 708.210 1796.210 ;
        RECT 709.050 1792.000 711.430 1796.210 ;
        RECT 712.270 1792.000 714.650 1796.210 ;
        RECT 715.490 1792.000 717.870 1796.210 ;
        RECT 718.710 1792.000 721.090 1796.210 ;
        RECT 721.930 1792.000 724.310 1796.210 ;
        RECT 725.150 1792.000 727.530 1796.210 ;
        RECT 728.370 1792.000 730.750 1796.210 ;
        RECT 731.590 1792.000 733.970 1796.210 ;
        RECT 734.810 1792.000 737.190 1796.210 ;
        RECT 738.030 1792.000 740.410 1796.210 ;
        RECT 741.250 1792.000 743.630 1796.210 ;
        RECT 744.470 1792.000 746.850 1796.210 ;
        RECT 747.690 1792.000 750.070 1796.210 ;
        RECT 750.910 1792.000 753.290 1796.210 ;
        RECT 754.130 1792.000 756.510 1796.210 ;
        RECT 757.350 1792.000 759.730 1796.210 ;
        RECT 760.570 1792.000 762.950 1796.210 ;
        RECT 763.790 1792.000 766.170 1796.210 ;
        RECT 767.010 1792.000 769.390 1796.210 ;
        RECT 770.230 1792.000 772.610 1796.210 ;
        RECT 773.450 1792.000 775.830 1796.210 ;
        RECT 776.670 1792.000 779.050 1796.210 ;
        RECT 779.890 1792.000 782.270 1796.210 ;
        RECT 783.110 1792.000 785.490 1796.210 ;
        RECT 786.330 1792.000 788.710 1796.210 ;
        RECT 789.550 1792.000 791.930 1796.210 ;
        RECT 792.770 1792.000 795.150 1796.210 ;
        RECT 795.990 1792.000 798.370 1796.210 ;
        RECT 799.210 1792.000 801.590 1796.210 ;
        RECT 802.430 1792.000 804.810 1796.210 ;
        RECT 805.650 1792.000 808.030 1796.210 ;
        RECT 808.870 1792.000 811.250 1796.210 ;
        RECT 812.090 1792.000 814.930 1796.210 ;
        RECT 815.770 1792.000 818.150 1796.210 ;
        RECT 818.990 1792.000 821.370 1796.210 ;
        RECT 822.210 1792.000 824.590 1796.210 ;
        RECT 825.430 1792.000 827.810 1796.210 ;
        RECT 828.650 1792.000 831.030 1796.210 ;
        RECT 831.870 1792.000 834.250 1796.210 ;
        RECT 835.090 1792.000 837.470 1796.210 ;
        RECT 838.310 1792.000 840.690 1796.210 ;
        RECT 841.530 1792.000 843.910 1796.210 ;
        RECT 844.750 1792.000 847.130 1796.210 ;
        RECT 847.970 1792.000 850.350 1796.210 ;
        RECT 851.190 1792.000 853.570 1796.210 ;
        RECT 854.410 1792.000 856.790 1796.210 ;
        RECT 857.630 1792.000 860.010 1796.210 ;
        RECT 860.850 1792.000 863.230 1796.210 ;
        RECT 864.070 1792.000 866.450 1796.210 ;
        RECT 867.290 1792.000 869.670 1796.210 ;
        RECT 870.510 1792.000 872.890 1796.210 ;
        RECT 873.730 1792.000 876.110 1796.210 ;
        RECT 876.950 1792.000 879.330 1796.210 ;
        RECT 880.170 1792.000 882.550 1796.210 ;
        RECT 883.390 1792.000 885.770 1796.210 ;
        RECT 886.610 1792.000 888.990 1796.210 ;
        RECT 889.830 1792.000 892.210 1796.210 ;
        RECT 893.050 1792.000 895.430 1796.210 ;
        RECT 896.270 1792.000 898.650 1796.210 ;
        RECT 899.490 1792.000 901.870 1796.210 ;
        RECT 902.710 1792.000 905.090 1796.210 ;
        RECT 905.930 1792.000 908.310 1796.210 ;
        RECT 909.150 1792.000 911.530 1796.210 ;
        RECT 912.370 1792.000 914.750 1796.210 ;
        RECT 915.590 1792.000 917.970 1796.210 ;
        RECT 918.810 1792.000 921.190 1796.210 ;
        RECT 922.030 1792.000 924.410 1796.210 ;
        RECT 925.250 1792.000 927.630 1796.210 ;
        RECT 928.470 1792.000 930.850 1796.210 ;
        RECT 931.690 1792.000 934.070 1796.210 ;
        RECT 934.910 1792.000 937.290 1796.210 ;
        RECT 938.130 1792.000 940.510 1796.210 ;
        RECT 941.350 1792.000 943.730 1796.210 ;
        RECT 944.570 1792.000 946.950 1796.210 ;
        RECT 947.790 1792.000 950.170 1796.210 ;
        RECT 951.010 1792.000 953.390 1796.210 ;
        RECT 954.230 1792.000 956.610 1796.210 ;
        RECT 957.450 1792.000 959.830 1796.210 ;
        RECT 960.670 1792.000 963.050 1796.210 ;
        RECT 963.890 1792.000 966.270 1796.210 ;
        RECT 967.110 1792.000 969.490 1796.210 ;
        RECT 970.330 1792.000 972.710 1796.210 ;
        RECT 973.550 1792.000 976.390 1796.210 ;
        RECT 977.230 1792.000 979.610 1796.210 ;
        RECT 980.450 1792.000 982.830 1796.210 ;
        RECT 983.670 1792.000 986.050 1796.210 ;
        RECT 986.890 1792.000 989.270 1796.210 ;
        RECT 990.110 1792.000 992.490 1796.210 ;
        RECT 993.330 1792.000 995.710 1796.210 ;
        RECT 996.550 1792.000 998.930 1796.210 ;
        RECT 999.770 1792.000 1002.150 1796.210 ;
        RECT 1002.990 1792.000 1005.370 1796.210 ;
        RECT 1006.210 1792.000 1008.590 1796.210 ;
        RECT 1009.430 1792.000 1011.810 1796.210 ;
        RECT 1012.650 1792.000 1015.030 1796.210 ;
        RECT 1015.870 1792.000 1018.250 1796.210 ;
        RECT 1019.090 1792.000 1021.470 1796.210 ;
        RECT 1022.310 1792.000 1024.690 1796.210 ;
        RECT 1025.530 1792.000 1027.910 1796.210 ;
        RECT 1028.750 1792.000 1031.130 1796.210 ;
        RECT 1031.970 1792.000 1034.350 1796.210 ;
        RECT 1035.190 1792.000 1037.570 1796.210 ;
        RECT 1038.410 1792.000 1040.790 1796.210 ;
        RECT 1041.630 1792.000 1044.010 1796.210 ;
        RECT 1044.850 1792.000 1047.230 1796.210 ;
        RECT 1048.070 1792.000 1050.450 1796.210 ;
        RECT 1051.290 1792.000 1053.670 1796.210 ;
        RECT 1054.510 1792.000 1056.890 1796.210 ;
        RECT 1057.730 1792.000 1060.110 1796.210 ;
        RECT 1060.950 1792.000 1063.330 1796.210 ;
        RECT 1064.170 1792.000 1066.550 1796.210 ;
        RECT 1067.390 1792.000 1069.770 1796.210 ;
        RECT 1070.610 1792.000 1072.990 1796.210 ;
        RECT 1073.830 1792.000 1076.210 1796.210 ;
        RECT 1077.050 1792.000 1079.430 1796.210 ;
        RECT 1080.270 1792.000 1082.650 1796.210 ;
        RECT 1083.490 1792.000 1085.870 1796.210 ;
        RECT 1086.710 1792.000 1089.090 1796.210 ;
        RECT 1089.930 1792.000 1092.310 1796.210 ;
        RECT 1093.150 1792.000 1095.530 1796.210 ;
        RECT 1096.370 1792.000 1098.750 1796.210 ;
        RECT 1099.590 1792.000 1101.970 1796.210 ;
        RECT 1102.810 1792.000 1105.190 1796.210 ;
        RECT 1106.030 1792.000 1108.410 1796.210 ;
        RECT 1109.250 1792.000 1111.630 1796.210 ;
        RECT 1112.470 1792.000 1114.850 1796.210 ;
        RECT 1115.690 1792.000 1118.070 1796.210 ;
        RECT 1118.910 1792.000 1121.290 1796.210 ;
        RECT 1122.130 1792.000 1124.510 1796.210 ;
        RECT 1125.350 1792.000 1127.730 1796.210 ;
        RECT 1128.570 1792.000 1130.950 1796.210 ;
        RECT 1131.790 1792.000 1134.170 1796.210 ;
        RECT 1135.010 1792.000 1137.850 1796.210 ;
        RECT 1138.690 1792.000 1141.070 1796.210 ;
        RECT 1141.910 1792.000 1144.290 1796.210 ;
        RECT 1145.130 1792.000 1147.510 1796.210 ;
        RECT 1148.350 1792.000 1150.730 1796.210 ;
        RECT 1151.570 1792.000 1153.950 1796.210 ;
        RECT 1154.790 1792.000 1157.170 1796.210 ;
        RECT 1158.010 1792.000 1160.390 1796.210 ;
        RECT 1161.230 1792.000 1163.610 1796.210 ;
        RECT 1164.450 1792.000 1166.830 1796.210 ;
        RECT 1167.670 1792.000 1170.050 1796.210 ;
        RECT 1170.890 1792.000 1173.270 1796.210 ;
        RECT 1174.110 1792.000 1176.490 1796.210 ;
        RECT 1177.330 1792.000 1179.710 1796.210 ;
        RECT 1180.550 1792.000 1182.930 1796.210 ;
        RECT 1183.770 1792.000 1186.150 1796.210 ;
        RECT 1186.990 1792.000 1189.370 1796.210 ;
        RECT 1190.210 1792.000 1192.590 1796.210 ;
        RECT 1193.430 1792.000 1195.810 1796.210 ;
        RECT 1196.650 1792.000 1199.030 1796.210 ;
        RECT 1199.870 1792.000 1202.250 1796.210 ;
        RECT 1203.090 1792.000 1205.470 1796.210 ;
        RECT 1206.310 1792.000 1208.690 1796.210 ;
        RECT 1209.530 1792.000 1211.910 1796.210 ;
        RECT 1212.750 1792.000 1215.130 1796.210 ;
        RECT 1215.970 1792.000 1218.350 1796.210 ;
        RECT 1219.190 1792.000 1221.570 1796.210 ;
        RECT 1222.410 1792.000 1224.790 1796.210 ;
        RECT 1225.630 1792.000 1228.010 1796.210 ;
        RECT 1228.850 1792.000 1231.230 1796.210 ;
        RECT 1232.070 1792.000 1234.450 1796.210 ;
        RECT 1235.290 1792.000 1237.670 1796.210 ;
        RECT 1238.510 1792.000 1240.890 1796.210 ;
        RECT 1241.730 1792.000 1244.110 1796.210 ;
        RECT 1244.950 1792.000 1247.330 1796.210 ;
        RECT 1248.170 1792.000 1250.550 1796.210 ;
        RECT 1251.390 1792.000 1253.770 1796.210 ;
        RECT 1254.610 1792.000 1256.990 1796.210 ;
        RECT 1257.830 1792.000 1260.210 1796.210 ;
        RECT 1261.050 1792.000 1263.430 1796.210 ;
        RECT 1264.270 1792.000 1266.650 1796.210 ;
        RECT 1267.490 1792.000 1269.870 1796.210 ;
        RECT 1270.710 1792.000 1273.090 1796.210 ;
        RECT 1273.930 1792.000 1276.310 1796.210 ;
        RECT 1277.150 1792.000 1279.530 1796.210 ;
        RECT 1280.370 1792.000 1282.750 1796.210 ;
        RECT 1283.590 1792.000 1285.970 1796.210 ;
        RECT 1286.810 1792.000 1289.190 1796.210 ;
        RECT 1290.030 1792.000 1292.410 1796.210 ;
        RECT 1293.250 1792.000 1295.630 1796.210 ;
        RECT 1296.470 1792.000 1298.850 1796.210 ;
        RECT 1299.690 1792.000 1302.530 1796.210 ;
        RECT 1303.370 1792.000 1305.750 1796.210 ;
        RECT 1306.590 1792.000 1308.970 1796.210 ;
        RECT 1309.810 1792.000 1312.190 1796.210 ;
        RECT 1313.030 1792.000 1315.410 1796.210 ;
        RECT 1316.250 1792.000 1318.630 1796.210 ;
        RECT 1319.470 1792.000 1321.850 1796.210 ;
        RECT 1322.690 1792.000 1325.070 1796.210 ;
        RECT 1325.910 1792.000 1328.290 1796.210 ;
        RECT 1329.130 1792.000 1331.510 1796.210 ;
        RECT 1332.350 1792.000 1334.730 1796.210 ;
        RECT 1335.570 1792.000 1337.950 1796.210 ;
        RECT 1338.790 1792.000 1341.170 1796.210 ;
        RECT 1342.010 1792.000 1344.390 1796.210 ;
        RECT 1345.230 1792.000 1347.610 1796.210 ;
        RECT 1348.450 1792.000 1350.830 1796.210 ;
        RECT 1351.670 1792.000 1354.050 1796.210 ;
        RECT 1354.890 1792.000 1357.270 1796.210 ;
        RECT 1358.110 1792.000 1360.490 1796.210 ;
        RECT 1361.330 1792.000 1363.710 1796.210 ;
        RECT 1364.550 1792.000 1366.930 1796.210 ;
        RECT 1367.770 1792.000 1370.150 1796.210 ;
        RECT 1370.990 1792.000 1373.370 1796.210 ;
        RECT 1374.210 1792.000 1376.590 1796.210 ;
        RECT 1377.430 1792.000 1379.810 1796.210 ;
        RECT 1380.650 1792.000 1383.030 1796.210 ;
        RECT 1383.870 1792.000 1386.250 1796.210 ;
        RECT 1387.090 1792.000 1389.470 1796.210 ;
        RECT 1390.310 1792.000 1392.690 1796.210 ;
        RECT 1393.530 1792.000 1395.910 1796.210 ;
        RECT 1396.750 1792.000 1399.130 1796.210 ;
        RECT 1399.970 1792.000 1402.350 1796.210 ;
        RECT 1403.190 1792.000 1405.570 1796.210 ;
        RECT 1406.410 1792.000 1408.790 1796.210 ;
        RECT 1409.630 1792.000 1412.010 1796.210 ;
        RECT 1412.850 1792.000 1415.230 1796.210 ;
        RECT 1416.070 1792.000 1418.450 1796.210 ;
        RECT 1419.290 1792.000 1421.670 1796.210 ;
        RECT 1422.510 1792.000 1424.890 1796.210 ;
        RECT 1425.730 1792.000 1428.110 1796.210 ;
        RECT 1428.950 1792.000 1431.330 1796.210 ;
        RECT 1432.170 1792.000 1434.550 1796.210 ;
        RECT 1435.390 1792.000 1437.770 1796.210 ;
        RECT 1438.610 1792.000 1440.990 1796.210 ;
        RECT 1441.830 1792.000 1444.210 1796.210 ;
        RECT 1445.050 1792.000 1447.430 1796.210 ;
        RECT 1448.270 1792.000 1450.650 1796.210 ;
        RECT 1451.490 1792.000 1453.870 1796.210 ;
        RECT 1454.710 1792.000 1457.090 1796.210 ;
        RECT 1457.930 1792.000 1460.310 1796.210 ;
        RECT 1461.150 1792.000 1463.990 1796.210 ;
        RECT 1464.830 1792.000 1467.210 1796.210 ;
        RECT 1468.050 1792.000 1470.430 1796.210 ;
        RECT 1471.270 1792.000 1473.650 1796.210 ;
        RECT 1474.490 1792.000 1476.870 1796.210 ;
        RECT 1477.710 1792.000 1480.090 1796.210 ;
        RECT 1480.930 1792.000 1483.310 1796.210 ;
        RECT 1484.150 1792.000 1486.530 1796.210 ;
        RECT 1487.370 1792.000 1489.750 1796.210 ;
        RECT 1490.590 1792.000 1492.970 1796.210 ;
        RECT 1493.810 1792.000 1496.190 1796.210 ;
        RECT 1497.030 1792.000 1499.410 1796.210 ;
        RECT 1500.250 1792.000 1502.630 1796.210 ;
        RECT 1503.470 1792.000 1505.850 1796.210 ;
        RECT 1506.690 1792.000 1509.070 1796.210 ;
        RECT 1509.910 1792.000 1512.290 1796.210 ;
        RECT 1513.130 1792.000 1515.510 1796.210 ;
        RECT 1516.350 1792.000 1518.730 1796.210 ;
        RECT 1519.570 1792.000 1521.950 1796.210 ;
        RECT 1522.790 1792.000 1525.170 1796.210 ;
        RECT 1526.010 1792.000 1528.390 1796.210 ;
        RECT 1529.230 1792.000 1531.610 1796.210 ;
        RECT 1532.450 1792.000 1534.830 1796.210 ;
        RECT 1535.670 1792.000 1538.050 1796.210 ;
        RECT 1538.890 1792.000 1541.270 1796.210 ;
        RECT 1542.110 1792.000 1544.490 1796.210 ;
        RECT 1545.330 1792.000 1547.710 1796.210 ;
        RECT 1548.550 1792.000 1550.930 1796.210 ;
        RECT 1551.770 1792.000 1554.150 1796.210 ;
        RECT 1554.990 1792.000 1557.370 1796.210 ;
        RECT 1558.210 1792.000 1560.590 1796.210 ;
        RECT 1561.430 1792.000 1563.810 1796.210 ;
        RECT 1564.650 1792.000 1567.030 1796.210 ;
        RECT 1567.870 1792.000 1570.250 1796.210 ;
        RECT 1571.090 1792.000 1573.470 1796.210 ;
        RECT 1574.310 1792.000 1576.690 1796.210 ;
        RECT 1577.530 1792.000 1579.910 1796.210 ;
        RECT 1580.750 1792.000 1583.130 1796.210 ;
        RECT 1583.970 1792.000 1586.350 1796.210 ;
        RECT 1587.190 1792.000 1589.570 1796.210 ;
        RECT 1590.410 1792.000 1592.790 1796.210 ;
        RECT 1593.630 1792.000 1596.010 1796.210 ;
        RECT 1596.850 1792.000 1599.230 1796.210 ;
        RECT 1600.070 1792.000 1602.450 1796.210 ;
        RECT 1603.290 1792.000 1605.670 1796.210 ;
        RECT 1606.510 1792.000 1608.890 1796.210 ;
        RECT 1609.730 1792.000 1612.110 1796.210 ;
        RECT 1612.950 1792.000 1615.330 1796.210 ;
        RECT 1616.170 1792.000 1618.550 1796.210 ;
        RECT 1619.390 1792.000 1621.770 1796.210 ;
        RECT 1622.610 1792.000 1625.450 1796.210 ;
        RECT 1626.290 1792.000 1628.670 1796.210 ;
        RECT 1629.510 1792.000 1631.890 1796.210 ;
        RECT 1632.730 1792.000 1635.110 1796.210 ;
        RECT 1635.950 1792.000 1638.330 1796.210 ;
        RECT 1639.170 1792.000 1641.550 1796.210 ;
        RECT 1642.390 1792.000 1644.770 1796.210 ;
        RECT 1645.610 1792.000 1647.990 1796.210 ;
        RECT 1648.830 1792.000 1651.210 1796.210 ;
        RECT 1652.050 1792.000 1654.430 1796.210 ;
        RECT 1655.270 1792.000 1657.650 1796.210 ;
        RECT 1658.490 1792.000 1660.870 1796.210 ;
        RECT 1661.710 1792.000 1664.090 1796.210 ;
        RECT 1664.930 1792.000 1667.310 1796.210 ;
        RECT 1668.150 1792.000 1670.530 1796.210 ;
        RECT 1671.370 1792.000 1673.750 1796.210 ;
        RECT 1674.590 1792.000 1676.970 1796.210 ;
        RECT 1677.810 1792.000 1680.190 1796.210 ;
        RECT 1681.030 1792.000 1683.410 1796.210 ;
        RECT 1684.250 1792.000 1686.630 1796.210 ;
        RECT 1687.470 1792.000 1689.850 1796.210 ;
        RECT 1690.690 1792.000 1693.070 1796.210 ;
        RECT 1693.910 1792.000 1696.290 1796.210 ;
        RECT 1697.130 1792.000 1699.510 1796.210 ;
        RECT 1700.350 1792.000 1702.730 1796.210 ;
        RECT 1703.570 1792.000 1705.950 1796.210 ;
        RECT 1706.790 1792.000 1709.170 1796.210 ;
        RECT 1710.010 1792.000 1712.390 1796.210 ;
        RECT 1713.230 1792.000 1715.610 1796.210 ;
        RECT 1716.450 1792.000 1718.830 1796.210 ;
        RECT 1719.670 1792.000 1722.050 1796.210 ;
        RECT 1722.890 1792.000 1725.270 1796.210 ;
        RECT 1726.110 1792.000 1728.490 1796.210 ;
        RECT 1729.330 1792.000 1731.710 1796.210 ;
        RECT 1732.550 1792.000 1734.930 1796.210 ;
        RECT 1735.770 1792.000 1738.150 1796.210 ;
        RECT 1738.990 1792.000 1741.370 1796.210 ;
        RECT 1742.210 1792.000 1744.590 1796.210 ;
        RECT 1745.430 1792.000 1747.810 1796.210 ;
        RECT 1748.650 1792.000 1751.030 1796.210 ;
        RECT 1751.870 1792.000 1754.250 1796.210 ;
        RECT 1755.090 1792.000 1757.470 1796.210 ;
        RECT 1758.310 1792.000 1760.690 1796.210 ;
        RECT 1761.530 1792.000 1763.910 1796.210 ;
        RECT 1764.750 1792.000 1767.130 1796.210 ;
        RECT 1767.970 1792.000 1770.350 1796.210 ;
        RECT 1771.190 1792.000 1773.570 1796.210 ;
        RECT 1774.410 1792.000 1776.790 1796.210 ;
        RECT 1777.630 1792.000 1780.010 1796.210 ;
        RECT 1780.850 1792.000 1783.230 1796.210 ;
        RECT 0.090 4.280 1783.780 1792.000 ;
        RECT 0.090 2.390 1.190 4.280 ;
        RECT 2.030 2.390 4.410 4.280 ;
        RECT 5.250 2.390 8.090 4.280 ;
        RECT 8.930 2.390 11.770 4.280 ;
        RECT 12.610 2.390 15.450 4.280 ;
        RECT 16.290 2.390 19.130 4.280 ;
        RECT 19.970 2.390 22.810 4.280 ;
        RECT 23.650 2.390 26.490 4.280 ;
        RECT 27.330 2.390 29.710 4.280 ;
        RECT 30.550 2.390 33.390 4.280 ;
        RECT 34.230 2.390 37.070 4.280 ;
        RECT 37.910 2.390 40.750 4.280 ;
        RECT 41.590 2.390 44.430 4.280 ;
        RECT 45.270 2.390 48.110 4.280 ;
        RECT 48.950 2.390 51.790 4.280 ;
        RECT 52.630 2.390 55.470 4.280 ;
        RECT 56.310 2.390 58.690 4.280 ;
        RECT 59.530 2.390 62.370 4.280 ;
        RECT 63.210 2.390 66.050 4.280 ;
        RECT 66.890 2.390 69.730 4.280 ;
        RECT 70.570 2.390 73.410 4.280 ;
        RECT 74.250 2.390 77.090 4.280 ;
        RECT 77.930 2.390 80.770 4.280 ;
        RECT 81.610 2.390 84.450 4.280 ;
        RECT 85.290 2.390 87.670 4.280 ;
        RECT 88.510 2.390 91.350 4.280 ;
        RECT 92.190 2.390 95.030 4.280 ;
        RECT 95.870 2.390 98.710 4.280 ;
        RECT 99.550 2.390 102.390 4.280 ;
        RECT 103.230 2.390 106.070 4.280 ;
        RECT 106.910 2.390 109.750 4.280 ;
        RECT 110.590 2.390 113.430 4.280 ;
        RECT 114.270 2.390 116.650 4.280 ;
        RECT 117.490 2.390 120.330 4.280 ;
        RECT 121.170 2.390 124.010 4.280 ;
        RECT 124.850 2.390 127.690 4.280 ;
        RECT 128.530 2.390 131.370 4.280 ;
        RECT 132.210 2.390 135.050 4.280 ;
        RECT 135.890 2.390 138.730 4.280 ;
        RECT 139.570 2.390 142.410 4.280 ;
        RECT 143.250 2.390 145.630 4.280 ;
        RECT 146.470 2.390 149.310 4.280 ;
        RECT 150.150 2.390 152.990 4.280 ;
        RECT 153.830 2.390 156.670 4.280 ;
        RECT 157.510 2.390 160.350 4.280 ;
        RECT 161.190 2.390 164.030 4.280 ;
        RECT 164.870 2.390 167.710 4.280 ;
        RECT 168.550 2.390 171.390 4.280 ;
        RECT 172.230 2.390 174.610 4.280 ;
        RECT 175.450 2.390 178.290 4.280 ;
        RECT 179.130 2.390 181.970 4.280 ;
        RECT 182.810 2.390 185.650 4.280 ;
        RECT 186.490 2.390 189.330 4.280 ;
        RECT 190.170 2.390 193.010 4.280 ;
        RECT 193.850 2.390 196.690 4.280 ;
        RECT 197.530 2.390 200.370 4.280 ;
        RECT 201.210 2.390 203.590 4.280 ;
        RECT 204.430 2.390 207.270 4.280 ;
        RECT 208.110 2.390 210.950 4.280 ;
        RECT 211.790 2.390 214.630 4.280 ;
        RECT 215.470 2.390 218.310 4.280 ;
        RECT 219.150 2.390 221.990 4.280 ;
        RECT 222.830 2.390 225.670 4.280 ;
        RECT 226.510 2.390 229.350 4.280 ;
        RECT 230.190 2.390 232.570 4.280 ;
        RECT 233.410 2.390 236.250 4.280 ;
        RECT 237.090 2.390 239.930 4.280 ;
        RECT 240.770 2.390 243.610 4.280 ;
        RECT 244.450 2.390 247.290 4.280 ;
        RECT 248.130 2.390 250.970 4.280 ;
        RECT 251.810 2.390 254.650 4.280 ;
        RECT 255.490 2.390 258.330 4.280 ;
        RECT 259.170 2.390 261.550 4.280 ;
        RECT 262.390 2.390 265.230 4.280 ;
        RECT 266.070 2.390 268.910 4.280 ;
        RECT 269.750 2.390 272.590 4.280 ;
        RECT 273.430 2.390 276.270 4.280 ;
        RECT 277.110 2.390 279.950 4.280 ;
        RECT 280.790 2.390 283.630 4.280 ;
        RECT 284.470 2.390 287.310 4.280 ;
        RECT 288.150 2.390 290.530 4.280 ;
        RECT 291.370 2.390 294.210 4.280 ;
        RECT 295.050 2.390 297.890 4.280 ;
        RECT 298.730 2.390 301.570 4.280 ;
        RECT 302.410 2.390 305.250 4.280 ;
        RECT 306.090 2.390 308.930 4.280 ;
        RECT 309.770 2.390 312.610 4.280 ;
        RECT 313.450 2.390 316.290 4.280 ;
        RECT 317.130 2.390 319.510 4.280 ;
        RECT 320.350 2.390 323.190 4.280 ;
        RECT 324.030 2.390 326.870 4.280 ;
        RECT 327.710 2.390 330.550 4.280 ;
        RECT 331.390 2.390 334.230 4.280 ;
        RECT 335.070 2.390 337.910 4.280 ;
        RECT 338.750 2.390 341.590 4.280 ;
        RECT 342.430 2.390 345.270 4.280 ;
        RECT 346.110 2.390 348.490 4.280 ;
        RECT 349.330 2.390 352.170 4.280 ;
        RECT 353.010 2.390 355.850 4.280 ;
        RECT 356.690 2.390 359.530 4.280 ;
        RECT 360.370 2.390 363.210 4.280 ;
        RECT 364.050 2.390 366.890 4.280 ;
        RECT 367.730 2.390 370.570 4.280 ;
        RECT 371.410 2.390 374.250 4.280 ;
        RECT 375.090 2.390 377.470 4.280 ;
        RECT 378.310 2.390 381.150 4.280 ;
        RECT 381.990 2.390 384.830 4.280 ;
        RECT 385.670 2.390 388.510 4.280 ;
        RECT 389.350 2.390 392.190 4.280 ;
        RECT 393.030 2.390 395.870 4.280 ;
        RECT 396.710 2.390 399.550 4.280 ;
        RECT 400.390 2.390 403.230 4.280 ;
        RECT 404.070 2.390 406.450 4.280 ;
        RECT 407.290 2.390 410.130 4.280 ;
        RECT 410.970 2.390 413.810 4.280 ;
        RECT 414.650 2.390 417.490 4.280 ;
        RECT 418.330 2.390 421.170 4.280 ;
        RECT 422.010 2.390 424.850 4.280 ;
        RECT 425.690 2.390 428.530 4.280 ;
        RECT 429.370 2.390 432.210 4.280 ;
        RECT 433.050 2.390 435.430 4.280 ;
        RECT 436.270 2.390 439.110 4.280 ;
        RECT 439.950 2.390 442.790 4.280 ;
        RECT 443.630 2.390 446.470 4.280 ;
        RECT 447.310 2.390 450.150 4.280 ;
        RECT 450.990 2.390 453.830 4.280 ;
        RECT 454.670 2.390 457.510 4.280 ;
        RECT 458.350 2.390 461.190 4.280 ;
        RECT 462.030 2.390 464.410 4.280 ;
        RECT 465.250 2.390 468.090 4.280 ;
        RECT 468.930 2.390 471.770 4.280 ;
        RECT 472.610 2.390 475.450 4.280 ;
        RECT 476.290 2.390 479.130 4.280 ;
        RECT 479.970 2.390 482.810 4.280 ;
        RECT 483.650 2.390 486.490 4.280 ;
        RECT 487.330 2.390 490.170 4.280 ;
        RECT 491.010 2.390 493.390 4.280 ;
        RECT 494.230 2.390 497.070 4.280 ;
        RECT 497.910 2.390 500.750 4.280 ;
        RECT 501.590 2.390 504.430 4.280 ;
        RECT 505.270 2.390 508.110 4.280 ;
        RECT 508.950 2.390 511.790 4.280 ;
        RECT 512.630 2.390 515.470 4.280 ;
        RECT 516.310 2.390 519.150 4.280 ;
        RECT 519.990 2.390 522.370 4.280 ;
        RECT 523.210 2.390 526.050 4.280 ;
        RECT 526.890 2.390 529.730 4.280 ;
        RECT 530.570 2.390 533.410 4.280 ;
        RECT 534.250 2.390 537.090 4.280 ;
        RECT 537.930 2.390 540.770 4.280 ;
        RECT 541.610 2.390 544.450 4.280 ;
        RECT 545.290 2.390 548.130 4.280 ;
        RECT 548.970 2.390 551.350 4.280 ;
        RECT 552.190 2.390 555.030 4.280 ;
        RECT 555.870 2.390 558.710 4.280 ;
        RECT 559.550 2.390 562.390 4.280 ;
        RECT 563.230 2.390 566.070 4.280 ;
        RECT 566.910 2.390 569.750 4.280 ;
        RECT 570.590 2.390 573.430 4.280 ;
        RECT 574.270 2.390 577.110 4.280 ;
        RECT 577.950 2.390 580.330 4.280 ;
        RECT 581.170 2.390 584.010 4.280 ;
        RECT 584.850 2.390 587.690 4.280 ;
        RECT 588.530 2.390 591.370 4.280 ;
        RECT 592.210 2.390 595.050 4.280 ;
        RECT 595.890 2.390 598.730 4.280 ;
        RECT 599.570 2.390 602.410 4.280 ;
        RECT 603.250 2.390 605.630 4.280 ;
        RECT 606.470 2.390 609.310 4.280 ;
        RECT 610.150 2.390 612.990 4.280 ;
        RECT 613.830 2.390 616.670 4.280 ;
        RECT 617.510 2.390 620.350 4.280 ;
        RECT 621.190 2.390 624.030 4.280 ;
        RECT 624.870 2.390 627.710 4.280 ;
        RECT 628.550 2.390 631.390 4.280 ;
        RECT 632.230 2.390 634.610 4.280 ;
        RECT 635.450 2.390 638.290 4.280 ;
        RECT 639.130 2.390 641.970 4.280 ;
        RECT 642.810 2.390 645.650 4.280 ;
        RECT 646.490 2.390 649.330 4.280 ;
        RECT 650.170 2.390 653.010 4.280 ;
        RECT 653.850 2.390 656.690 4.280 ;
        RECT 657.530 2.390 660.370 4.280 ;
        RECT 661.210 2.390 663.590 4.280 ;
        RECT 664.430 2.390 667.270 4.280 ;
        RECT 668.110 2.390 670.950 4.280 ;
        RECT 671.790 2.390 674.630 4.280 ;
        RECT 675.470 2.390 678.310 4.280 ;
        RECT 679.150 2.390 681.990 4.280 ;
        RECT 682.830 2.390 685.670 4.280 ;
        RECT 686.510 2.390 689.350 4.280 ;
        RECT 690.190 2.390 692.570 4.280 ;
        RECT 693.410 2.390 696.250 4.280 ;
        RECT 697.090 2.390 699.930 4.280 ;
        RECT 700.770 2.390 703.610 4.280 ;
        RECT 704.450 2.390 707.290 4.280 ;
        RECT 708.130 2.390 710.970 4.280 ;
        RECT 711.810 2.390 714.650 4.280 ;
        RECT 715.490 2.390 718.330 4.280 ;
        RECT 719.170 2.390 721.550 4.280 ;
        RECT 722.390 2.390 725.230 4.280 ;
        RECT 726.070 2.390 728.910 4.280 ;
        RECT 729.750 2.390 732.590 4.280 ;
        RECT 733.430 2.390 736.270 4.280 ;
        RECT 737.110 2.390 739.950 4.280 ;
        RECT 740.790 2.390 743.630 4.280 ;
        RECT 744.470 2.390 747.310 4.280 ;
        RECT 748.150 2.390 750.530 4.280 ;
        RECT 751.370 2.390 754.210 4.280 ;
        RECT 755.050 2.390 757.890 4.280 ;
        RECT 758.730 2.390 761.570 4.280 ;
        RECT 762.410 2.390 765.250 4.280 ;
        RECT 766.090 2.390 768.930 4.280 ;
        RECT 769.770 2.390 772.610 4.280 ;
        RECT 773.450 2.390 776.290 4.280 ;
        RECT 777.130 2.390 779.510 4.280 ;
        RECT 780.350 2.390 783.190 4.280 ;
        RECT 784.030 2.390 786.870 4.280 ;
        RECT 787.710 2.390 790.550 4.280 ;
        RECT 791.390 2.390 794.230 4.280 ;
        RECT 795.070 2.390 797.910 4.280 ;
        RECT 798.750 2.390 801.590 4.280 ;
        RECT 802.430 2.390 805.270 4.280 ;
        RECT 806.110 2.390 808.490 4.280 ;
        RECT 809.330 2.390 812.170 4.280 ;
        RECT 813.010 2.390 815.850 4.280 ;
        RECT 816.690 2.390 819.530 4.280 ;
        RECT 820.370 2.390 823.210 4.280 ;
        RECT 824.050 2.390 826.890 4.280 ;
        RECT 827.730 2.390 830.570 4.280 ;
        RECT 831.410 2.390 834.250 4.280 ;
        RECT 835.090 2.390 837.470 4.280 ;
        RECT 838.310 2.390 841.150 4.280 ;
        RECT 841.990 2.390 844.830 4.280 ;
        RECT 845.670 2.390 848.510 4.280 ;
        RECT 849.350 2.390 852.190 4.280 ;
        RECT 853.030 2.390 855.870 4.280 ;
        RECT 856.710 2.390 859.550 4.280 ;
        RECT 860.390 2.390 863.230 4.280 ;
        RECT 864.070 2.390 866.450 4.280 ;
        RECT 867.290 2.390 870.130 4.280 ;
        RECT 870.970 2.390 873.810 4.280 ;
        RECT 874.650 2.390 877.490 4.280 ;
        RECT 878.330 2.390 881.170 4.280 ;
        RECT 882.010 2.390 884.850 4.280 ;
        RECT 885.690 2.390 888.530 4.280 ;
        RECT 889.370 2.390 892.210 4.280 ;
        RECT 893.050 2.390 895.430 4.280 ;
        RECT 896.270 2.390 899.110 4.280 ;
        RECT 899.950 2.390 902.790 4.280 ;
        RECT 903.630 2.390 906.470 4.280 ;
        RECT 907.310 2.390 910.150 4.280 ;
        RECT 910.990 2.390 913.830 4.280 ;
        RECT 914.670 2.390 917.510 4.280 ;
        RECT 918.350 2.390 921.190 4.280 ;
        RECT 922.030 2.390 924.410 4.280 ;
        RECT 925.250 2.390 928.090 4.280 ;
        RECT 928.930 2.390 931.770 4.280 ;
        RECT 932.610 2.390 935.450 4.280 ;
        RECT 936.290 2.390 939.130 4.280 ;
        RECT 939.970 2.390 942.810 4.280 ;
        RECT 943.650 2.390 946.490 4.280 ;
        RECT 947.330 2.390 950.170 4.280 ;
        RECT 951.010 2.390 953.390 4.280 ;
        RECT 954.230 2.390 957.070 4.280 ;
        RECT 957.910 2.390 960.750 4.280 ;
        RECT 961.590 2.390 964.430 4.280 ;
        RECT 965.270 2.390 968.110 4.280 ;
        RECT 968.950 2.390 971.790 4.280 ;
        RECT 972.630 2.390 975.470 4.280 ;
        RECT 976.310 2.390 979.150 4.280 ;
        RECT 979.990 2.390 982.370 4.280 ;
        RECT 983.210 2.390 986.050 4.280 ;
        RECT 986.890 2.390 989.730 4.280 ;
        RECT 990.570 2.390 993.410 4.280 ;
        RECT 994.250 2.390 997.090 4.280 ;
        RECT 997.930 2.390 1000.770 4.280 ;
        RECT 1001.610 2.390 1004.450 4.280 ;
        RECT 1005.290 2.390 1008.130 4.280 ;
        RECT 1008.970 2.390 1011.350 4.280 ;
        RECT 1012.190 2.390 1015.030 4.280 ;
        RECT 1015.870 2.390 1018.710 4.280 ;
        RECT 1019.550 2.390 1022.390 4.280 ;
        RECT 1023.230 2.390 1026.070 4.280 ;
        RECT 1026.910 2.390 1029.750 4.280 ;
        RECT 1030.590 2.390 1033.430 4.280 ;
        RECT 1034.270 2.390 1037.110 4.280 ;
        RECT 1037.950 2.390 1040.330 4.280 ;
        RECT 1041.170 2.390 1044.010 4.280 ;
        RECT 1044.850 2.390 1047.690 4.280 ;
        RECT 1048.530 2.390 1051.370 4.280 ;
        RECT 1052.210 2.390 1055.050 4.280 ;
        RECT 1055.890 2.390 1058.730 4.280 ;
        RECT 1059.570 2.390 1062.410 4.280 ;
        RECT 1063.250 2.390 1066.090 4.280 ;
        RECT 1066.930 2.390 1069.310 4.280 ;
        RECT 1070.150 2.390 1072.990 4.280 ;
        RECT 1073.830 2.390 1076.670 4.280 ;
        RECT 1077.510 2.390 1080.350 4.280 ;
        RECT 1081.190 2.390 1084.030 4.280 ;
        RECT 1084.870 2.390 1087.710 4.280 ;
        RECT 1088.550 2.390 1091.390 4.280 ;
        RECT 1092.230 2.390 1095.070 4.280 ;
        RECT 1095.910 2.390 1098.290 4.280 ;
        RECT 1099.130 2.390 1101.970 4.280 ;
        RECT 1102.810 2.390 1105.650 4.280 ;
        RECT 1106.490 2.390 1109.330 4.280 ;
        RECT 1110.170 2.390 1113.010 4.280 ;
        RECT 1113.850 2.390 1116.690 4.280 ;
        RECT 1117.530 2.390 1120.370 4.280 ;
        RECT 1121.210 2.390 1124.050 4.280 ;
        RECT 1124.890 2.390 1127.270 4.280 ;
        RECT 1128.110 2.390 1130.950 4.280 ;
        RECT 1131.790 2.390 1134.630 4.280 ;
        RECT 1135.470 2.390 1138.310 4.280 ;
        RECT 1139.150 2.390 1141.990 4.280 ;
        RECT 1142.830 2.390 1145.670 4.280 ;
        RECT 1146.510 2.390 1149.350 4.280 ;
        RECT 1150.190 2.390 1153.030 4.280 ;
        RECT 1153.870 2.390 1156.250 4.280 ;
        RECT 1157.090 2.390 1159.930 4.280 ;
        RECT 1160.770 2.390 1163.610 4.280 ;
        RECT 1164.450 2.390 1167.290 4.280 ;
        RECT 1168.130 2.390 1170.970 4.280 ;
        RECT 1171.810 2.390 1174.650 4.280 ;
        RECT 1175.490 2.390 1178.330 4.280 ;
        RECT 1179.170 2.390 1182.010 4.280 ;
        RECT 1182.850 2.390 1185.230 4.280 ;
        RECT 1186.070 2.390 1188.910 4.280 ;
        RECT 1189.750 2.390 1192.590 4.280 ;
        RECT 1193.430 2.390 1196.270 4.280 ;
        RECT 1197.110 2.390 1199.950 4.280 ;
        RECT 1200.790 2.390 1203.630 4.280 ;
        RECT 1204.470 2.390 1207.310 4.280 ;
        RECT 1208.150 2.390 1210.530 4.280 ;
        RECT 1211.370 2.390 1214.210 4.280 ;
        RECT 1215.050 2.390 1217.890 4.280 ;
        RECT 1218.730 2.390 1221.570 4.280 ;
        RECT 1222.410 2.390 1225.250 4.280 ;
        RECT 1226.090 2.390 1228.930 4.280 ;
        RECT 1229.770 2.390 1232.610 4.280 ;
        RECT 1233.450 2.390 1236.290 4.280 ;
        RECT 1237.130 2.390 1239.510 4.280 ;
        RECT 1240.350 2.390 1243.190 4.280 ;
        RECT 1244.030 2.390 1246.870 4.280 ;
        RECT 1247.710 2.390 1250.550 4.280 ;
        RECT 1251.390 2.390 1254.230 4.280 ;
        RECT 1255.070 2.390 1257.910 4.280 ;
        RECT 1258.750 2.390 1261.590 4.280 ;
        RECT 1262.430 2.390 1265.270 4.280 ;
        RECT 1266.110 2.390 1268.490 4.280 ;
        RECT 1269.330 2.390 1272.170 4.280 ;
        RECT 1273.010 2.390 1275.850 4.280 ;
        RECT 1276.690 2.390 1279.530 4.280 ;
        RECT 1280.370 2.390 1283.210 4.280 ;
        RECT 1284.050 2.390 1286.890 4.280 ;
        RECT 1287.730 2.390 1290.570 4.280 ;
        RECT 1291.410 2.390 1294.250 4.280 ;
        RECT 1295.090 2.390 1297.470 4.280 ;
        RECT 1298.310 2.390 1301.150 4.280 ;
        RECT 1301.990 2.390 1304.830 4.280 ;
        RECT 1305.670 2.390 1308.510 4.280 ;
        RECT 1309.350 2.390 1312.190 4.280 ;
        RECT 1313.030 2.390 1315.870 4.280 ;
        RECT 1316.710 2.390 1319.550 4.280 ;
        RECT 1320.390 2.390 1323.230 4.280 ;
        RECT 1324.070 2.390 1326.450 4.280 ;
        RECT 1327.290 2.390 1330.130 4.280 ;
        RECT 1330.970 2.390 1333.810 4.280 ;
        RECT 1334.650 2.390 1337.490 4.280 ;
        RECT 1338.330 2.390 1341.170 4.280 ;
        RECT 1342.010 2.390 1344.850 4.280 ;
        RECT 1345.690 2.390 1348.530 4.280 ;
        RECT 1349.370 2.390 1352.210 4.280 ;
        RECT 1353.050 2.390 1355.430 4.280 ;
        RECT 1356.270 2.390 1359.110 4.280 ;
        RECT 1359.950 2.390 1362.790 4.280 ;
        RECT 1363.630 2.390 1366.470 4.280 ;
        RECT 1367.310 2.390 1370.150 4.280 ;
        RECT 1370.990 2.390 1373.830 4.280 ;
        RECT 1374.670 2.390 1377.510 4.280 ;
        RECT 1378.350 2.390 1381.190 4.280 ;
        RECT 1382.030 2.390 1384.410 4.280 ;
        RECT 1385.250 2.390 1388.090 4.280 ;
        RECT 1388.930 2.390 1391.770 4.280 ;
        RECT 1392.610 2.390 1395.450 4.280 ;
        RECT 1396.290 2.390 1399.130 4.280 ;
        RECT 1399.970 2.390 1402.810 4.280 ;
        RECT 1403.650 2.390 1406.490 4.280 ;
        RECT 1407.330 2.390 1410.170 4.280 ;
        RECT 1411.010 2.390 1413.390 4.280 ;
        RECT 1414.230 2.390 1417.070 4.280 ;
        RECT 1417.910 2.390 1420.750 4.280 ;
        RECT 1421.590 2.390 1424.430 4.280 ;
        RECT 1425.270 2.390 1428.110 4.280 ;
        RECT 1428.950 2.390 1431.790 4.280 ;
        RECT 1432.630 2.390 1435.470 4.280 ;
        RECT 1436.310 2.390 1439.150 4.280 ;
        RECT 1439.990 2.390 1442.370 4.280 ;
        RECT 1443.210 2.390 1446.050 4.280 ;
        RECT 1446.890 2.390 1449.730 4.280 ;
        RECT 1450.570 2.390 1453.410 4.280 ;
        RECT 1454.250 2.390 1457.090 4.280 ;
        RECT 1457.930 2.390 1460.770 4.280 ;
        RECT 1461.610 2.390 1464.450 4.280 ;
        RECT 1465.290 2.390 1468.130 4.280 ;
        RECT 1468.970 2.390 1471.350 4.280 ;
        RECT 1472.190 2.390 1475.030 4.280 ;
        RECT 1475.870 2.390 1478.710 4.280 ;
        RECT 1479.550 2.390 1482.390 4.280 ;
        RECT 1483.230 2.390 1486.070 4.280 ;
        RECT 1486.910 2.390 1489.750 4.280 ;
        RECT 1490.590 2.390 1493.430 4.280 ;
        RECT 1494.270 2.390 1497.110 4.280 ;
        RECT 1497.950 2.390 1500.330 4.280 ;
        RECT 1501.170 2.390 1504.010 4.280 ;
        RECT 1504.850 2.390 1507.690 4.280 ;
        RECT 1508.530 2.390 1511.370 4.280 ;
        RECT 1512.210 2.390 1515.050 4.280 ;
        RECT 1515.890 2.390 1518.730 4.280 ;
        RECT 1519.570 2.390 1522.410 4.280 ;
        RECT 1523.250 2.390 1526.090 4.280 ;
        RECT 1526.930 2.390 1529.310 4.280 ;
        RECT 1530.150 2.390 1532.990 4.280 ;
        RECT 1533.830 2.390 1536.670 4.280 ;
        RECT 1537.510 2.390 1540.350 4.280 ;
        RECT 1541.190 2.390 1544.030 4.280 ;
        RECT 1544.870 2.390 1547.710 4.280 ;
        RECT 1548.550 2.390 1551.390 4.280 ;
        RECT 1552.230 2.390 1555.070 4.280 ;
        RECT 1555.910 2.390 1558.290 4.280 ;
        RECT 1559.130 2.390 1561.970 4.280 ;
        RECT 1562.810 2.390 1565.650 4.280 ;
        RECT 1566.490 2.390 1569.330 4.280 ;
        RECT 1570.170 2.390 1573.010 4.280 ;
        RECT 1573.850 2.390 1576.690 4.280 ;
        RECT 1577.530 2.390 1580.370 4.280 ;
        RECT 1581.210 2.390 1584.050 4.280 ;
        RECT 1584.890 2.390 1587.270 4.280 ;
        RECT 1588.110 2.390 1590.950 4.280 ;
        RECT 1591.790 2.390 1594.630 4.280 ;
        RECT 1595.470 2.390 1598.310 4.280 ;
        RECT 1599.150 2.390 1601.990 4.280 ;
        RECT 1602.830 2.390 1605.670 4.280 ;
        RECT 1606.510 2.390 1609.350 4.280 ;
        RECT 1610.190 2.390 1613.030 4.280 ;
        RECT 1613.870 2.390 1616.250 4.280 ;
        RECT 1617.090 2.390 1619.930 4.280 ;
        RECT 1620.770 2.390 1623.610 4.280 ;
        RECT 1624.450 2.390 1627.290 4.280 ;
        RECT 1628.130 2.390 1630.970 4.280 ;
        RECT 1631.810 2.390 1634.650 4.280 ;
        RECT 1635.490 2.390 1638.330 4.280 ;
        RECT 1639.170 2.390 1642.010 4.280 ;
        RECT 1642.850 2.390 1645.230 4.280 ;
        RECT 1646.070 2.390 1648.910 4.280 ;
        RECT 1649.750 2.390 1652.590 4.280 ;
        RECT 1653.430 2.390 1656.270 4.280 ;
        RECT 1657.110 2.390 1659.950 4.280 ;
        RECT 1660.790 2.390 1663.630 4.280 ;
        RECT 1664.470 2.390 1667.310 4.280 ;
        RECT 1668.150 2.390 1670.990 4.280 ;
        RECT 1671.830 2.390 1674.210 4.280 ;
        RECT 1675.050 2.390 1677.890 4.280 ;
        RECT 1678.730 2.390 1681.570 4.280 ;
        RECT 1682.410 2.390 1685.250 4.280 ;
        RECT 1686.090 2.390 1688.930 4.280 ;
        RECT 1689.770 2.390 1692.610 4.280 ;
        RECT 1693.450 2.390 1696.290 4.280 ;
        RECT 1697.130 2.390 1699.970 4.280 ;
        RECT 1700.810 2.390 1703.190 4.280 ;
        RECT 1704.030 2.390 1706.870 4.280 ;
        RECT 1707.710 2.390 1710.550 4.280 ;
        RECT 1711.390 2.390 1714.230 4.280 ;
        RECT 1715.070 2.390 1717.910 4.280 ;
        RECT 1718.750 2.390 1721.590 4.280 ;
        RECT 1722.430 2.390 1725.270 4.280 ;
        RECT 1726.110 2.390 1728.950 4.280 ;
        RECT 1729.790 2.390 1732.170 4.280 ;
        RECT 1733.010 2.390 1735.850 4.280 ;
        RECT 1736.690 2.390 1739.530 4.280 ;
        RECT 1740.370 2.390 1743.210 4.280 ;
        RECT 1744.050 2.390 1746.890 4.280 ;
        RECT 1747.730 2.390 1750.570 4.280 ;
        RECT 1751.410 2.390 1754.250 4.280 ;
        RECT 1755.090 2.390 1757.930 4.280 ;
        RECT 1758.770 2.390 1761.150 4.280 ;
        RECT 1761.990 2.390 1764.830 4.280 ;
        RECT 1765.670 2.390 1768.510 4.280 ;
        RECT 1769.350 2.390 1772.190 4.280 ;
        RECT 1773.030 2.390 1775.870 4.280 ;
        RECT 1776.710 2.390 1779.550 4.280 ;
        RECT 1780.390 2.390 1783.230 4.280 ;
      LAYER met3 ;
        RECT 0.065 1794.200 1781.560 1794.345 ;
        RECT 4.400 1792.800 1781.560 1794.200 ;
        RECT 0.065 1788.080 1781.560 1792.800 ;
        RECT 4.400 1786.680 1781.560 1788.080 ;
        RECT 0.065 1781.960 1781.560 1786.680 ;
        RECT 4.400 1780.560 1781.560 1781.960 ;
        RECT 0.065 1777.200 1781.560 1780.560 ;
        RECT 0.065 1776.520 1781.160 1777.200 ;
        RECT 4.400 1775.800 1781.160 1776.520 ;
        RECT 4.400 1775.120 1781.560 1775.800 ;
        RECT 0.065 1770.400 1781.560 1775.120 ;
        RECT 4.400 1769.000 1781.560 1770.400 ;
        RECT 0.065 1764.280 1781.560 1769.000 ;
        RECT 4.400 1762.880 1781.560 1764.280 ;
        RECT 0.065 1758.160 1781.560 1762.880 ;
        RECT 4.400 1756.760 1781.560 1758.160 ;
        RECT 0.065 1752.720 1781.560 1756.760 ;
        RECT 4.400 1751.320 1781.560 1752.720 ;
        RECT 0.065 1746.600 1781.560 1751.320 ;
        RECT 4.400 1745.200 1781.560 1746.600 ;
        RECT 0.065 1740.480 1781.560 1745.200 ;
        RECT 4.400 1739.080 1781.560 1740.480 ;
        RECT 0.065 1737.080 1781.560 1739.080 ;
        RECT 0.065 1735.680 1781.160 1737.080 ;
        RECT 0.065 1735.040 1781.560 1735.680 ;
        RECT 4.400 1733.640 1781.560 1735.040 ;
        RECT 0.065 1728.920 1781.560 1733.640 ;
        RECT 4.400 1727.520 1781.560 1728.920 ;
        RECT 0.065 1722.800 1781.560 1727.520 ;
        RECT 4.400 1721.400 1781.560 1722.800 ;
        RECT 0.065 1716.680 1781.560 1721.400 ;
        RECT 4.400 1715.280 1781.560 1716.680 ;
        RECT 0.065 1711.240 1781.560 1715.280 ;
        RECT 4.400 1709.840 1781.560 1711.240 ;
        RECT 0.065 1705.120 1781.560 1709.840 ;
        RECT 4.400 1703.720 1781.560 1705.120 ;
        RECT 0.065 1699.000 1781.560 1703.720 ;
        RECT 4.400 1697.600 1781.560 1699.000 ;
        RECT 0.065 1696.960 1781.560 1697.600 ;
        RECT 0.065 1695.560 1781.160 1696.960 ;
        RECT 0.065 1693.560 1781.560 1695.560 ;
        RECT 4.400 1692.160 1781.560 1693.560 ;
        RECT 0.065 1687.440 1781.560 1692.160 ;
        RECT 4.400 1686.040 1781.560 1687.440 ;
        RECT 0.065 1681.320 1781.560 1686.040 ;
        RECT 4.400 1679.920 1781.560 1681.320 ;
        RECT 0.065 1675.200 1781.560 1679.920 ;
        RECT 4.400 1673.800 1781.560 1675.200 ;
        RECT 0.065 1669.760 1781.560 1673.800 ;
        RECT 4.400 1668.360 1781.560 1669.760 ;
        RECT 0.065 1663.640 1781.560 1668.360 ;
        RECT 4.400 1662.240 1781.560 1663.640 ;
        RECT 0.065 1657.520 1781.560 1662.240 ;
        RECT 4.400 1656.120 1781.160 1657.520 ;
        RECT 0.065 1652.080 1781.560 1656.120 ;
        RECT 4.400 1650.680 1781.560 1652.080 ;
        RECT 0.065 1645.960 1781.560 1650.680 ;
        RECT 4.400 1644.560 1781.560 1645.960 ;
        RECT 0.065 1639.840 1781.560 1644.560 ;
        RECT 4.400 1638.440 1781.560 1639.840 ;
        RECT 0.065 1633.720 1781.560 1638.440 ;
        RECT 4.400 1632.320 1781.560 1633.720 ;
        RECT 0.065 1628.280 1781.560 1632.320 ;
        RECT 4.400 1626.880 1781.560 1628.280 ;
        RECT 0.065 1622.160 1781.560 1626.880 ;
        RECT 4.400 1620.760 1781.560 1622.160 ;
        RECT 0.065 1617.400 1781.560 1620.760 ;
        RECT 0.065 1616.040 1781.160 1617.400 ;
        RECT 4.400 1616.000 1781.160 1616.040 ;
        RECT 4.400 1614.640 1781.560 1616.000 ;
        RECT 0.065 1609.920 1781.560 1614.640 ;
        RECT 4.400 1608.520 1781.560 1609.920 ;
        RECT 0.065 1604.480 1781.560 1608.520 ;
        RECT 4.400 1603.080 1781.560 1604.480 ;
        RECT 0.065 1598.360 1781.560 1603.080 ;
        RECT 4.400 1596.960 1781.560 1598.360 ;
        RECT 0.065 1592.240 1781.560 1596.960 ;
        RECT 4.400 1590.840 1781.560 1592.240 ;
        RECT 0.065 1586.800 1781.560 1590.840 ;
        RECT 4.400 1585.400 1781.560 1586.800 ;
        RECT 0.065 1580.680 1781.560 1585.400 ;
        RECT 4.400 1579.280 1781.560 1580.680 ;
        RECT 0.065 1577.280 1781.560 1579.280 ;
        RECT 0.065 1575.880 1781.160 1577.280 ;
        RECT 0.065 1574.560 1781.560 1575.880 ;
        RECT 4.400 1573.160 1781.560 1574.560 ;
        RECT 0.065 1568.440 1781.560 1573.160 ;
        RECT 4.400 1567.040 1781.560 1568.440 ;
        RECT 0.065 1563.000 1781.560 1567.040 ;
        RECT 4.400 1561.600 1781.560 1563.000 ;
        RECT 0.065 1556.880 1781.560 1561.600 ;
        RECT 4.400 1555.480 1781.560 1556.880 ;
        RECT 0.065 1550.760 1781.560 1555.480 ;
        RECT 4.400 1549.360 1781.560 1550.760 ;
        RECT 0.065 1545.320 1781.560 1549.360 ;
        RECT 4.400 1543.920 1781.560 1545.320 ;
        RECT 0.065 1539.200 1781.560 1543.920 ;
        RECT 4.400 1537.840 1781.560 1539.200 ;
        RECT 4.400 1537.800 1781.160 1537.840 ;
        RECT 0.065 1536.440 1781.160 1537.800 ;
        RECT 0.065 1533.080 1781.560 1536.440 ;
        RECT 4.400 1531.680 1781.560 1533.080 ;
        RECT 0.065 1526.960 1781.560 1531.680 ;
        RECT 4.400 1525.560 1781.560 1526.960 ;
        RECT 0.065 1521.520 1781.560 1525.560 ;
        RECT 4.400 1520.120 1781.560 1521.520 ;
        RECT 0.065 1515.400 1781.560 1520.120 ;
        RECT 4.400 1514.000 1781.560 1515.400 ;
        RECT 0.065 1509.280 1781.560 1514.000 ;
        RECT 4.400 1507.880 1781.560 1509.280 ;
        RECT 0.065 1503.840 1781.560 1507.880 ;
        RECT 4.400 1502.440 1781.560 1503.840 ;
        RECT 0.065 1497.720 1781.560 1502.440 ;
        RECT 4.400 1496.320 1781.160 1497.720 ;
        RECT 0.065 1491.600 1781.560 1496.320 ;
        RECT 4.400 1490.200 1781.560 1491.600 ;
        RECT 0.065 1485.480 1781.560 1490.200 ;
        RECT 4.400 1484.080 1781.560 1485.480 ;
        RECT 0.065 1480.040 1781.560 1484.080 ;
        RECT 4.400 1478.640 1781.560 1480.040 ;
        RECT 0.065 1473.920 1781.560 1478.640 ;
        RECT 4.400 1472.520 1781.560 1473.920 ;
        RECT 0.065 1467.800 1781.560 1472.520 ;
        RECT 4.400 1466.400 1781.560 1467.800 ;
        RECT 0.065 1461.680 1781.560 1466.400 ;
        RECT 4.400 1460.280 1781.560 1461.680 ;
        RECT 0.065 1457.600 1781.560 1460.280 ;
        RECT 0.065 1456.240 1781.160 1457.600 ;
        RECT 4.400 1456.200 1781.160 1456.240 ;
        RECT 4.400 1454.840 1781.560 1456.200 ;
        RECT 0.065 1450.120 1781.560 1454.840 ;
        RECT 4.400 1448.720 1781.560 1450.120 ;
        RECT 0.065 1444.000 1781.560 1448.720 ;
        RECT 4.400 1442.600 1781.560 1444.000 ;
        RECT 0.065 1438.560 1781.560 1442.600 ;
        RECT 4.400 1437.160 1781.560 1438.560 ;
        RECT 0.065 1432.440 1781.560 1437.160 ;
        RECT 4.400 1431.040 1781.560 1432.440 ;
        RECT 0.065 1426.320 1781.560 1431.040 ;
        RECT 4.400 1424.920 1781.560 1426.320 ;
        RECT 0.065 1420.200 1781.560 1424.920 ;
        RECT 4.400 1418.800 1781.560 1420.200 ;
        RECT 0.065 1417.480 1781.560 1418.800 ;
        RECT 0.065 1416.080 1781.160 1417.480 ;
        RECT 0.065 1414.760 1781.560 1416.080 ;
        RECT 4.400 1413.360 1781.560 1414.760 ;
        RECT 0.065 1408.640 1781.560 1413.360 ;
        RECT 4.400 1407.240 1781.560 1408.640 ;
        RECT 0.065 1402.520 1781.560 1407.240 ;
        RECT 4.400 1401.120 1781.560 1402.520 ;
        RECT 0.065 1397.080 1781.560 1401.120 ;
        RECT 4.400 1395.680 1781.560 1397.080 ;
        RECT 0.065 1390.960 1781.560 1395.680 ;
        RECT 4.400 1389.560 1781.560 1390.960 ;
        RECT 0.065 1384.840 1781.560 1389.560 ;
        RECT 4.400 1383.440 1781.560 1384.840 ;
        RECT 0.065 1378.720 1781.560 1383.440 ;
        RECT 4.400 1378.040 1781.560 1378.720 ;
        RECT 4.400 1377.320 1781.160 1378.040 ;
        RECT 0.065 1376.640 1781.160 1377.320 ;
        RECT 0.065 1373.280 1781.560 1376.640 ;
        RECT 4.400 1371.880 1781.560 1373.280 ;
        RECT 0.065 1367.160 1781.560 1371.880 ;
        RECT 4.400 1365.760 1781.560 1367.160 ;
        RECT 0.065 1361.040 1781.560 1365.760 ;
        RECT 4.400 1359.640 1781.560 1361.040 ;
        RECT 0.065 1355.600 1781.560 1359.640 ;
        RECT 4.400 1354.200 1781.560 1355.600 ;
        RECT 0.065 1349.480 1781.560 1354.200 ;
        RECT 4.400 1348.080 1781.560 1349.480 ;
        RECT 0.065 1343.360 1781.560 1348.080 ;
        RECT 4.400 1341.960 1781.560 1343.360 ;
        RECT 0.065 1337.920 1781.560 1341.960 ;
        RECT 0.065 1337.240 1781.160 1337.920 ;
        RECT 4.400 1336.520 1781.160 1337.240 ;
        RECT 4.400 1335.840 1781.560 1336.520 ;
        RECT 0.065 1331.800 1781.560 1335.840 ;
        RECT 4.400 1330.400 1781.560 1331.800 ;
        RECT 0.065 1325.680 1781.560 1330.400 ;
        RECT 4.400 1324.280 1781.560 1325.680 ;
        RECT 0.065 1319.560 1781.560 1324.280 ;
        RECT 4.400 1318.160 1781.560 1319.560 ;
        RECT 0.065 1314.120 1781.560 1318.160 ;
        RECT 4.400 1312.720 1781.560 1314.120 ;
        RECT 0.065 1308.000 1781.560 1312.720 ;
        RECT 4.400 1306.600 1781.560 1308.000 ;
        RECT 0.065 1301.880 1781.560 1306.600 ;
        RECT 4.400 1300.480 1781.560 1301.880 ;
        RECT 0.065 1297.800 1781.560 1300.480 ;
        RECT 0.065 1296.400 1781.160 1297.800 ;
        RECT 0.065 1295.760 1781.560 1296.400 ;
        RECT 4.400 1294.360 1781.560 1295.760 ;
        RECT 0.065 1290.320 1781.560 1294.360 ;
        RECT 4.400 1288.920 1781.560 1290.320 ;
        RECT 0.065 1284.200 1781.560 1288.920 ;
        RECT 4.400 1282.800 1781.560 1284.200 ;
        RECT 0.065 1278.080 1781.560 1282.800 ;
        RECT 4.400 1276.680 1781.560 1278.080 ;
        RECT 0.065 1271.960 1781.560 1276.680 ;
        RECT 4.400 1270.560 1781.560 1271.960 ;
        RECT 0.065 1266.520 1781.560 1270.560 ;
        RECT 4.400 1265.120 1781.560 1266.520 ;
        RECT 0.065 1260.400 1781.560 1265.120 ;
        RECT 4.400 1259.000 1781.560 1260.400 ;
        RECT 0.065 1258.360 1781.560 1259.000 ;
        RECT 0.065 1256.960 1781.160 1258.360 ;
        RECT 0.065 1254.280 1781.560 1256.960 ;
        RECT 4.400 1252.880 1781.560 1254.280 ;
        RECT 0.065 1248.840 1781.560 1252.880 ;
        RECT 4.400 1247.440 1781.560 1248.840 ;
        RECT 0.065 1242.720 1781.560 1247.440 ;
        RECT 4.400 1241.320 1781.560 1242.720 ;
        RECT 0.065 1236.600 1781.560 1241.320 ;
        RECT 4.400 1235.200 1781.560 1236.600 ;
        RECT 0.065 1230.480 1781.560 1235.200 ;
        RECT 4.400 1229.080 1781.560 1230.480 ;
        RECT 0.065 1225.040 1781.560 1229.080 ;
        RECT 4.400 1223.640 1781.560 1225.040 ;
        RECT 0.065 1218.920 1781.560 1223.640 ;
        RECT 4.400 1218.240 1781.560 1218.920 ;
        RECT 4.400 1217.520 1781.160 1218.240 ;
        RECT 0.065 1216.840 1781.160 1217.520 ;
        RECT 0.065 1212.800 1781.560 1216.840 ;
        RECT 4.400 1211.400 1781.560 1212.800 ;
        RECT 0.065 1207.360 1781.560 1211.400 ;
        RECT 4.400 1205.960 1781.560 1207.360 ;
        RECT 0.065 1201.240 1781.560 1205.960 ;
        RECT 4.400 1199.840 1781.560 1201.240 ;
        RECT 0.065 1195.120 1781.560 1199.840 ;
        RECT 4.400 1193.720 1781.560 1195.120 ;
        RECT 0.065 1189.000 1781.560 1193.720 ;
        RECT 4.400 1187.600 1781.560 1189.000 ;
        RECT 0.065 1183.560 1781.560 1187.600 ;
        RECT 4.400 1182.160 1781.560 1183.560 ;
        RECT 0.065 1178.120 1781.560 1182.160 ;
        RECT 0.065 1177.440 1781.160 1178.120 ;
        RECT 4.400 1176.720 1781.160 1177.440 ;
        RECT 4.400 1176.040 1781.560 1176.720 ;
        RECT 0.065 1171.320 1781.560 1176.040 ;
        RECT 4.400 1169.920 1781.560 1171.320 ;
        RECT 0.065 1165.880 1781.560 1169.920 ;
        RECT 4.400 1164.480 1781.560 1165.880 ;
        RECT 0.065 1159.760 1781.560 1164.480 ;
        RECT 4.400 1158.360 1781.560 1159.760 ;
        RECT 0.065 1153.640 1781.560 1158.360 ;
        RECT 4.400 1152.240 1781.560 1153.640 ;
        RECT 0.065 1147.520 1781.560 1152.240 ;
        RECT 4.400 1146.120 1781.560 1147.520 ;
        RECT 0.065 1142.080 1781.560 1146.120 ;
        RECT 4.400 1140.680 1781.560 1142.080 ;
        RECT 0.065 1138.000 1781.560 1140.680 ;
        RECT 0.065 1136.600 1781.160 1138.000 ;
        RECT 0.065 1135.960 1781.560 1136.600 ;
        RECT 4.400 1134.560 1781.560 1135.960 ;
        RECT 0.065 1129.840 1781.560 1134.560 ;
        RECT 4.400 1128.440 1781.560 1129.840 ;
        RECT 0.065 1123.720 1781.560 1128.440 ;
        RECT 4.400 1122.320 1781.560 1123.720 ;
        RECT 0.065 1118.280 1781.560 1122.320 ;
        RECT 4.400 1116.880 1781.560 1118.280 ;
        RECT 0.065 1112.160 1781.560 1116.880 ;
        RECT 4.400 1110.760 1781.560 1112.160 ;
        RECT 0.065 1106.040 1781.560 1110.760 ;
        RECT 4.400 1104.640 1781.560 1106.040 ;
        RECT 0.065 1100.600 1781.560 1104.640 ;
        RECT 4.400 1099.200 1781.560 1100.600 ;
        RECT 0.065 1098.560 1781.560 1099.200 ;
        RECT 0.065 1097.160 1781.160 1098.560 ;
        RECT 0.065 1094.480 1781.560 1097.160 ;
        RECT 4.400 1093.080 1781.560 1094.480 ;
        RECT 0.065 1088.360 1781.560 1093.080 ;
        RECT 4.400 1086.960 1781.560 1088.360 ;
        RECT 0.065 1082.240 1781.560 1086.960 ;
        RECT 4.400 1080.840 1781.560 1082.240 ;
        RECT 0.065 1076.800 1781.560 1080.840 ;
        RECT 4.400 1075.400 1781.560 1076.800 ;
        RECT 0.065 1070.680 1781.560 1075.400 ;
        RECT 4.400 1069.280 1781.560 1070.680 ;
        RECT 0.065 1064.560 1781.560 1069.280 ;
        RECT 4.400 1063.160 1781.560 1064.560 ;
        RECT 0.065 1059.120 1781.560 1063.160 ;
        RECT 4.400 1058.440 1781.560 1059.120 ;
        RECT 4.400 1057.720 1781.160 1058.440 ;
        RECT 0.065 1057.040 1781.160 1057.720 ;
        RECT 0.065 1053.000 1781.560 1057.040 ;
        RECT 4.400 1051.600 1781.560 1053.000 ;
        RECT 0.065 1046.880 1781.560 1051.600 ;
        RECT 4.400 1045.480 1781.560 1046.880 ;
        RECT 0.065 1040.760 1781.560 1045.480 ;
        RECT 4.400 1039.360 1781.560 1040.760 ;
        RECT 0.065 1035.320 1781.560 1039.360 ;
        RECT 4.400 1033.920 1781.560 1035.320 ;
        RECT 0.065 1029.200 1781.560 1033.920 ;
        RECT 4.400 1027.800 1781.560 1029.200 ;
        RECT 0.065 1023.080 1781.560 1027.800 ;
        RECT 4.400 1021.680 1781.560 1023.080 ;
        RECT 0.065 1018.320 1781.560 1021.680 ;
        RECT 0.065 1017.640 1781.160 1018.320 ;
        RECT 4.400 1016.920 1781.160 1017.640 ;
        RECT 4.400 1016.240 1781.560 1016.920 ;
        RECT 0.065 1011.520 1781.560 1016.240 ;
        RECT 4.400 1010.120 1781.560 1011.520 ;
        RECT 0.065 1005.400 1781.560 1010.120 ;
        RECT 4.400 1004.000 1781.560 1005.400 ;
        RECT 0.065 999.280 1781.560 1004.000 ;
        RECT 4.400 997.880 1781.560 999.280 ;
        RECT 0.065 993.840 1781.560 997.880 ;
        RECT 4.400 992.440 1781.560 993.840 ;
        RECT 0.065 987.720 1781.560 992.440 ;
        RECT 4.400 986.320 1781.560 987.720 ;
        RECT 0.065 981.600 1781.560 986.320 ;
        RECT 4.400 980.200 1781.560 981.600 ;
        RECT 0.065 978.880 1781.560 980.200 ;
        RECT 0.065 977.480 1781.160 978.880 ;
        RECT 0.065 975.480 1781.560 977.480 ;
        RECT 4.400 974.080 1781.560 975.480 ;
        RECT 0.065 970.040 1781.560 974.080 ;
        RECT 4.400 968.640 1781.560 970.040 ;
        RECT 0.065 963.920 1781.560 968.640 ;
        RECT 4.400 962.520 1781.560 963.920 ;
        RECT 0.065 957.800 1781.560 962.520 ;
        RECT 4.400 956.400 1781.560 957.800 ;
        RECT 0.065 952.360 1781.560 956.400 ;
        RECT 4.400 950.960 1781.560 952.360 ;
        RECT 0.065 946.240 1781.560 950.960 ;
        RECT 4.400 944.840 1781.560 946.240 ;
        RECT 0.065 940.120 1781.560 944.840 ;
        RECT 4.400 938.760 1781.560 940.120 ;
        RECT 4.400 938.720 1781.160 938.760 ;
        RECT 0.065 937.360 1781.160 938.720 ;
        RECT 0.065 934.000 1781.560 937.360 ;
        RECT 4.400 932.600 1781.560 934.000 ;
        RECT 0.065 928.560 1781.560 932.600 ;
        RECT 4.400 927.160 1781.560 928.560 ;
        RECT 0.065 922.440 1781.560 927.160 ;
        RECT 4.400 921.040 1781.560 922.440 ;
        RECT 0.065 916.320 1781.560 921.040 ;
        RECT 4.400 914.920 1781.560 916.320 ;
        RECT 0.065 910.880 1781.560 914.920 ;
        RECT 4.400 909.480 1781.560 910.880 ;
        RECT 0.065 904.760 1781.560 909.480 ;
        RECT 4.400 903.360 1781.560 904.760 ;
        RECT 0.065 898.640 1781.560 903.360 ;
        RECT 4.400 897.240 1781.160 898.640 ;
        RECT 0.065 892.520 1781.560 897.240 ;
        RECT 4.400 891.120 1781.560 892.520 ;
        RECT 0.065 887.080 1781.560 891.120 ;
        RECT 4.400 885.680 1781.560 887.080 ;
        RECT 0.065 880.960 1781.560 885.680 ;
        RECT 4.400 879.560 1781.560 880.960 ;
        RECT 0.065 874.840 1781.560 879.560 ;
        RECT 4.400 873.440 1781.560 874.840 ;
        RECT 0.065 869.400 1781.560 873.440 ;
        RECT 4.400 868.000 1781.560 869.400 ;
        RECT 0.065 863.280 1781.560 868.000 ;
        RECT 4.400 861.880 1781.560 863.280 ;
        RECT 0.065 858.520 1781.560 861.880 ;
        RECT 0.065 857.160 1781.160 858.520 ;
        RECT 4.400 857.120 1781.160 857.160 ;
        RECT 4.400 855.760 1781.560 857.120 ;
        RECT 0.065 851.040 1781.560 855.760 ;
        RECT 4.400 849.640 1781.560 851.040 ;
        RECT 0.065 845.600 1781.560 849.640 ;
        RECT 4.400 844.200 1781.560 845.600 ;
        RECT 0.065 839.480 1781.560 844.200 ;
        RECT 4.400 838.080 1781.560 839.480 ;
        RECT 0.065 833.360 1781.560 838.080 ;
        RECT 4.400 831.960 1781.560 833.360 ;
        RECT 0.065 827.920 1781.560 831.960 ;
        RECT 4.400 826.520 1781.560 827.920 ;
        RECT 0.065 821.800 1781.560 826.520 ;
        RECT 4.400 820.400 1781.560 821.800 ;
        RECT 0.065 819.080 1781.560 820.400 ;
        RECT 0.065 817.680 1781.160 819.080 ;
        RECT 0.065 815.680 1781.560 817.680 ;
        RECT 4.400 814.280 1781.560 815.680 ;
        RECT 0.065 809.560 1781.560 814.280 ;
        RECT 4.400 808.160 1781.560 809.560 ;
        RECT 0.065 804.120 1781.560 808.160 ;
        RECT 4.400 802.720 1781.560 804.120 ;
        RECT 0.065 798.000 1781.560 802.720 ;
        RECT 4.400 796.600 1781.560 798.000 ;
        RECT 0.065 791.880 1781.560 796.600 ;
        RECT 4.400 790.480 1781.560 791.880 ;
        RECT 0.065 785.760 1781.560 790.480 ;
        RECT 4.400 784.360 1781.560 785.760 ;
        RECT 0.065 780.320 1781.560 784.360 ;
        RECT 4.400 778.960 1781.560 780.320 ;
        RECT 4.400 778.920 1781.160 778.960 ;
        RECT 0.065 777.560 1781.160 778.920 ;
        RECT 0.065 774.200 1781.560 777.560 ;
        RECT 4.400 772.800 1781.560 774.200 ;
        RECT 0.065 768.080 1781.560 772.800 ;
        RECT 4.400 766.680 1781.560 768.080 ;
        RECT 0.065 762.640 1781.560 766.680 ;
        RECT 4.400 761.240 1781.560 762.640 ;
        RECT 0.065 756.520 1781.560 761.240 ;
        RECT 4.400 755.120 1781.560 756.520 ;
        RECT 0.065 750.400 1781.560 755.120 ;
        RECT 4.400 749.000 1781.560 750.400 ;
        RECT 0.065 744.280 1781.560 749.000 ;
        RECT 4.400 742.880 1781.560 744.280 ;
        RECT 0.065 738.840 1781.560 742.880 ;
        RECT 4.400 737.440 1781.160 738.840 ;
        RECT 0.065 732.720 1781.560 737.440 ;
        RECT 4.400 731.320 1781.560 732.720 ;
        RECT 0.065 726.600 1781.560 731.320 ;
        RECT 4.400 725.200 1781.560 726.600 ;
        RECT 0.065 721.160 1781.560 725.200 ;
        RECT 4.400 719.760 1781.560 721.160 ;
        RECT 0.065 715.040 1781.560 719.760 ;
        RECT 4.400 713.640 1781.560 715.040 ;
        RECT 0.065 708.920 1781.560 713.640 ;
        RECT 4.400 707.520 1781.560 708.920 ;
        RECT 0.065 702.800 1781.560 707.520 ;
        RECT 4.400 701.400 1781.560 702.800 ;
        RECT 0.065 699.400 1781.560 701.400 ;
        RECT 0.065 698.000 1781.160 699.400 ;
        RECT 0.065 697.360 1781.560 698.000 ;
        RECT 4.400 695.960 1781.560 697.360 ;
        RECT 0.065 691.240 1781.560 695.960 ;
        RECT 4.400 689.840 1781.560 691.240 ;
        RECT 0.065 685.120 1781.560 689.840 ;
        RECT 4.400 683.720 1781.560 685.120 ;
        RECT 0.065 679.680 1781.560 683.720 ;
        RECT 4.400 678.280 1781.560 679.680 ;
        RECT 0.065 673.560 1781.560 678.280 ;
        RECT 4.400 672.160 1781.560 673.560 ;
        RECT 0.065 667.440 1781.560 672.160 ;
        RECT 4.400 666.040 1781.560 667.440 ;
        RECT 0.065 661.320 1781.560 666.040 ;
        RECT 4.400 659.920 1781.560 661.320 ;
        RECT 0.065 659.280 1781.560 659.920 ;
        RECT 0.065 657.880 1781.160 659.280 ;
        RECT 0.065 655.880 1781.560 657.880 ;
        RECT 4.400 654.480 1781.560 655.880 ;
        RECT 0.065 649.760 1781.560 654.480 ;
        RECT 4.400 648.360 1781.560 649.760 ;
        RECT 0.065 643.640 1781.560 648.360 ;
        RECT 4.400 642.240 1781.560 643.640 ;
        RECT 0.065 637.520 1781.560 642.240 ;
        RECT 4.400 636.120 1781.560 637.520 ;
        RECT 0.065 632.080 1781.560 636.120 ;
        RECT 4.400 630.680 1781.560 632.080 ;
        RECT 0.065 625.960 1781.560 630.680 ;
        RECT 4.400 624.560 1781.560 625.960 ;
        RECT 0.065 619.840 1781.560 624.560 ;
        RECT 4.400 619.160 1781.560 619.840 ;
        RECT 4.400 618.440 1781.160 619.160 ;
        RECT 0.065 617.760 1781.160 618.440 ;
        RECT 0.065 614.400 1781.560 617.760 ;
        RECT 4.400 613.000 1781.560 614.400 ;
        RECT 0.065 608.280 1781.560 613.000 ;
        RECT 4.400 606.880 1781.560 608.280 ;
        RECT 0.065 602.160 1781.560 606.880 ;
        RECT 4.400 600.760 1781.560 602.160 ;
        RECT 0.065 596.040 1781.560 600.760 ;
        RECT 4.400 594.640 1781.560 596.040 ;
        RECT 0.065 590.600 1781.560 594.640 ;
        RECT 4.400 589.200 1781.560 590.600 ;
        RECT 0.065 584.480 1781.560 589.200 ;
        RECT 4.400 583.080 1781.560 584.480 ;
        RECT 0.065 579.040 1781.560 583.080 ;
        RECT 0.065 578.360 1781.160 579.040 ;
        RECT 4.400 577.640 1781.160 578.360 ;
        RECT 4.400 576.960 1781.560 577.640 ;
        RECT 0.065 572.920 1781.560 576.960 ;
        RECT 4.400 571.520 1781.560 572.920 ;
        RECT 0.065 566.800 1781.560 571.520 ;
        RECT 4.400 565.400 1781.560 566.800 ;
        RECT 0.065 560.680 1781.560 565.400 ;
        RECT 4.400 559.280 1781.560 560.680 ;
        RECT 0.065 554.560 1781.560 559.280 ;
        RECT 4.400 553.160 1781.560 554.560 ;
        RECT 0.065 549.120 1781.560 553.160 ;
        RECT 4.400 547.720 1781.560 549.120 ;
        RECT 0.065 543.000 1781.560 547.720 ;
        RECT 4.400 541.600 1781.560 543.000 ;
        RECT 0.065 539.600 1781.560 541.600 ;
        RECT 0.065 538.200 1781.160 539.600 ;
        RECT 0.065 536.880 1781.560 538.200 ;
        RECT 4.400 535.480 1781.560 536.880 ;
        RECT 0.065 531.440 1781.560 535.480 ;
        RECT 4.400 530.040 1781.560 531.440 ;
        RECT 0.065 525.320 1781.560 530.040 ;
        RECT 4.400 523.920 1781.560 525.320 ;
        RECT 0.065 519.200 1781.560 523.920 ;
        RECT 4.400 517.800 1781.560 519.200 ;
        RECT 0.065 513.080 1781.560 517.800 ;
        RECT 4.400 511.680 1781.560 513.080 ;
        RECT 0.065 507.640 1781.560 511.680 ;
        RECT 4.400 506.240 1781.560 507.640 ;
        RECT 0.065 501.520 1781.560 506.240 ;
        RECT 4.400 500.120 1781.560 501.520 ;
        RECT 0.065 499.480 1781.560 500.120 ;
        RECT 0.065 498.080 1781.160 499.480 ;
        RECT 0.065 495.400 1781.560 498.080 ;
        RECT 4.400 494.000 1781.560 495.400 ;
        RECT 0.065 489.280 1781.560 494.000 ;
        RECT 4.400 487.880 1781.560 489.280 ;
        RECT 0.065 483.840 1781.560 487.880 ;
        RECT 4.400 482.440 1781.560 483.840 ;
        RECT 0.065 477.720 1781.560 482.440 ;
        RECT 4.400 476.320 1781.560 477.720 ;
        RECT 0.065 471.600 1781.560 476.320 ;
        RECT 4.400 470.200 1781.560 471.600 ;
        RECT 0.065 466.160 1781.560 470.200 ;
        RECT 4.400 464.760 1781.560 466.160 ;
        RECT 0.065 460.040 1781.560 464.760 ;
        RECT 4.400 459.360 1781.560 460.040 ;
        RECT 4.400 458.640 1781.160 459.360 ;
        RECT 0.065 457.960 1781.160 458.640 ;
        RECT 0.065 453.920 1781.560 457.960 ;
        RECT 4.400 452.520 1781.560 453.920 ;
        RECT 0.065 447.800 1781.560 452.520 ;
        RECT 4.400 446.400 1781.560 447.800 ;
        RECT 0.065 442.360 1781.560 446.400 ;
        RECT 4.400 440.960 1781.560 442.360 ;
        RECT 0.065 436.240 1781.560 440.960 ;
        RECT 4.400 434.840 1781.560 436.240 ;
        RECT 0.065 430.120 1781.560 434.840 ;
        RECT 4.400 428.720 1781.560 430.120 ;
        RECT 0.065 424.680 1781.560 428.720 ;
        RECT 4.400 423.280 1781.560 424.680 ;
        RECT 0.065 419.920 1781.560 423.280 ;
        RECT 0.065 418.560 1781.160 419.920 ;
        RECT 4.400 418.520 1781.160 418.560 ;
        RECT 4.400 417.160 1781.560 418.520 ;
        RECT 0.065 412.440 1781.560 417.160 ;
        RECT 4.400 411.040 1781.560 412.440 ;
        RECT 0.065 406.320 1781.560 411.040 ;
        RECT 4.400 404.920 1781.560 406.320 ;
        RECT 0.065 400.880 1781.560 404.920 ;
        RECT 4.400 399.480 1781.560 400.880 ;
        RECT 0.065 394.760 1781.560 399.480 ;
        RECT 4.400 393.360 1781.560 394.760 ;
        RECT 0.065 388.640 1781.560 393.360 ;
        RECT 4.400 387.240 1781.560 388.640 ;
        RECT 0.065 383.200 1781.560 387.240 ;
        RECT 4.400 381.800 1781.560 383.200 ;
        RECT 0.065 379.800 1781.560 381.800 ;
        RECT 0.065 378.400 1781.160 379.800 ;
        RECT 0.065 377.080 1781.560 378.400 ;
        RECT 4.400 375.680 1781.560 377.080 ;
        RECT 0.065 370.960 1781.560 375.680 ;
        RECT 4.400 369.560 1781.560 370.960 ;
        RECT 0.065 364.840 1781.560 369.560 ;
        RECT 4.400 363.440 1781.560 364.840 ;
        RECT 0.065 359.400 1781.560 363.440 ;
        RECT 4.400 358.000 1781.560 359.400 ;
        RECT 0.065 353.280 1781.560 358.000 ;
        RECT 4.400 351.880 1781.560 353.280 ;
        RECT 0.065 347.160 1781.560 351.880 ;
        RECT 4.400 345.760 1781.560 347.160 ;
        RECT 0.065 341.720 1781.560 345.760 ;
        RECT 4.400 340.320 1781.560 341.720 ;
        RECT 0.065 339.680 1781.560 340.320 ;
        RECT 0.065 338.280 1781.160 339.680 ;
        RECT 0.065 335.600 1781.560 338.280 ;
        RECT 4.400 334.200 1781.560 335.600 ;
        RECT 0.065 329.480 1781.560 334.200 ;
        RECT 4.400 328.080 1781.560 329.480 ;
        RECT 0.065 323.360 1781.560 328.080 ;
        RECT 4.400 321.960 1781.560 323.360 ;
        RECT 0.065 317.920 1781.560 321.960 ;
        RECT 4.400 316.520 1781.560 317.920 ;
        RECT 0.065 311.800 1781.560 316.520 ;
        RECT 4.400 310.400 1781.560 311.800 ;
        RECT 0.065 305.680 1781.560 310.400 ;
        RECT 4.400 304.280 1781.560 305.680 ;
        RECT 0.065 299.560 1781.560 304.280 ;
        RECT 4.400 298.160 1781.160 299.560 ;
        RECT 0.065 294.120 1781.560 298.160 ;
        RECT 4.400 292.720 1781.560 294.120 ;
        RECT 0.065 288.000 1781.560 292.720 ;
        RECT 4.400 286.600 1781.560 288.000 ;
        RECT 0.065 281.880 1781.560 286.600 ;
        RECT 4.400 280.480 1781.560 281.880 ;
        RECT 0.065 276.440 1781.560 280.480 ;
        RECT 4.400 275.040 1781.560 276.440 ;
        RECT 0.065 270.320 1781.560 275.040 ;
        RECT 4.400 268.920 1781.560 270.320 ;
        RECT 0.065 264.200 1781.560 268.920 ;
        RECT 4.400 262.800 1781.560 264.200 ;
        RECT 0.065 260.120 1781.560 262.800 ;
        RECT 0.065 258.720 1781.160 260.120 ;
        RECT 0.065 258.080 1781.560 258.720 ;
        RECT 4.400 256.680 1781.560 258.080 ;
        RECT 0.065 252.640 1781.560 256.680 ;
        RECT 4.400 251.240 1781.560 252.640 ;
        RECT 0.065 246.520 1781.560 251.240 ;
        RECT 4.400 245.120 1781.560 246.520 ;
        RECT 0.065 240.400 1781.560 245.120 ;
        RECT 4.400 239.000 1781.560 240.400 ;
        RECT 0.065 234.960 1781.560 239.000 ;
        RECT 4.400 233.560 1781.560 234.960 ;
        RECT 0.065 228.840 1781.560 233.560 ;
        RECT 4.400 227.440 1781.560 228.840 ;
        RECT 0.065 222.720 1781.560 227.440 ;
        RECT 4.400 221.320 1781.560 222.720 ;
        RECT 0.065 220.000 1781.560 221.320 ;
        RECT 0.065 218.600 1781.160 220.000 ;
        RECT 0.065 216.600 1781.560 218.600 ;
        RECT 4.400 215.200 1781.560 216.600 ;
        RECT 0.065 211.160 1781.560 215.200 ;
        RECT 4.400 209.760 1781.560 211.160 ;
        RECT 0.065 205.040 1781.560 209.760 ;
        RECT 4.400 203.640 1781.560 205.040 ;
        RECT 0.065 198.920 1781.560 203.640 ;
        RECT 4.400 197.520 1781.560 198.920 ;
        RECT 0.065 193.480 1781.560 197.520 ;
        RECT 4.400 192.080 1781.560 193.480 ;
        RECT 0.065 187.360 1781.560 192.080 ;
        RECT 4.400 185.960 1781.560 187.360 ;
        RECT 0.065 181.240 1781.560 185.960 ;
        RECT 4.400 179.880 1781.560 181.240 ;
        RECT 4.400 179.840 1781.160 179.880 ;
        RECT 0.065 178.480 1781.160 179.840 ;
        RECT 0.065 175.120 1781.560 178.480 ;
        RECT 4.400 173.720 1781.560 175.120 ;
        RECT 0.065 169.680 1781.560 173.720 ;
        RECT 4.400 168.280 1781.560 169.680 ;
        RECT 0.065 163.560 1781.560 168.280 ;
        RECT 4.400 162.160 1781.560 163.560 ;
        RECT 0.065 157.440 1781.560 162.160 ;
        RECT 4.400 156.040 1781.560 157.440 ;
        RECT 0.065 151.320 1781.560 156.040 ;
        RECT 4.400 149.920 1781.560 151.320 ;
        RECT 0.065 145.880 1781.560 149.920 ;
        RECT 4.400 144.480 1781.560 145.880 ;
        RECT 0.065 140.440 1781.560 144.480 ;
        RECT 0.065 139.760 1781.160 140.440 ;
        RECT 4.400 139.040 1781.160 139.760 ;
        RECT 4.400 138.360 1781.560 139.040 ;
        RECT 0.065 133.640 1781.560 138.360 ;
        RECT 4.400 132.240 1781.560 133.640 ;
        RECT 0.065 128.200 1781.560 132.240 ;
        RECT 4.400 126.800 1781.560 128.200 ;
        RECT 0.065 122.080 1781.560 126.800 ;
        RECT 4.400 120.680 1781.560 122.080 ;
        RECT 0.065 115.960 1781.560 120.680 ;
        RECT 4.400 114.560 1781.560 115.960 ;
        RECT 0.065 109.840 1781.560 114.560 ;
        RECT 4.400 108.440 1781.560 109.840 ;
        RECT 0.065 104.400 1781.560 108.440 ;
        RECT 4.400 103.000 1781.560 104.400 ;
        RECT 0.065 100.320 1781.560 103.000 ;
        RECT 0.065 98.920 1781.160 100.320 ;
        RECT 0.065 98.280 1781.560 98.920 ;
        RECT 4.400 96.880 1781.560 98.280 ;
        RECT 0.065 92.160 1781.560 96.880 ;
        RECT 4.400 90.760 1781.560 92.160 ;
        RECT 0.065 86.720 1781.560 90.760 ;
        RECT 4.400 85.320 1781.560 86.720 ;
        RECT 0.065 80.600 1781.560 85.320 ;
        RECT 4.400 79.200 1781.560 80.600 ;
        RECT 0.065 74.480 1781.560 79.200 ;
        RECT 4.400 73.080 1781.560 74.480 ;
        RECT 0.065 68.360 1781.560 73.080 ;
        RECT 4.400 66.960 1781.560 68.360 ;
        RECT 0.065 62.920 1781.560 66.960 ;
        RECT 4.400 61.520 1781.560 62.920 ;
        RECT 0.065 60.200 1781.560 61.520 ;
        RECT 0.065 58.800 1781.160 60.200 ;
        RECT 0.065 56.800 1781.560 58.800 ;
        RECT 4.400 55.400 1781.560 56.800 ;
        RECT 0.065 50.680 1781.560 55.400 ;
        RECT 4.400 49.280 1781.560 50.680 ;
        RECT 0.065 45.240 1781.560 49.280 ;
        RECT 4.400 43.840 1781.560 45.240 ;
        RECT 0.065 39.120 1781.560 43.840 ;
        RECT 4.400 37.720 1781.560 39.120 ;
        RECT 0.065 33.000 1781.560 37.720 ;
        RECT 4.400 31.600 1781.560 33.000 ;
        RECT 0.065 26.880 1781.560 31.600 ;
        RECT 4.400 25.480 1781.560 26.880 ;
        RECT 0.065 21.440 1781.560 25.480 ;
        RECT 4.400 20.760 1781.560 21.440 ;
        RECT 4.400 20.040 1781.160 20.760 ;
        RECT 0.065 19.360 1781.160 20.040 ;
        RECT 0.065 15.320 1781.560 19.360 ;
        RECT 4.400 13.920 1781.560 15.320 ;
        RECT 0.065 9.200 1781.560 13.920 ;
        RECT 4.400 7.800 1781.560 9.200 ;
        RECT 0.065 3.760 1781.560 7.800 ;
        RECT 4.400 2.895 1781.560 3.760 ;
      LAYER met4 ;
        RECT 2.135 1784.960 1686.065 1786.185 ;
        RECT 2.135 10.240 20.640 1784.960 ;
        RECT 23.040 10.240 97.440 1784.960 ;
        RECT 99.840 10.240 174.240 1784.960 ;
        RECT 176.640 10.240 251.040 1784.960 ;
        RECT 253.440 10.240 327.840 1784.960 ;
        RECT 330.240 10.240 404.640 1784.960 ;
        RECT 407.040 10.240 481.440 1784.960 ;
        RECT 483.840 10.240 558.240 1784.960 ;
        RECT 560.640 10.240 635.040 1784.960 ;
        RECT 637.440 10.240 711.840 1784.960 ;
        RECT 714.240 10.240 788.640 1784.960 ;
        RECT 791.040 10.240 865.440 1784.960 ;
        RECT 867.840 10.240 942.240 1784.960 ;
        RECT 944.640 10.240 1019.040 1784.960 ;
        RECT 1021.440 10.240 1095.840 1784.960 ;
        RECT 1098.240 10.240 1172.640 1784.960 ;
        RECT 1175.040 10.240 1249.440 1784.960 ;
        RECT 1251.840 10.240 1326.240 1784.960 ;
        RECT 1328.640 10.240 1403.040 1784.960 ;
        RECT 1405.440 10.240 1479.840 1784.960 ;
        RECT 1482.240 10.240 1556.640 1784.960 ;
        RECT 1559.040 10.240 1633.440 1784.960 ;
        RECT 1635.840 10.240 1686.065 1784.960 ;
        RECT 2.135 9.015 1686.065 10.240 ;
  END
END Marmot
END LIBRARY

