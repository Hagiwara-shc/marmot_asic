VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Marmot
  CLASS BLOCK ;
  FOREIGN Marmot ;
  ORIGIN 0.000 0.000 ;
  SIZE 1756.380 BY 1767.100 ;
  PIN data_arrays_0_0_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END data_arrays_0_0_ext_ram_addr1[0]
  PIN data_arrays_0_0_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END data_arrays_0_0_ext_ram_addr1[1]
  PIN data_arrays_0_0_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.280 4.000 947.880 ;
    END
  END data_arrays_0_0_ext_ram_addr1[2]
  PIN data_arrays_0_0_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 953.400 4.000 954.000 ;
    END
  END data_arrays_0_0_ext_ram_addr1[3]
  PIN data_arrays_0_0_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 959.520 4.000 960.120 ;
    END
  END data_arrays_0_0_ext_ram_addr1[4]
  PIN data_arrays_0_0_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END data_arrays_0_0_ext_ram_addr1[5]
  PIN data_arrays_0_0_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END data_arrays_0_0_ext_ram_addr1[6]
  PIN data_arrays_0_0_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.200 4.000 977.800 ;
    END
  END data_arrays_0_0_ext_ram_addr1[7]
  PIN data_arrays_0_0_ext_ram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END data_arrays_0_0_ext_ram_addr1[8]
  PIN data_arrays_0_0_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END data_arrays_0_0_ext_ram_addr[0]
  PIN data_arrays_0_0_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END data_arrays_0_0_ext_ram_addr[1]
  PIN data_arrays_0_0_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END data_arrays_0_0_ext_ram_addr[2]
  PIN data_arrays_0_0_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END data_arrays_0_0_ext_ram_addr[3]
  PIN data_arrays_0_0_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 4.000 417.480 ;
    END
  END data_arrays_0_0_ext_ram_addr[4]
  PIN data_arrays_0_0_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END data_arrays_0_0_ext_ram_addr[5]
  PIN data_arrays_0_0_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END data_arrays_0_0_ext_ram_addr[6]
  PIN data_arrays_0_0_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END data_arrays_0_0_ext_ram_addr[7]
  PIN data_arrays_0_0_ext_ram_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END data_arrays_0_0_ext_ram_addr[8]
  PIN data_arrays_0_0_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END data_arrays_0_0_ext_ram_clk
  PIN data_arrays_0_0_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END data_arrays_0_0_ext_ram_csb1[0]
  PIN data_arrays_0_0_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END data_arrays_0_0_ext_ram_csb1[1]
  PIN data_arrays_0_0_ext_ram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 898.320 4.000 898.920 ;
    END
  END data_arrays_0_0_ext_ram_csb1[2]
  PIN data_arrays_0_0_ext_ram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END data_arrays_0_0_ext_ram_csb1[3]
  PIN data_arrays_0_0_ext_ram_csb1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 910.560 4.000 911.160 ;
    END
  END data_arrays_0_0_ext_ram_csb1[4]
  PIN data_arrays_0_0_ext_ram_csb1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END data_arrays_0_0_ext_ram_csb1[5]
  PIN data_arrays_0_0_ext_ram_csb1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.800 4.000 923.400 ;
    END
  END data_arrays_0_0_ext_ram_csb1[6]
  PIN data_arrays_0_0_ext_ram_csb1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.920 4.000 929.520 ;
    END
  END data_arrays_0_0_ext_ram_csb1[7]
  PIN data_arrays_0_0_ext_ram_csb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END data_arrays_0_0_ext_ram_csb[0]
  PIN data_arrays_0_0_ext_ram_csb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 861.600 4.000 862.200 ;
    END
  END data_arrays_0_0_ext_ram_csb[1]
  PIN data_arrays_0_0_ext_ram_csb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 4.000 868.320 ;
    END
  END data_arrays_0_0_ext_ram_csb[2]
  PIN data_arrays_0_0_ext_ram_csb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END data_arrays_0_0_ext_ram_csb[3]
  PIN data_arrays_0_0_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[0]
  PIN data_arrays_0_0_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[10]
  PIN data_arrays_0_0_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[11]
  PIN data_arrays_0_0_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[12]
  PIN data_arrays_0_0_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[13]
  PIN data_arrays_0_0_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[14]
  PIN data_arrays_0_0_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[15]
  PIN data_arrays_0_0_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[16]
  PIN data_arrays_0_0_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[17]
  PIN data_arrays_0_0_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[18]
  PIN data_arrays_0_0_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[19]
  PIN data_arrays_0_0_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[1]
  PIN data_arrays_0_0_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[20]
  PIN data_arrays_0_0_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[21]
  PIN data_arrays_0_0_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[22]
  PIN data_arrays_0_0_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[23]
  PIN data_arrays_0_0_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[24]
  PIN data_arrays_0_0_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[25]
  PIN data_arrays_0_0_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[26]
  PIN data_arrays_0_0_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[27]
  PIN data_arrays_0_0_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[28]
  PIN data_arrays_0_0_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[29]
  PIN data_arrays_0_0_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[2]
  PIN data_arrays_0_0_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[30]
  PIN data_arrays_0_0_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[31]
  PIN data_arrays_0_0_ext_ram_rdata0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[32]
  PIN data_arrays_0_0_ext_ram_rdata0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[33]
  PIN data_arrays_0_0_ext_ram_rdata0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[34]
  PIN data_arrays_0_0_ext_ram_rdata0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[35]
  PIN data_arrays_0_0_ext_ram_rdata0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[36]
  PIN data_arrays_0_0_ext_ram_rdata0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[37]
  PIN data_arrays_0_0_ext_ram_rdata0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[38]
  PIN data_arrays_0_0_ext_ram_rdata0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[39]
  PIN data_arrays_0_0_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[3]
  PIN data_arrays_0_0_ext_ram_rdata0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[40]
  PIN data_arrays_0_0_ext_ram_rdata0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[41]
  PIN data_arrays_0_0_ext_ram_rdata0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[42]
  PIN data_arrays_0_0_ext_ram_rdata0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[43]
  PIN data_arrays_0_0_ext_ram_rdata0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[44]
  PIN data_arrays_0_0_ext_ram_rdata0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[45]
  PIN data_arrays_0_0_ext_ram_rdata0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[46]
  PIN data_arrays_0_0_ext_ram_rdata0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[47]
  PIN data_arrays_0_0_ext_ram_rdata0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[48]
  PIN data_arrays_0_0_ext_ram_rdata0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[49]
  PIN data_arrays_0_0_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[4]
  PIN data_arrays_0_0_ext_ram_rdata0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[50]
  PIN data_arrays_0_0_ext_ram_rdata0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[51]
  PIN data_arrays_0_0_ext_ram_rdata0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[52]
  PIN data_arrays_0_0_ext_ram_rdata0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[53]
  PIN data_arrays_0_0_ext_ram_rdata0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[54]
  PIN data_arrays_0_0_ext_ram_rdata0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[55]
  PIN data_arrays_0_0_ext_ram_rdata0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[56]
  PIN data_arrays_0_0_ext_ram_rdata0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[57]
  PIN data_arrays_0_0_ext_ram_rdata0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[58]
  PIN data_arrays_0_0_ext_ram_rdata0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[59]
  PIN data_arrays_0_0_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[5]
  PIN data_arrays_0_0_ext_ram_rdata0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[60]
  PIN data_arrays_0_0_ext_ram_rdata0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[61]
  PIN data_arrays_0_0_ext_ram_rdata0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[62]
  PIN data_arrays_0_0_ext_ram_rdata0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[63]
  PIN data_arrays_0_0_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[6]
  PIN data_arrays_0_0_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[7]
  PIN data_arrays_0_0_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[8]
  PIN data_arrays_0_0_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[9]
  PIN data_arrays_0_0_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[0]
  PIN data_arrays_0_0_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[10]
  PIN data_arrays_0_0_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.760 4.000 1057.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[11]
  PIN data_arrays_0_0_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.880 4.000 1063.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[12]
  PIN data_arrays_0_0_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1069.000 4.000 1069.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[13]
  PIN data_arrays_0_0_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.120 4.000 1075.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[14]
  PIN data_arrays_0_0_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[15]
  PIN data_arrays_0_0_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1087.360 4.000 1087.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[16]
  PIN data_arrays_0_0_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1093.480 4.000 1094.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[17]
  PIN data_arrays_0_0_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[18]
  PIN data_arrays_0_0_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.720 4.000 1106.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[19]
  PIN data_arrays_0_0_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 995.560 4.000 996.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[1]
  PIN data_arrays_0_0_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[20]
  PIN data_arrays_0_0_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.960 4.000 1118.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[21]
  PIN data_arrays_0_0_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.080 4.000 1124.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[22]
  PIN data_arrays_0_0_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1129.520 4.000 1130.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[23]
  PIN data_arrays_0_0_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[24]
  PIN data_arrays_0_0_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.760 4.000 1142.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[25]
  PIN data_arrays_0_0_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.880 4.000 1148.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[26]
  PIN data_arrays_0_0_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.000 4.000 1154.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[27]
  PIN data_arrays_0_0_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1160.120 4.000 1160.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[28]
  PIN data_arrays_0_0_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[29]
  PIN data_arrays_0_0_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.680 4.000 1002.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[2]
  PIN data_arrays_0_0_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1172.360 4.000 1172.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[30]
  PIN data_arrays_0_0_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1178.480 4.000 1179.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[31]
  PIN data_arrays_0_0_ext_ram_rdata1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1184.600 4.000 1185.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[32]
  PIN data_arrays_0_0_ext_ram_rdata1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.720 4.000 1191.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[33]
  PIN data_arrays_0_0_ext_ram_rdata1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1196.840 4.000 1197.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[34]
  PIN data_arrays_0_0_ext_ram_rdata1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.960 4.000 1203.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[35]
  PIN data_arrays_0_0_ext_ram_rdata1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1209.080 4.000 1209.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[36]
  PIN data_arrays_0_0_ext_ram_rdata1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1215.200 4.000 1215.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[37]
  PIN data_arrays_0_0_ext_ram_rdata1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1221.320 4.000 1221.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[38]
  PIN data_arrays_0_0_ext_ram_rdata1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[39]
  PIN data_arrays_0_0_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[3]
  PIN data_arrays_0_0_ext_ram_rdata1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1233.560 4.000 1234.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[40]
  PIN data_arrays_0_0_ext_ram_rdata1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.680 4.000 1240.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[41]
  PIN data_arrays_0_0_ext_ram_rdata1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1245.800 4.000 1246.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[42]
  PIN data_arrays_0_0_ext_ram_rdata1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.920 4.000 1252.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[43]
  PIN data_arrays_0_0_ext_ram_rdata1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[44]
  PIN data_arrays_0_0_ext_ram_rdata1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.160 4.000 1264.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[45]
  PIN data_arrays_0_0_ext_ram_rdata1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.280 4.000 1270.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[46]
  PIN data_arrays_0_0_ext_ram_rdata1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1276.400 4.000 1277.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[47]
  PIN data_arrays_0_0_ext_ram_rdata1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1282.520 4.000 1283.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[48]
  PIN data_arrays_0_0_ext_ram_rdata1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1287.960 4.000 1288.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[49]
  PIN data_arrays_0_0_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.920 4.000 1014.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[4]
  PIN data_arrays_0_0_ext_ram_rdata1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1294.080 4.000 1294.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[50]
  PIN data_arrays_0_0_ext_ram_rdata1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.200 4.000 1300.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[51]
  PIN data_arrays_0_0_ext_ram_rdata1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1306.320 4.000 1306.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[52]
  PIN data_arrays_0_0_ext_ram_rdata1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1312.440 4.000 1313.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[53]
  PIN data_arrays_0_0_ext_ram_rdata1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1318.560 4.000 1319.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[54]
  PIN data_arrays_0_0_ext_ram_rdata1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1324.680 4.000 1325.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[55]
  PIN data_arrays_0_0_ext_ram_rdata1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1330.800 4.000 1331.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[56]
  PIN data_arrays_0_0_ext_ram_rdata1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1336.920 4.000 1337.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[57]
  PIN data_arrays_0_0_ext_ram_rdata1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[58]
  PIN data_arrays_0_0_ext_ram_rdata1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.160 4.000 1349.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[59]
  PIN data_arrays_0_0_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[5]
  PIN data_arrays_0_0_ext_ram_rdata1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1355.280 4.000 1355.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[60]
  PIN data_arrays_0_0_ext_ram_rdata1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1361.400 4.000 1362.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[61]
  PIN data_arrays_0_0_ext_ram_rdata1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1367.520 4.000 1368.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[62]
  PIN data_arrays_0_0_ext_ram_rdata1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[63]
  PIN data_arrays_0_0_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.160 4.000 1026.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[6]
  PIN data_arrays_0_0_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.280 4.000 1032.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[7]
  PIN data_arrays_0_0_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1038.400 4.000 1039.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[8]
  PIN data_arrays_0_0_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1044.520 4.000 1045.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[9]
  PIN data_arrays_0_0_ext_ram_rdata2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1379.760 4.000 1380.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[0]
  PIN data_arrays_0_0_ext_ram_rdata2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1440.960 4.000 1441.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[10]
  PIN data_arrays_0_0_ext_ram_rdata2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1447.080 4.000 1447.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[11]
  PIN data_arrays_0_0_ext_ram_rdata2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1452.520 4.000 1453.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[12]
  PIN data_arrays_0_0_ext_ram_rdata2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[13]
  PIN data_arrays_0_0_ext_ram_rdata2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1464.760 4.000 1465.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[14]
  PIN data_arrays_0_0_ext_ram_rdata2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1470.880 4.000 1471.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[15]
  PIN data_arrays_0_0_ext_ram_rdata2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1477.000 4.000 1477.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[16]
  PIN data_arrays_0_0_ext_ram_rdata2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1483.120 4.000 1483.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[17]
  PIN data_arrays_0_0_ext_ram_rdata2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[18]
  PIN data_arrays_0_0_ext_ram_rdata2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1495.360 4.000 1495.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[19]
  PIN data_arrays_0_0_ext_ram_rdata2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1385.880 4.000 1386.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[1]
  PIN data_arrays_0_0_ext_ram_rdata2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1501.480 4.000 1502.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[20]
  PIN data_arrays_0_0_ext_ram_rdata2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1507.600 4.000 1508.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[21]
  PIN data_arrays_0_0_ext_ram_rdata2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1513.720 4.000 1514.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[22]
  PIN data_arrays_0_0_ext_ram_rdata2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1519.840 4.000 1520.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[23]
  PIN data_arrays_0_0_ext_ram_rdata2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1525.960 4.000 1526.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[24]
  PIN data_arrays_0_0_ext_ram_rdata2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1532.080 4.000 1532.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[25]
  PIN data_arrays_0_0_ext_ram_rdata2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1538.200 4.000 1538.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[26]
  PIN data_arrays_0_0_ext_ram_rdata2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1544.320 4.000 1544.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[27]
  PIN data_arrays_0_0_ext_ram_rdata2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[28]
  PIN data_arrays_0_0_ext_ram_rdata2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1556.560 4.000 1557.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[29]
  PIN data_arrays_0_0_ext_ram_rdata2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.000 4.000 1392.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[2]
  PIN data_arrays_0_0_ext_ram_rdata2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1562.680 4.000 1563.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[30]
  PIN data_arrays_0_0_ext_ram_rdata2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1568.800 4.000 1569.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[31]
  PIN data_arrays_0_0_ext_ram_rdata2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.920 4.000 1575.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[32]
  PIN data_arrays_0_0_ext_ram_rdata2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1581.040 4.000 1581.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[33]
  PIN data_arrays_0_0_ext_ram_rdata2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1587.160 4.000 1587.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[34]
  PIN data_arrays_0_0_ext_ram_rdata2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1593.280 4.000 1593.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[35]
  PIN data_arrays_0_0_ext_ram_rdata2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1599.400 4.000 1600.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[36]
  PIN data_arrays_0_0_ext_ram_rdata2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1605.520 4.000 1606.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[37]
  PIN data_arrays_0_0_ext_ram_rdata2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1610.960 4.000 1611.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[38]
  PIN data_arrays_0_0_ext_ram_rdata2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1617.080 4.000 1617.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[39]
  PIN data_arrays_0_0_ext_ram_rdata2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1398.120 4.000 1398.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[3]
  PIN data_arrays_0_0_ext_ram_rdata2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1623.200 4.000 1623.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[40]
  PIN data_arrays_0_0_ext_ram_rdata2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1629.320 4.000 1629.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[41]
  PIN data_arrays_0_0_ext_ram_rdata2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1635.440 4.000 1636.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[42]
  PIN data_arrays_0_0_ext_ram_rdata2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1641.560 4.000 1642.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[43]
  PIN data_arrays_0_0_ext_ram_rdata2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1647.680 4.000 1648.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[44]
  PIN data_arrays_0_0_ext_ram_rdata2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1653.800 4.000 1654.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[45]
  PIN data_arrays_0_0_ext_ram_rdata2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.920 4.000 1660.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[46]
  PIN data_arrays_0_0_ext_ram_rdata2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.040 4.000 1666.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[47]
  PIN data_arrays_0_0_ext_ram_rdata2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1672.160 4.000 1672.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[48]
  PIN data_arrays_0_0_ext_ram_rdata2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1678.280 4.000 1678.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[49]
  PIN data_arrays_0_0_ext_ram_rdata2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.240 4.000 1404.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[4]
  PIN data_arrays_0_0_ext_ram_rdata2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1684.400 4.000 1685.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[50]
  PIN data_arrays_0_0_ext_ram_rdata2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1690.520 4.000 1691.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[51]
  PIN data_arrays_0_0_ext_ram_rdata2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1696.640 4.000 1697.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[52]
  PIN data_arrays_0_0_ext_ram_rdata2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1702.760 4.000 1703.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[53]
  PIN data_arrays_0_0_ext_ram_rdata2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1708.880 4.000 1709.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[54]
  PIN data_arrays_0_0_ext_ram_rdata2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.000 4.000 1715.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[55]
  PIN data_arrays_0_0_ext_ram_rdata2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1721.120 4.000 1721.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[56]
  PIN data_arrays_0_0_ext_ram_rdata2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[57]
  PIN data_arrays_0_0_ext_ram_rdata2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1733.360 4.000 1733.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[58]
  PIN data_arrays_0_0_ext_ram_rdata2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1739.480 4.000 1740.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[59]
  PIN data_arrays_0_0_ext_ram_rdata2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1410.360 4.000 1410.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[5]
  PIN data_arrays_0_0_ext_ram_rdata2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1745.600 4.000 1746.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[60]
  PIN data_arrays_0_0_ext_ram_rdata2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.720 4.000 1752.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[61]
  PIN data_arrays_0_0_ext_ram_rdata2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.840 4.000 1758.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[62]
  PIN data_arrays_0_0_ext_ram_rdata2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1763.960 4.000 1764.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[63]
  PIN data_arrays_0_0_ext_ram_rdata2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1416.480 4.000 1417.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[6]
  PIN data_arrays_0_0_ext_ram_rdata2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1422.600 4.000 1423.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[7]
  PIN data_arrays_0_0_ext_ram_rdata2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.720 4.000 1429.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[8]
  PIN data_arrays_0_0_ext_ram_rdata2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.840 4.000 1435.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[9]
  PIN data_arrays_0_0_ext_ram_rdata3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.070 1763.100 1363.350 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[0]
  PIN data_arrays_0_0_ext_ram_rdata3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.170 1763.100 1425.450 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[10]
  PIN data_arrays_0_0_ext_ram_rdata3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.150 1763.100 1431.430 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[11]
  PIN data_arrays_0_0_ext_ram_rdata3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.130 1763.100 1437.410 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[12]
  PIN data_arrays_0_0_ext_ram_rdata3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.570 1763.100 1443.850 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[13]
  PIN data_arrays_0_0_ext_ram_rdata3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.550 1763.100 1449.830 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[14]
  PIN data_arrays_0_0_ext_ram_rdata3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 1763.100 1456.270 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[15]
  PIN data_arrays_0_0_ext_ram_rdata3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 1763.100 1462.250 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[16]
  PIN data_arrays_0_0_ext_ram_rdata3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 1763.100 1468.690 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[17]
  PIN data_arrays_0_0_ext_ram_rdata3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.390 1763.100 1474.670 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[18]
  PIN data_arrays_0_0_ext_ram_rdata3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.830 1763.100 1481.110 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[19]
  PIN data_arrays_0_0_ext_ram_rdata3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.510 1763.100 1369.790 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[1]
  PIN data_arrays_0_0_ext_ram_rdata3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.810 1763.100 1487.090 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[20]
  PIN data_arrays_0_0_ext_ram_rdata3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 1763.100 1493.070 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[21]
  PIN data_arrays_0_0_ext_ram_rdata3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.230 1763.100 1499.510 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[22]
  PIN data_arrays_0_0_ext_ram_rdata3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1505.210 1763.100 1505.490 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[23]
  PIN data_arrays_0_0_ext_ram_rdata3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.650 1763.100 1511.930 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[24]
  PIN data_arrays_0_0_ext_ram_rdata3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.630 1763.100 1517.910 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[25]
  PIN data_arrays_0_0_ext_ram_rdata3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.070 1763.100 1524.350 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[26]
  PIN data_arrays_0_0_ext_ram_rdata3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.050 1763.100 1530.330 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[27]
  PIN data_arrays_0_0_ext_ram_rdata3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.490 1763.100 1536.770 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[28]
  PIN data_arrays_0_0_ext_ram_rdata3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 1763.100 1542.750 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[29]
  PIN data_arrays_0_0_ext_ram_rdata3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.490 1763.100 1375.770 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[2]
  PIN data_arrays_0_0_ext_ram_rdata3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.450 1763.100 1548.730 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[30]
  PIN data_arrays_0_0_ext_ram_rdata3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.890 1763.100 1555.170 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[31]
  PIN data_arrays_0_0_ext_ram_rdata3[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.870 1763.100 1561.150 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[32]
  PIN data_arrays_0_0_ext_ram_rdata3[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.310 1763.100 1567.590 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[33]
  PIN data_arrays_0_0_ext_ram_rdata3[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.290 1763.100 1573.570 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[34]
  PIN data_arrays_0_0_ext_ram_rdata3[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.730 1763.100 1580.010 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[35]
  PIN data_arrays_0_0_ext_ram_rdata3[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.710 1763.100 1585.990 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[36]
  PIN data_arrays_0_0_ext_ram_rdata3[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.150 1763.100 1592.430 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[37]
  PIN data_arrays_0_0_ext_ram_rdata3[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.130 1763.100 1598.410 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[38]
  PIN data_arrays_0_0_ext_ram_rdata3[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.110 1763.100 1604.390 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[39]
  PIN data_arrays_0_0_ext_ram_rdata3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 1763.100 1381.750 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[3]
  PIN data_arrays_0_0_ext_ram_rdata3[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.550 1763.100 1610.830 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[40]
  PIN data_arrays_0_0_ext_ram_rdata3[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 1763.100 1616.810 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[41]
  PIN data_arrays_0_0_ext_ram_rdata3[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 1763.100 1623.250 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[42]
  PIN data_arrays_0_0_ext_ram_rdata3[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.950 1763.100 1629.230 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[43]
  PIN data_arrays_0_0_ext_ram_rdata3[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.390 1763.100 1635.670 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[44]
  PIN data_arrays_0_0_ext_ram_rdata3[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.370 1763.100 1641.650 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[45]
  PIN data_arrays_0_0_ext_ram_rdata3[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.810 1763.100 1648.090 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[46]
  PIN data_arrays_0_0_ext_ram_rdata3[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.790 1763.100 1654.070 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[47]
  PIN data_arrays_0_0_ext_ram_rdata3[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1659.770 1763.100 1660.050 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[48]
  PIN data_arrays_0_0_ext_ram_rdata3[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.210 1763.100 1666.490 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[49]
  PIN data_arrays_0_0_ext_ram_rdata3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 1763.100 1388.190 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[4]
  PIN data_arrays_0_0_ext_ram_rdata3[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 1763.100 1672.470 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[50]
  PIN data_arrays_0_0_ext_ram_rdata3[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.630 1763.100 1678.910 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[51]
  PIN data_arrays_0_0_ext_ram_rdata3[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.610 1763.100 1684.890 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[52]
  PIN data_arrays_0_0_ext_ram_rdata3[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.050 1763.100 1691.330 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[53]
  PIN data_arrays_0_0_ext_ram_rdata3[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.030 1763.100 1697.310 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[54]
  PIN data_arrays_0_0_ext_ram_rdata3[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 1763.100 1703.750 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[55]
  PIN data_arrays_0_0_ext_ram_rdata3[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.450 1763.100 1709.730 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[56]
  PIN data_arrays_0_0_ext_ram_rdata3[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.430 1763.100 1715.710 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[57]
  PIN data_arrays_0_0_ext_ram_rdata3[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.870 1763.100 1722.150 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[58]
  PIN data_arrays_0_0_ext_ram_rdata3[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.850 1763.100 1728.130 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[59]
  PIN data_arrays_0_0_ext_ram_rdata3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.890 1763.100 1394.170 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[5]
  PIN data_arrays_0_0_ext_ram_rdata3[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.290 1763.100 1734.570 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[60]
  PIN data_arrays_0_0_ext_ram_rdata3[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.270 1763.100 1740.550 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[61]
  PIN data_arrays_0_0_ext_ram_rdata3[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.710 1763.100 1746.990 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[62]
  PIN data_arrays_0_0_ext_ram_rdata3[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.690 1763.100 1752.970 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[63]
  PIN data_arrays_0_0_ext_ram_rdata3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.330 1763.100 1400.610 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[6]
  PIN data_arrays_0_0_ext_ram_rdata3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.310 1763.100 1406.590 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[7]
  PIN data_arrays_0_0_ext_ram_rdata3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.750 1763.100 1413.030 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[8]
  PIN data_arrays_0_0_ext_ram_rdata3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 1763.100 1419.010 1767.100 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[9]
  PIN data_arrays_0_0_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[0]
  PIN data_arrays_0_0_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata[10]
  PIN data_arrays_0_0_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata[11]
  PIN data_arrays_0_0_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata[12]
  PIN data_arrays_0_0_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 532.480 4.000 533.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[13]
  PIN data_arrays_0_0_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[14]
  PIN data_arrays_0_0_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[15]
  PIN data_arrays_0_0_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata[16]
  PIN data_arrays_0_0_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata[17]
  PIN data_arrays_0_0_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[18]
  PIN data_arrays_0_0_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.200 4.000 569.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[19]
  PIN data_arrays_0_0_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[1]
  PIN data_arrays_0_0_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[20]
  PIN data_arrays_0_0_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata[21]
  PIN data_arrays_0_0_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[22]
  PIN data_arrays_0_0_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 4.000 594.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata[23]
  PIN data_arrays_0_0_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[24]
  PIN data_arrays_0_0_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[25]
  PIN data_arrays_0_0_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata[26]
  PIN data_arrays_0_0_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.160 4.000 618.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[27]
  PIN data_arrays_0_0_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata[28]
  PIN data_arrays_0_0_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[29]
  PIN data_arrays_0_0_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata[2]
  PIN data_arrays_0_0_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[30]
  PIN data_arrays_0_0_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[31]
  PIN data_arrays_0_0_ext_ram_wdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 4.000 648.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[32]
  PIN data_arrays_0_0_ext_ram_wdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[33]
  PIN data_arrays_0_0_ext_ram_wdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[34]
  PIN data_arrays_0_0_ext_ram_wdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata[35]
  PIN data_arrays_0_0_ext_ram_wdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 672.560 4.000 673.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[36]
  PIN data_arrays_0_0_ext_ram_wdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata[37]
  PIN data_arrays_0_0_ext_ram_wdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[38]
  PIN data_arrays_0_0_ext_ram_wdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[39]
  PIN data_arrays_0_0_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata[3]
  PIN data_arrays_0_0_ext_ram_wdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata[40]
  PIN data_arrays_0_0_ext_ram_wdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[41]
  PIN data_arrays_0_0_ext_ram_wdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.280 4.000 709.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata[42]
  PIN data_arrays_0_0_ext_ram_wdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[43]
  PIN data_arrays_0_0_ext_ram_wdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 721.520 4.000 722.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[44]
  PIN data_arrays_0_0_ext_ram_wdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[45]
  PIN data_arrays_0_0_ext_ram_wdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.760 4.000 734.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata[46]
  PIN data_arrays_0_0_ext_ram_wdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[47]
  PIN data_arrays_0_0_ext_ram_wdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.000 4.000 746.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[48]
  PIN data_arrays_0_0_ext_ram_wdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata[49]
  PIN data_arrays_0_0_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[4]
  PIN data_arrays_0_0_ext_ram_wdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata[50]
  PIN data_arrays_0_0_ext_ram_wdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata[51]
  PIN data_arrays_0_0_ext_ram_wdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 770.480 4.000 771.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[52]
  PIN data_arrays_0_0_ext_ram_wdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[53]
  PIN data_arrays_0_0_ext_ram_wdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[54]
  PIN data_arrays_0_0_ext_ram_wdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata[55]
  PIN data_arrays_0_0_ext_ram_wdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.960 4.000 795.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata[56]
  PIN data_arrays_0_0_ext_ram_wdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[57]
  PIN data_arrays_0_0_ext_ram_wdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 806.520 4.000 807.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[58]
  PIN data_arrays_0_0_ext_ram_wdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[59]
  PIN data_arrays_0_0_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[5]
  PIN data_arrays_0_0_ext_ram_wdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.760 4.000 819.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata[60]
  PIN data_arrays_0_0_ext_ram_wdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.880 4.000 825.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[61]
  PIN data_arrays_0_0_ext_ram_wdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.000 4.000 831.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[62]
  PIN data_arrays_0_0_ext_ram_wdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.120 4.000 837.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata[63]
  PIN data_arrays_0_0_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[6]
  PIN data_arrays_0_0_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.760 4.000 496.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata[7]
  PIN data_arrays_0_0_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[8]
  PIN data_arrays_0_0_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[9]
  PIN data_arrays_0_0_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.960 4.000 880.560 ;
    END
  END data_arrays_0_0_ext_ram_web
  PIN data_arrays_0_0_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END data_arrays_0_0_ext_ram_wmask[0]
  PIN data_arrays_0_0_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 849.360 4.000 849.960 ;
    END
  END data_arrays_0_0_ext_ram_wmask[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 19.080 1756.380 19.680 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1196.840 1756.380 1197.440 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1314.480 1756.380 1315.080 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1432.800 1756.380 1433.400 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1550.440 1756.380 1551.040 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1668.080 1756.380 1668.680 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.670 1763.100 1344.950 1767.100 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.810 1763.100 1326.090 1767.100 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 1763.100 1307.690 1767.100 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 1763.100 1289.290 1767.100 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1270.150 1763.100 1270.430 1767.100 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 136.720 1756.380 137.320 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.750 1763.100 1252.030 1767.100 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1763.100 1233.630 1767.100 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 1763.100 1214.770 1767.100 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.090 1763.100 1196.370 1767.100 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.690 1763.100 1177.970 1767.100 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.830 1763.100 1159.110 1767.100 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.430 1763.100 1140.710 1767.100 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.030 1763.100 1122.310 1767.100 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.170 1763.100 1103.450 1767.100 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.770 1763.100 1085.050 1767.100 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 254.360 1756.380 254.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 1763.100 1066.650 1767.100 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 1763.100 1047.790 1767.100 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 1763.100 1029.390 1767.100 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.710 1763.100 1010.990 1767.100 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 1763.100 992.130 1767.100 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.450 1763.100 973.730 1767.100 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 1763.100 955.330 1767.100 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 1763.100 936.470 1767.100 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 372.000 1756.380 372.600 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 490.320 1756.380 490.920 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 607.960 1756.380 608.560 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 725.600 1756.380 726.200 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 843.240 1756.380 843.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 961.560 1756.380 962.160 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1079.200 1756.380 1079.800 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 57.840 1756.380 58.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1236.280 1756.380 1236.880 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1353.920 1756.380 1354.520 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1471.560 1756.380 1472.160 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1589.880 1756.380 1590.480 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1707.520 1756.380 1708.120 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.650 1763.100 1350.930 1767.100 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.250 1763.100 1332.530 1767.100 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 1763.100 1314.130 1767.100 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.990 1763.100 1295.270 1767.100 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.590 1763.100 1276.870 1767.100 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 176.160 1756.380 176.760 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.190 1763.100 1258.470 1767.100 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.330 1763.100 1239.610 1767.100 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.930 1763.100 1221.210 1767.100 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.530 1763.100 1202.810 1767.100 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 1763.100 1183.950 1767.100 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.270 1763.100 1165.550 1767.100 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.870 1763.100 1147.150 1767.100 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 1763.100 1128.290 1767.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 1763.100 1109.890 1767.100 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 1763.100 1091.490 1767.100 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 293.800 1756.380 294.400 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1763.100 1072.630 1767.100 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 1763.100 1054.230 1767.100 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.550 1763.100 1035.830 1767.100 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 1763.100 1016.970 1767.100 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 1763.100 998.570 1767.100 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 1763.100 980.170 1767.100 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 1763.100 961.310 1767.100 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 1763.100 942.910 1767.100 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 411.440 1756.380 412.040 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 529.080 1756.380 529.680 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 647.400 1756.380 648.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 765.040 1756.380 765.640 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 882.680 1756.380 883.280 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1000.320 1756.380 1000.920 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1118.640 1756.380 1119.240 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 97.280 1756.380 97.880 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1275.720 1756.380 1276.320 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1393.360 1756.380 1393.960 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1511.000 1756.380 1511.600 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1628.640 1756.380 1629.240 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1746.960 1756.380 1747.560 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.090 1763.100 1357.370 1767.100 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.230 1763.100 1338.510 1767.100 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.830 1763.100 1320.110 1767.100 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 1763.100 1301.710 1767.100 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.570 1763.100 1282.850 1767.100 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 214.920 1756.380 215.520 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 1763.100 1264.450 1767.100 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.770 1763.100 1246.050 1767.100 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 1763.100 1227.190 1767.100 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 1763.100 1208.790 1767.100 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.110 1763.100 1190.390 1767.100 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.250 1763.100 1171.530 1767.100 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 1763.100 1153.130 1767.100 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 1763.100 1134.730 1767.100 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.590 1763.100 1115.870 1767.100 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.190 1763.100 1097.470 1767.100 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 333.240 1756.380 333.840 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 1763.100 1079.070 1767.100 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 1763.100 1060.210 1767.100 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.530 1763.100 1041.810 1767.100 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 1763.100 1023.410 1767.100 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.270 1763.100 1004.550 1767.100 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.870 1763.100 986.150 1767.100 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 1763.100 967.750 1767.100 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 1763.100 948.890 1767.100 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 450.880 1756.380 451.480 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 568.520 1756.380 569.120 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 686.160 1756.380 686.760 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 804.480 1756.380 805.080 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 922.120 1756.380 922.720 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1039.760 1756.380 1040.360 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1752.380 1157.400 1756.380 1158.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.710 0.000 1746.990 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.390 0.000 1750.670 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.070 0.000 1754.350 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.710 0.000 1447.990 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.290 0.000 1458.570 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.870 0.000 1469.150 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.450 0.000 1479.730 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 0.000 1490.770 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.070 0.000 1501.350 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.650 0.000 1511.930 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.230 0.000 1522.510 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.270 0.000 1533.550 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.850 0.000 1544.130 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.430 0.000 1554.710 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 0.000 1565.290 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.050 0.000 1576.330 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.630 0.000 1586.910 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 0.000 1597.490 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.790 0.000 1608.070 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.370 0.000 1618.650 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.410 0.000 1629.690 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.990 0.000 1640.270 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.570 0.000 1650.850 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.150 0.000 1661.430 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 0.000 1672.470 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.770 0.000 1683.050 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.350 0.000 1693.630 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.930 0.000 1704.210 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.970 0.000 1715.250 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.550 0.000 1725.830 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.130 0.000 1736.410 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 0.000 753.390 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 0.000 774.550 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 0.000 806.750 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.250 0.000 849.530 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.190 0.000 913.470 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 0.000 924.050 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 0.000 956.250 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 0.000 966.830 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 0.000 988.450 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 0.000 1020.190 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 0.000 1031.230 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.530 0.000 1041.810 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 0.000 1052.390 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 0.000 1074.010 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 0.000 1084.590 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.470 0.000 1105.750 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 0.000 1116.790 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.670 0.000 1137.950 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.250 0.000 1148.530 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.830 0.000 1159.110 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 0.000 1170.150 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.450 0.000 1180.730 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.030 0.000 1191.310 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.610 0.000 1201.890 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.650 0.000 1212.930 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.230 0.000 1223.510 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 0.000 1234.090 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.390 0.000 1244.670 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.430 0.000 1255.710 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.590 0.000 1276.870 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.170 0.000 1287.450 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.790 0.000 1309.070 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 0.000 1319.650 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.530 0.000 1340.810 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.570 0.000 1351.850 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 0.000 1362.430 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.730 0.000 1373.010 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.310 0.000 1383.590 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.930 0.000 1405.210 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.510 0.000 1415.790 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.090 0.000 1426.370 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.130 0.000 1437.410 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.930 0.000 1451.210 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 0.000 1462.250 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.550 0.000 1472.830 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.130 0.000 1483.410 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.710 0.000 1493.990 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.750 0.000 1505.030 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.330 0.000 1515.610 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.910 0.000 1526.190 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.490 0.000 1536.770 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.530 0.000 1547.810 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.110 0.000 1558.390 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.690 0.000 1568.970 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.270 0.000 1579.550 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.310 0.000 1590.590 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.890 0.000 1601.170 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.050 0.000 1622.330 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 0.000 1632.910 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.670 0.000 1643.950 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.250 0.000 1654.530 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.830 0.000 1665.110 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.410 0.000 1675.690 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.450 0.000 1686.730 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.030 0.000 1697.310 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1707.610 0.000 1707.890 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 0.000 1718.470 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 0.000 1729.510 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.810 0.000 1740.090 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 0.000 639.310 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 0.000 703.250 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 0.000 735.450 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 0.000 746.030 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 0.000 756.610 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 0.000 799.390 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 0.000 821.010 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 0.000 852.750 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 0.000 874.370 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 0.000 884.950 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.290 0.000 906.570 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 0.000 938.310 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 0.000 949.350 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 0.000 970.510 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 0.000 981.090 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 0.000 991.670 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 0.000 1023.870 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 0.000 1034.450 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.210 0.000 1045.490 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 0.000 1066.650 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 0.000 1077.230 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.990 0.000 1088.270 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 0.000 1109.430 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.730 0.000 1120.010 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 0.000 1141.630 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 0.000 1173.370 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.130 0.000 1184.410 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 0.000 1194.990 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290 0.000 1205.570 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.870 0.000 1216.150 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.490 0.000 1237.770 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.070 0.000 1248.350 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.650 0.000 1258.930 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 0.000 1269.970 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 0.000 1280.550 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.850 0.000 1291.130 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 0.000 1301.710 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.010 0.000 1312.290 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 0.000 1323.330 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 0.000 1333.910 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 0.000 1344.490 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.790 0.000 1355.070 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.830 0.000 1366.110 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.410 0.000 1376.690 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.990 0.000 1387.270 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 0.000 1397.850 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.610 0.000 1408.890 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.190 0.000 1419.470 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.350 0.000 1440.630 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.610 0.000 1454.890 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 0.000 1465.470 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.230 0.000 1476.510 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.810 0.000 1487.090 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 0.000 1497.670 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.970 0.000 1508.250 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.010 0.000 1519.290 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 0.000 1529.870 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.170 0.000 1540.450 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.750 0.000 1551.030 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 0.000 1562.070 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.370 0.000 1572.650 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.950 0.000 1583.230 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.530 0.000 1593.810 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.110 0.000 1604.390 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.150 0.000 1615.430 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 0.000 1626.010 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.310 0.000 1636.590 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.890 0.000 1647.170 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.930 0.000 1658.210 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.510 0.000 1668.790 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.090 0.000 1679.370 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.670 0.000 1689.950 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.710 0.000 1700.990 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.290 0.000 1711.570 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.870 0.000 1722.150 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 0.000 1732.730 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.490 0.000 1743.770 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 0.000 642.530 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 0.000 685.310 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 0.000 717.510 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 0.000 781.910 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 0.000 803.070 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 0.000 813.650 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 0.000 824.230 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 0.000 835.270 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 0.000 856.430 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 0.000 878.050 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 0.000 899.210 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 0.000 920.830 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 0.000 931.410 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.710 0.000 941.990 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 0.000 952.570 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.910 0.000 974.190 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 0.000 984.770 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.650 0.000 1005.930 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 0.000 1038.130 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 0.000 1070.330 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 0.000 1080.910 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.830 0.000 1113.110 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.410 0.000 1123.690 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.990 0.000 1134.270 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.570 0.000 1144.850 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.610 0.000 1155.890 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.190 0.000 1166.470 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.350 0.000 1187.630 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 0.000 1198.670 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 0.000 1209.250 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 0.000 1219.830 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 0.000 1230.410 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.750 0.000 1252.030 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.910 0.000 1273.190 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.490 0.000 1283.770 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.110 0.000 1305.390 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.690 0.000 1315.970 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.270 0.000 1326.550 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.310 0.000 1337.590 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.890 0.000 1348.170 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.470 0.000 1358.750 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.050 0.000 1369.330 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 0.000 1380.370 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.670 0.000 1390.950 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.250 0.000 1401.530 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.830 0.000 1412.110 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.450 0.000 1433.730 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.030 0.000 1444.310 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END la_oenb[9]
  PIN tag_array_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1763.100 689.450 1767.100 ;
    END
  END tag_array_ext_ram_addr1[0]
  PIN tag_array_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 1763.100 695.430 1767.100 ;
    END
  END tag_array_ext_ram_addr1[1]
  PIN tag_array_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 1763.100 701.870 1767.100 ;
    END
  END tag_array_ext_ram_addr1[2]
  PIN tag_array_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 1763.100 707.850 1767.100 ;
    END
  END tag_array_ext_ram_addr1[3]
  PIN tag_array_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 1763.100 714.290 1767.100 ;
    END
  END tag_array_ext_ram_addr1[4]
  PIN tag_array_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 1763.100 720.270 1767.100 ;
    END
  END tag_array_ext_ram_addr1[5]
  PIN tag_array_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 1763.100 726.250 1767.100 ;
    END
  END tag_array_ext_ram_addr1[6]
  PIN tag_array_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 1763.100 732.690 1767.100 ;
    END
  END tag_array_ext_ram_addr1[7]
  PIN tag_array_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 1763.100 200.930 1767.100 ;
    END
  END tag_array_ext_ram_addr[0]
  PIN tag_array_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 1763.100 206.910 1767.100 ;
    END
  END tag_array_ext_ram_addr[1]
  PIN tag_array_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 1763.100 213.350 1767.100 ;
    END
  END tag_array_ext_ram_addr[2]
  PIN tag_array_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 1763.100 219.330 1767.100 ;
    END
  END tag_array_ext_ram_addr[3]
  PIN tag_array_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 1763.100 225.310 1767.100 ;
    END
  END tag_array_ext_ram_addr[4]
  PIN tag_array_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 1763.100 231.750 1767.100 ;
    END
  END tag_array_ext_ram_addr[5]
  PIN tag_array_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 1763.100 237.730 1767.100 ;
    END
  END tag_array_ext_ram_addr[6]
  PIN tag_array_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 1763.100 244.170 1767.100 ;
    END
  END tag_array_ext_ram_addr[7]
  PIN tag_array_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 1763.100 250.150 1767.100 ;
    END
  END tag_array_ext_ram_clk
  PIN tag_array_ext_ram_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 1763.100 664.610 1767.100 ;
    END
  END tag_array_ext_ram_csb
  PIN tag_array_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 1763.100 677.030 1767.100 ;
    END
  END tag_array_ext_ram_csb1[0]
  PIN tag_array_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 1763.100 683.010 1767.100 ;
    END
  END tag_array_ext_ram_csb1[1]
  PIN tag_array_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 1763.100 3.130 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[0]
  PIN tag_array_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1763.100 64.770 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[10]
  PIN tag_array_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 1763.100 70.750 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[11]
  PIN tag_array_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 1763.100 77.190 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[12]
  PIN tag_array_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 1763.100 83.170 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[13]
  PIN tag_array_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 1763.100 89.610 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[14]
  PIN tag_array_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 1763.100 95.590 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[15]
  PIN tag_array_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 1763.100 102.030 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[16]
  PIN tag_array_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 1763.100 108.010 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[17]
  PIN tag_array_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 1763.100 113.990 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[18]
  PIN tag_array_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 1763.100 120.430 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[19]
  PIN tag_array_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 1763.100 9.110 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[1]
  PIN tag_array_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 1763.100 126.410 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[20]
  PIN tag_array_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 1763.100 132.850 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[21]
  PIN tag_array_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 1763.100 138.830 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[22]
  PIN tag_array_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1763.100 145.270 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[23]
  PIN tag_array_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 1763.100 151.250 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[24]
  PIN tag_array_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 1763.100 157.690 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[25]
  PIN tag_array_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 1763.100 163.670 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[26]
  PIN tag_array_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 1763.100 169.650 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[27]
  PIN tag_array_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 1763.100 176.090 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[28]
  PIN tag_array_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 1763.100 182.070 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[29]
  PIN tag_array_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 1763.100 15.090 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[2]
  PIN tag_array_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 1763.100 188.510 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[30]
  PIN tag_array_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 1763.100 194.490 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[31]
  PIN tag_array_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 1763.100 21.530 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[3]
  PIN tag_array_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 1763.100 27.510 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[4]
  PIN tag_array_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 1763.100 33.950 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[5]
  PIN tag_array_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 1763.100 39.930 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[6]
  PIN tag_array_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 1763.100 46.370 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[7]
  PIN tag_array_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 1763.100 52.350 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[8]
  PIN tag_array_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1763.100 58.330 1767.100 ;
    END
  END tag_array_ext_ram_rdata0[9]
  PIN tag_array_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 1763.100 738.670 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[0]
  PIN tag_array_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 1763.100 800.770 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[10]
  PIN tag_array_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 1763.100 806.750 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[11]
  PIN tag_array_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.910 1763.100 813.190 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[12]
  PIN tag_array_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 1763.100 819.170 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[13]
  PIN tag_array_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 1763.100 825.610 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[14]
  PIN tag_array_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 1763.100 831.590 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[15]
  PIN tag_array_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 1763.100 837.570 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[16]
  PIN tag_array_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 1763.100 844.010 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[17]
  PIN tag_array_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 1763.100 849.990 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[18]
  PIN tag_array_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 1763.100 856.430 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[19]
  PIN tag_array_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 1763.100 745.110 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[1]
  PIN tag_array_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 1763.100 862.410 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[20]
  PIN tag_array_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 1763.100 868.850 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[21]
  PIN tag_array_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 1763.100 874.830 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[22]
  PIN tag_array_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 1763.100 881.270 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[23]
  PIN tag_array_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 1763.100 887.250 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[24]
  PIN tag_array_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 1763.100 893.230 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[25]
  PIN tag_array_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 1763.100 899.670 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[26]
  PIN tag_array_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 1763.100 905.650 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[27]
  PIN tag_array_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 1763.100 912.090 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[28]
  PIN tag_array_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 1763.100 918.070 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[29]
  PIN tag_array_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 1763.100 751.090 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[2]
  PIN tag_array_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 1763.100 924.510 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[30]
  PIN tag_array_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 1763.100 930.490 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[31]
  PIN tag_array_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 1763.100 757.530 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[3]
  PIN tag_array_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1763.100 763.510 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[4]
  PIN tag_array_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 1763.100 769.950 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[5]
  PIN tag_array_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 1763.100 775.930 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[6]
  PIN tag_array_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 1763.100 781.910 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[7]
  PIN tag_array_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 1763.100 788.350 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[8]
  PIN tag_array_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 1763.100 794.330 1767.100 ;
    END
  END tag_array_ext_ram_rdata1[9]
  PIN tag_array_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 1763.100 256.590 1767.100 ;
    END
  END tag_array_ext_ram_wdata[0]
  PIN tag_array_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 1763.100 318.230 1767.100 ;
    END
  END tag_array_ext_ram_wdata[10]
  PIN tag_array_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 1763.100 324.670 1767.100 ;
    END
  END tag_array_ext_ram_wdata[11]
  PIN tag_array_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 1763.100 330.650 1767.100 ;
    END
  END tag_array_ext_ram_wdata[12]
  PIN tag_array_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 1763.100 336.630 1767.100 ;
    END
  END tag_array_ext_ram_wdata[13]
  PIN tag_array_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 1763.100 343.070 1767.100 ;
    END
  END tag_array_ext_ram_wdata[14]
  PIN tag_array_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 1763.100 349.050 1767.100 ;
    END
  END tag_array_ext_ram_wdata[15]
  PIN tag_array_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 1763.100 355.490 1767.100 ;
    END
  END tag_array_ext_ram_wdata[16]
  PIN tag_array_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 1763.100 361.470 1767.100 ;
    END
  END tag_array_ext_ram_wdata[17]
  PIN tag_array_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 1763.100 367.910 1767.100 ;
    END
  END tag_array_ext_ram_wdata[18]
  PIN tag_array_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 1763.100 373.890 1767.100 ;
    END
  END tag_array_ext_ram_wdata[19]
  PIN tag_array_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 1763.100 262.570 1767.100 ;
    END
  END tag_array_ext_ram_wdata[1]
  PIN tag_array_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 1763.100 380.330 1767.100 ;
    END
  END tag_array_ext_ram_wdata[20]
  PIN tag_array_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 1763.100 386.310 1767.100 ;
    END
  END tag_array_ext_ram_wdata[21]
  PIN tag_array_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 1763.100 392.290 1767.100 ;
    END
  END tag_array_ext_ram_wdata[22]
  PIN tag_array_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 1763.100 398.730 1767.100 ;
    END
  END tag_array_ext_ram_wdata[23]
  PIN tag_array_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 1763.100 404.710 1767.100 ;
    END
  END tag_array_ext_ram_wdata[24]
  PIN tag_array_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 1763.100 411.150 1767.100 ;
    END
  END tag_array_ext_ram_wdata[25]
  PIN tag_array_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 1763.100 417.130 1767.100 ;
    END
  END tag_array_ext_ram_wdata[26]
  PIN tag_array_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 1763.100 423.570 1767.100 ;
    END
  END tag_array_ext_ram_wdata[27]
  PIN tag_array_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 1763.100 429.550 1767.100 ;
    END
  END tag_array_ext_ram_wdata[28]
  PIN tag_array_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 1763.100 435.990 1767.100 ;
    END
  END tag_array_ext_ram_wdata[29]
  PIN tag_array_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 1763.100 269.010 1767.100 ;
    END
  END tag_array_ext_ram_wdata[2]
  PIN tag_array_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 1763.100 441.970 1767.100 ;
    END
  END tag_array_ext_ram_wdata[30]
  PIN tag_array_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 1763.100 447.950 1767.100 ;
    END
  END tag_array_ext_ram_wdata[31]
  PIN tag_array_ext_ram_wdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1763.100 454.390 1767.100 ;
    END
  END tag_array_ext_ram_wdata[32]
  PIN tag_array_ext_ram_wdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 1763.100 460.370 1767.100 ;
    END
  END tag_array_ext_ram_wdata[33]
  PIN tag_array_ext_ram_wdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 1763.100 466.810 1767.100 ;
    END
  END tag_array_ext_ram_wdata[34]
  PIN tag_array_ext_ram_wdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 1763.100 472.790 1767.100 ;
    END
  END tag_array_ext_ram_wdata[35]
  PIN tag_array_ext_ram_wdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 1763.100 479.230 1767.100 ;
    END
  END tag_array_ext_ram_wdata[36]
  PIN tag_array_ext_ram_wdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 1763.100 485.210 1767.100 ;
    END
  END tag_array_ext_ram_wdata[37]
  PIN tag_array_ext_ram_wdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 1763.100 491.650 1767.100 ;
    END
  END tag_array_ext_ram_wdata[38]
  PIN tag_array_ext_ram_wdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 1763.100 497.630 1767.100 ;
    END
  END tag_array_ext_ram_wdata[39]
  PIN tag_array_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 1763.100 274.990 1767.100 ;
    END
  END tag_array_ext_ram_wdata[3]
  PIN tag_array_ext_ram_wdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 1763.100 503.610 1767.100 ;
    END
  END tag_array_ext_ram_wdata[40]
  PIN tag_array_ext_ram_wdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 1763.100 510.050 1767.100 ;
    END
  END tag_array_ext_ram_wdata[41]
  PIN tag_array_ext_ram_wdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 1763.100 516.030 1767.100 ;
    END
  END tag_array_ext_ram_wdata[42]
  PIN tag_array_ext_ram_wdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 1763.100 522.470 1767.100 ;
    END
  END tag_array_ext_ram_wdata[43]
  PIN tag_array_ext_ram_wdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1763.100 528.450 1767.100 ;
    END
  END tag_array_ext_ram_wdata[44]
  PIN tag_array_ext_ram_wdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 1763.100 534.890 1767.100 ;
    END
  END tag_array_ext_ram_wdata[45]
  PIN tag_array_ext_ram_wdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 1763.100 540.870 1767.100 ;
    END
  END tag_array_ext_ram_wdata[46]
  PIN tag_array_ext_ram_wdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 1763.100 547.310 1767.100 ;
    END
  END tag_array_ext_ram_wdata[47]
  PIN tag_array_ext_ram_wdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 1763.100 553.290 1767.100 ;
    END
  END tag_array_ext_ram_wdata[48]
  PIN tag_array_ext_ram_wdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 1763.100 559.270 1767.100 ;
    END
  END tag_array_ext_ram_wdata[49]
  PIN tag_array_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 1763.100 280.970 1767.100 ;
    END
  END tag_array_ext_ram_wdata[4]
  PIN tag_array_ext_ram_wdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 1763.100 565.710 1767.100 ;
    END
  END tag_array_ext_ram_wdata[50]
  PIN tag_array_ext_ram_wdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 1763.100 571.690 1767.100 ;
    END
  END tag_array_ext_ram_wdata[51]
  PIN tag_array_ext_ram_wdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 1763.100 578.130 1767.100 ;
    END
  END tag_array_ext_ram_wdata[52]
  PIN tag_array_ext_ram_wdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 1763.100 584.110 1767.100 ;
    END
  END tag_array_ext_ram_wdata[53]
  PIN tag_array_ext_ram_wdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 1763.100 590.550 1767.100 ;
    END
  END tag_array_ext_ram_wdata[54]
  PIN tag_array_ext_ram_wdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 1763.100 596.530 1767.100 ;
    END
  END tag_array_ext_ram_wdata[55]
  PIN tag_array_ext_ram_wdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 1763.100 602.970 1767.100 ;
    END
  END tag_array_ext_ram_wdata[56]
  PIN tag_array_ext_ram_wdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 1763.100 608.950 1767.100 ;
    END
  END tag_array_ext_ram_wdata[57]
  PIN tag_array_ext_ram_wdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 1763.100 614.930 1767.100 ;
    END
  END tag_array_ext_ram_wdata[58]
  PIN tag_array_ext_ram_wdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 1763.100 621.370 1767.100 ;
    END
  END tag_array_ext_ram_wdata[59]
  PIN tag_array_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 1763.100 287.410 1767.100 ;
    END
  END tag_array_ext_ram_wdata[5]
  PIN tag_array_ext_ram_wdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 1763.100 627.350 1767.100 ;
    END
  END tag_array_ext_ram_wdata[60]
  PIN tag_array_ext_ram_wdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 1763.100 633.790 1767.100 ;
    END
  END tag_array_ext_ram_wdata[61]
  PIN tag_array_ext_ram_wdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 1763.100 639.770 1767.100 ;
    END
  END tag_array_ext_ram_wdata[62]
  PIN tag_array_ext_ram_wdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 1763.100 646.210 1767.100 ;
    END
  END tag_array_ext_ram_wdata[63]
  PIN tag_array_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 1763.100 293.390 1767.100 ;
    END
  END tag_array_ext_ram_wdata[6]
  PIN tag_array_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1763.100 299.830 1767.100 ;
    END
  END tag_array_ext_ram_wdata[7]
  PIN tag_array_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 1763.100 305.810 1767.100 ;
    END
  END tag_array_ext_ram_wdata[8]
  PIN tag_array_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 1763.100 312.250 1767.100 ;
    END
  END tag_array_ext_ram_wdata[9]
  PIN tag_array_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 1763.100 670.590 1767.100 ;
    END
  END tag_array_ext_ram_web
  PIN tag_array_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 1763.100 652.190 1767.100 ;
    END
  END tag_array_ext_ram_wmask[0]
  PIN tag_array_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 1763.100 658.630 1767.100 ;
    END
  END tag_array_ext_ram_wmask[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1754.640 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1754.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1754.640 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1750.760 1754.485 ;
      LAYER met1 ;
        RECT 1.910 10.640 1754.370 1763.540 ;
      LAYER met2 ;
        RECT 1.470 1762.820 2.570 1766.485 ;
        RECT 3.410 1762.820 8.550 1766.485 ;
        RECT 9.390 1762.820 14.530 1766.485 ;
        RECT 15.370 1762.820 20.970 1766.485 ;
        RECT 21.810 1762.820 26.950 1766.485 ;
        RECT 27.790 1762.820 33.390 1766.485 ;
        RECT 34.230 1762.820 39.370 1766.485 ;
        RECT 40.210 1762.820 45.810 1766.485 ;
        RECT 46.650 1762.820 51.790 1766.485 ;
        RECT 52.630 1762.820 57.770 1766.485 ;
        RECT 58.610 1762.820 64.210 1766.485 ;
        RECT 65.050 1762.820 70.190 1766.485 ;
        RECT 71.030 1762.820 76.630 1766.485 ;
        RECT 77.470 1762.820 82.610 1766.485 ;
        RECT 83.450 1762.820 89.050 1766.485 ;
        RECT 89.890 1762.820 95.030 1766.485 ;
        RECT 95.870 1762.820 101.470 1766.485 ;
        RECT 102.310 1762.820 107.450 1766.485 ;
        RECT 108.290 1762.820 113.430 1766.485 ;
        RECT 114.270 1762.820 119.870 1766.485 ;
        RECT 120.710 1762.820 125.850 1766.485 ;
        RECT 126.690 1762.820 132.290 1766.485 ;
        RECT 133.130 1762.820 138.270 1766.485 ;
        RECT 139.110 1762.820 144.710 1766.485 ;
        RECT 145.550 1762.820 150.690 1766.485 ;
        RECT 151.530 1762.820 157.130 1766.485 ;
        RECT 157.970 1762.820 163.110 1766.485 ;
        RECT 163.950 1762.820 169.090 1766.485 ;
        RECT 169.930 1762.820 175.530 1766.485 ;
        RECT 176.370 1762.820 181.510 1766.485 ;
        RECT 182.350 1762.820 187.950 1766.485 ;
        RECT 188.790 1762.820 193.930 1766.485 ;
        RECT 194.770 1762.820 200.370 1766.485 ;
        RECT 201.210 1762.820 206.350 1766.485 ;
        RECT 207.190 1762.820 212.790 1766.485 ;
        RECT 213.630 1762.820 218.770 1766.485 ;
        RECT 219.610 1762.820 224.750 1766.485 ;
        RECT 225.590 1762.820 231.190 1766.485 ;
        RECT 232.030 1762.820 237.170 1766.485 ;
        RECT 238.010 1762.820 243.610 1766.485 ;
        RECT 244.450 1762.820 249.590 1766.485 ;
        RECT 250.430 1762.820 256.030 1766.485 ;
        RECT 256.870 1762.820 262.010 1766.485 ;
        RECT 262.850 1762.820 268.450 1766.485 ;
        RECT 269.290 1762.820 274.430 1766.485 ;
        RECT 275.270 1762.820 280.410 1766.485 ;
        RECT 281.250 1762.820 286.850 1766.485 ;
        RECT 287.690 1762.820 292.830 1766.485 ;
        RECT 293.670 1762.820 299.270 1766.485 ;
        RECT 300.110 1762.820 305.250 1766.485 ;
        RECT 306.090 1762.820 311.690 1766.485 ;
        RECT 312.530 1762.820 317.670 1766.485 ;
        RECT 318.510 1762.820 324.110 1766.485 ;
        RECT 324.950 1762.820 330.090 1766.485 ;
        RECT 330.930 1762.820 336.070 1766.485 ;
        RECT 336.910 1762.820 342.510 1766.485 ;
        RECT 343.350 1762.820 348.490 1766.485 ;
        RECT 349.330 1762.820 354.930 1766.485 ;
        RECT 355.770 1762.820 360.910 1766.485 ;
        RECT 361.750 1762.820 367.350 1766.485 ;
        RECT 368.190 1762.820 373.330 1766.485 ;
        RECT 374.170 1762.820 379.770 1766.485 ;
        RECT 380.610 1762.820 385.750 1766.485 ;
        RECT 386.590 1762.820 391.730 1766.485 ;
        RECT 392.570 1762.820 398.170 1766.485 ;
        RECT 399.010 1762.820 404.150 1766.485 ;
        RECT 404.990 1762.820 410.590 1766.485 ;
        RECT 411.430 1762.820 416.570 1766.485 ;
        RECT 417.410 1762.820 423.010 1766.485 ;
        RECT 423.850 1762.820 428.990 1766.485 ;
        RECT 429.830 1762.820 435.430 1766.485 ;
        RECT 436.270 1762.820 441.410 1766.485 ;
        RECT 442.250 1762.820 447.390 1766.485 ;
        RECT 448.230 1762.820 453.830 1766.485 ;
        RECT 454.670 1762.820 459.810 1766.485 ;
        RECT 460.650 1762.820 466.250 1766.485 ;
        RECT 467.090 1762.820 472.230 1766.485 ;
        RECT 473.070 1762.820 478.670 1766.485 ;
        RECT 479.510 1762.820 484.650 1766.485 ;
        RECT 485.490 1762.820 491.090 1766.485 ;
        RECT 491.930 1762.820 497.070 1766.485 ;
        RECT 497.910 1762.820 503.050 1766.485 ;
        RECT 503.890 1762.820 509.490 1766.485 ;
        RECT 510.330 1762.820 515.470 1766.485 ;
        RECT 516.310 1762.820 521.910 1766.485 ;
        RECT 522.750 1762.820 527.890 1766.485 ;
        RECT 528.730 1762.820 534.330 1766.485 ;
        RECT 535.170 1762.820 540.310 1766.485 ;
        RECT 541.150 1762.820 546.750 1766.485 ;
        RECT 547.590 1762.820 552.730 1766.485 ;
        RECT 553.570 1762.820 558.710 1766.485 ;
        RECT 559.550 1762.820 565.150 1766.485 ;
        RECT 565.990 1762.820 571.130 1766.485 ;
        RECT 571.970 1762.820 577.570 1766.485 ;
        RECT 578.410 1762.820 583.550 1766.485 ;
        RECT 584.390 1762.820 589.990 1766.485 ;
        RECT 590.830 1762.820 595.970 1766.485 ;
        RECT 596.810 1762.820 602.410 1766.485 ;
        RECT 603.250 1762.820 608.390 1766.485 ;
        RECT 609.230 1762.820 614.370 1766.485 ;
        RECT 615.210 1762.820 620.810 1766.485 ;
        RECT 621.650 1762.820 626.790 1766.485 ;
        RECT 627.630 1762.820 633.230 1766.485 ;
        RECT 634.070 1762.820 639.210 1766.485 ;
        RECT 640.050 1762.820 645.650 1766.485 ;
        RECT 646.490 1762.820 651.630 1766.485 ;
        RECT 652.470 1762.820 658.070 1766.485 ;
        RECT 658.910 1762.820 664.050 1766.485 ;
        RECT 664.890 1762.820 670.030 1766.485 ;
        RECT 670.870 1762.820 676.470 1766.485 ;
        RECT 677.310 1762.820 682.450 1766.485 ;
        RECT 683.290 1762.820 688.890 1766.485 ;
        RECT 689.730 1762.820 694.870 1766.485 ;
        RECT 695.710 1762.820 701.310 1766.485 ;
        RECT 702.150 1762.820 707.290 1766.485 ;
        RECT 708.130 1762.820 713.730 1766.485 ;
        RECT 714.570 1762.820 719.710 1766.485 ;
        RECT 720.550 1762.820 725.690 1766.485 ;
        RECT 726.530 1762.820 732.130 1766.485 ;
        RECT 732.970 1762.820 738.110 1766.485 ;
        RECT 738.950 1762.820 744.550 1766.485 ;
        RECT 745.390 1762.820 750.530 1766.485 ;
        RECT 751.370 1762.820 756.970 1766.485 ;
        RECT 757.810 1762.820 762.950 1766.485 ;
        RECT 763.790 1762.820 769.390 1766.485 ;
        RECT 770.230 1762.820 775.370 1766.485 ;
        RECT 776.210 1762.820 781.350 1766.485 ;
        RECT 782.190 1762.820 787.790 1766.485 ;
        RECT 788.630 1762.820 793.770 1766.485 ;
        RECT 794.610 1762.820 800.210 1766.485 ;
        RECT 801.050 1762.820 806.190 1766.485 ;
        RECT 807.030 1762.820 812.630 1766.485 ;
        RECT 813.470 1762.820 818.610 1766.485 ;
        RECT 819.450 1762.820 825.050 1766.485 ;
        RECT 825.890 1762.820 831.030 1766.485 ;
        RECT 831.870 1762.820 837.010 1766.485 ;
        RECT 837.850 1762.820 843.450 1766.485 ;
        RECT 844.290 1762.820 849.430 1766.485 ;
        RECT 850.270 1762.820 855.870 1766.485 ;
        RECT 856.710 1762.820 861.850 1766.485 ;
        RECT 862.690 1762.820 868.290 1766.485 ;
        RECT 869.130 1762.820 874.270 1766.485 ;
        RECT 875.110 1762.820 880.710 1766.485 ;
        RECT 881.550 1762.820 886.690 1766.485 ;
        RECT 887.530 1762.820 892.670 1766.485 ;
        RECT 893.510 1762.820 899.110 1766.485 ;
        RECT 899.950 1762.820 905.090 1766.485 ;
        RECT 905.930 1762.820 911.530 1766.485 ;
        RECT 912.370 1762.820 917.510 1766.485 ;
        RECT 918.350 1762.820 923.950 1766.485 ;
        RECT 924.790 1762.820 929.930 1766.485 ;
        RECT 930.770 1762.820 935.910 1766.485 ;
        RECT 936.750 1762.820 942.350 1766.485 ;
        RECT 943.190 1762.820 948.330 1766.485 ;
        RECT 949.170 1762.820 954.770 1766.485 ;
        RECT 955.610 1762.820 960.750 1766.485 ;
        RECT 961.590 1762.820 967.190 1766.485 ;
        RECT 968.030 1762.820 973.170 1766.485 ;
        RECT 974.010 1762.820 979.610 1766.485 ;
        RECT 980.450 1762.820 985.590 1766.485 ;
        RECT 986.430 1762.820 991.570 1766.485 ;
        RECT 992.410 1762.820 998.010 1766.485 ;
        RECT 998.850 1762.820 1003.990 1766.485 ;
        RECT 1004.830 1762.820 1010.430 1766.485 ;
        RECT 1011.270 1762.820 1016.410 1766.485 ;
        RECT 1017.250 1762.820 1022.850 1766.485 ;
        RECT 1023.690 1762.820 1028.830 1766.485 ;
        RECT 1029.670 1762.820 1035.270 1766.485 ;
        RECT 1036.110 1762.820 1041.250 1766.485 ;
        RECT 1042.090 1762.820 1047.230 1766.485 ;
        RECT 1048.070 1762.820 1053.670 1766.485 ;
        RECT 1054.510 1762.820 1059.650 1766.485 ;
        RECT 1060.490 1762.820 1066.090 1766.485 ;
        RECT 1066.930 1762.820 1072.070 1766.485 ;
        RECT 1072.910 1762.820 1078.510 1766.485 ;
        RECT 1079.350 1762.820 1084.490 1766.485 ;
        RECT 1085.330 1762.820 1090.930 1766.485 ;
        RECT 1091.770 1762.820 1096.910 1766.485 ;
        RECT 1097.750 1762.820 1102.890 1766.485 ;
        RECT 1103.730 1762.820 1109.330 1766.485 ;
        RECT 1110.170 1762.820 1115.310 1766.485 ;
        RECT 1116.150 1762.820 1121.750 1766.485 ;
        RECT 1122.590 1762.820 1127.730 1766.485 ;
        RECT 1128.570 1762.820 1134.170 1766.485 ;
        RECT 1135.010 1762.820 1140.150 1766.485 ;
        RECT 1140.990 1762.820 1146.590 1766.485 ;
        RECT 1147.430 1762.820 1152.570 1766.485 ;
        RECT 1153.410 1762.820 1158.550 1766.485 ;
        RECT 1159.390 1762.820 1164.990 1766.485 ;
        RECT 1165.830 1762.820 1170.970 1766.485 ;
        RECT 1171.810 1762.820 1177.410 1766.485 ;
        RECT 1178.250 1762.820 1183.390 1766.485 ;
        RECT 1184.230 1762.820 1189.830 1766.485 ;
        RECT 1190.670 1762.820 1195.810 1766.485 ;
        RECT 1196.650 1762.820 1202.250 1766.485 ;
        RECT 1203.090 1762.820 1208.230 1766.485 ;
        RECT 1209.070 1762.820 1214.210 1766.485 ;
        RECT 1215.050 1762.820 1220.650 1766.485 ;
        RECT 1221.490 1762.820 1226.630 1766.485 ;
        RECT 1227.470 1762.820 1233.070 1766.485 ;
        RECT 1233.910 1762.820 1239.050 1766.485 ;
        RECT 1239.890 1762.820 1245.490 1766.485 ;
        RECT 1246.330 1762.820 1251.470 1766.485 ;
        RECT 1252.310 1762.820 1257.910 1766.485 ;
        RECT 1258.750 1762.820 1263.890 1766.485 ;
        RECT 1264.730 1762.820 1269.870 1766.485 ;
        RECT 1270.710 1762.820 1276.310 1766.485 ;
        RECT 1277.150 1762.820 1282.290 1766.485 ;
        RECT 1283.130 1762.820 1288.730 1766.485 ;
        RECT 1289.570 1762.820 1294.710 1766.485 ;
        RECT 1295.550 1762.820 1301.150 1766.485 ;
        RECT 1301.990 1762.820 1307.130 1766.485 ;
        RECT 1307.970 1762.820 1313.570 1766.485 ;
        RECT 1314.410 1762.820 1319.550 1766.485 ;
        RECT 1320.390 1762.820 1325.530 1766.485 ;
        RECT 1326.370 1762.820 1331.970 1766.485 ;
        RECT 1332.810 1762.820 1337.950 1766.485 ;
        RECT 1338.790 1762.820 1344.390 1766.485 ;
        RECT 1345.230 1762.820 1350.370 1766.485 ;
        RECT 1351.210 1762.820 1356.810 1766.485 ;
        RECT 1357.650 1762.820 1362.790 1766.485 ;
        RECT 1363.630 1762.820 1369.230 1766.485 ;
        RECT 1370.070 1762.820 1375.210 1766.485 ;
        RECT 1376.050 1762.820 1381.190 1766.485 ;
        RECT 1382.030 1762.820 1387.630 1766.485 ;
        RECT 1388.470 1762.820 1393.610 1766.485 ;
        RECT 1394.450 1762.820 1400.050 1766.485 ;
        RECT 1400.890 1762.820 1406.030 1766.485 ;
        RECT 1406.870 1762.820 1412.470 1766.485 ;
        RECT 1413.310 1762.820 1418.450 1766.485 ;
        RECT 1419.290 1762.820 1424.890 1766.485 ;
        RECT 1425.730 1762.820 1430.870 1766.485 ;
        RECT 1431.710 1762.820 1436.850 1766.485 ;
        RECT 1437.690 1762.820 1443.290 1766.485 ;
        RECT 1444.130 1762.820 1449.270 1766.485 ;
        RECT 1450.110 1762.820 1455.710 1766.485 ;
        RECT 1456.550 1762.820 1461.690 1766.485 ;
        RECT 1462.530 1762.820 1468.130 1766.485 ;
        RECT 1468.970 1762.820 1474.110 1766.485 ;
        RECT 1474.950 1762.820 1480.550 1766.485 ;
        RECT 1481.390 1762.820 1486.530 1766.485 ;
        RECT 1487.370 1762.820 1492.510 1766.485 ;
        RECT 1493.350 1762.820 1498.950 1766.485 ;
        RECT 1499.790 1762.820 1504.930 1766.485 ;
        RECT 1505.770 1762.820 1511.370 1766.485 ;
        RECT 1512.210 1762.820 1517.350 1766.485 ;
        RECT 1518.190 1762.820 1523.790 1766.485 ;
        RECT 1524.630 1762.820 1529.770 1766.485 ;
        RECT 1530.610 1762.820 1536.210 1766.485 ;
        RECT 1537.050 1762.820 1542.190 1766.485 ;
        RECT 1543.030 1762.820 1548.170 1766.485 ;
        RECT 1549.010 1762.820 1554.610 1766.485 ;
        RECT 1555.450 1762.820 1560.590 1766.485 ;
        RECT 1561.430 1762.820 1567.030 1766.485 ;
        RECT 1567.870 1762.820 1573.010 1766.485 ;
        RECT 1573.850 1762.820 1579.450 1766.485 ;
        RECT 1580.290 1762.820 1585.430 1766.485 ;
        RECT 1586.270 1762.820 1591.870 1766.485 ;
        RECT 1592.710 1762.820 1597.850 1766.485 ;
        RECT 1598.690 1762.820 1603.830 1766.485 ;
        RECT 1604.670 1762.820 1610.270 1766.485 ;
        RECT 1611.110 1762.820 1616.250 1766.485 ;
        RECT 1617.090 1762.820 1622.690 1766.485 ;
        RECT 1623.530 1762.820 1628.670 1766.485 ;
        RECT 1629.510 1762.820 1635.110 1766.485 ;
        RECT 1635.950 1762.820 1641.090 1766.485 ;
        RECT 1641.930 1762.820 1647.530 1766.485 ;
        RECT 1648.370 1762.820 1653.510 1766.485 ;
        RECT 1654.350 1762.820 1659.490 1766.485 ;
        RECT 1660.330 1762.820 1665.930 1766.485 ;
        RECT 1666.770 1762.820 1671.910 1766.485 ;
        RECT 1672.750 1762.820 1678.350 1766.485 ;
        RECT 1679.190 1762.820 1684.330 1766.485 ;
        RECT 1685.170 1762.820 1690.770 1766.485 ;
        RECT 1691.610 1762.820 1696.750 1766.485 ;
        RECT 1697.590 1762.820 1703.190 1766.485 ;
        RECT 1704.030 1762.820 1709.170 1766.485 ;
        RECT 1710.010 1762.820 1715.150 1766.485 ;
        RECT 1715.990 1762.820 1721.590 1766.485 ;
        RECT 1722.430 1762.820 1727.570 1766.485 ;
        RECT 1728.410 1762.820 1734.010 1766.485 ;
        RECT 1734.850 1762.820 1739.990 1766.485 ;
        RECT 1740.830 1762.820 1746.430 1766.485 ;
        RECT 1747.270 1762.820 1752.410 1766.485 ;
        RECT 1753.250 1762.820 1754.340 1766.485 ;
        RECT 1.470 4.280 1754.340 1762.820 ;
        RECT 2.030 2.875 4.410 4.280 ;
        RECT 5.250 2.875 8.090 4.280 ;
        RECT 8.930 2.875 11.770 4.280 ;
        RECT 12.610 2.875 14.990 4.280 ;
        RECT 15.830 2.875 18.670 4.280 ;
        RECT 19.510 2.875 22.350 4.280 ;
        RECT 23.190 2.875 26.030 4.280 ;
        RECT 26.870 2.875 29.250 4.280 ;
        RECT 30.090 2.875 32.930 4.280 ;
        RECT 33.770 2.875 36.610 4.280 ;
        RECT 37.450 2.875 40.290 4.280 ;
        RECT 41.130 2.875 43.510 4.280 ;
        RECT 44.350 2.875 47.190 4.280 ;
        RECT 48.030 2.875 50.870 4.280 ;
        RECT 51.710 2.875 54.550 4.280 ;
        RECT 55.390 2.875 57.770 4.280 ;
        RECT 58.610 2.875 61.450 4.280 ;
        RECT 62.290 2.875 65.130 4.280 ;
        RECT 65.970 2.875 68.810 4.280 ;
        RECT 69.650 2.875 72.030 4.280 ;
        RECT 72.870 2.875 75.710 4.280 ;
        RECT 76.550 2.875 79.390 4.280 ;
        RECT 80.230 2.875 83.070 4.280 ;
        RECT 83.910 2.875 86.290 4.280 ;
        RECT 87.130 2.875 89.970 4.280 ;
        RECT 90.810 2.875 93.650 4.280 ;
        RECT 94.490 2.875 97.330 4.280 ;
        RECT 98.170 2.875 100.550 4.280 ;
        RECT 101.390 2.875 104.230 4.280 ;
        RECT 105.070 2.875 107.910 4.280 ;
        RECT 108.750 2.875 111.590 4.280 ;
        RECT 112.430 2.875 114.810 4.280 ;
        RECT 115.650 2.875 118.490 4.280 ;
        RECT 119.330 2.875 122.170 4.280 ;
        RECT 123.010 2.875 125.850 4.280 ;
        RECT 126.690 2.875 129.070 4.280 ;
        RECT 129.910 2.875 132.750 4.280 ;
        RECT 133.590 2.875 136.430 4.280 ;
        RECT 137.270 2.875 140.110 4.280 ;
        RECT 140.950 2.875 143.330 4.280 ;
        RECT 144.170 2.875 147.010 4.280 ;
        RECT 147.850 2.875 150.690 4.280 ;
        RECT 151.530 2.875 154.370 4.280 ;
        RECT 155.210 2.875 157.590 4.280 ;
        RECT 158.430 2.875 161.270 4.280 ;
        RECT 162.110 2.875 164.950 4.280 ;
        RECT 165.790 2.875 168.170 4.280 ;
        RECT 169.010 2.875 171.850 4.280 ;
        RECT 172.690 2.875 175.530 4.280 ;
        RECT 176.370 2.875 179.210 4.280 ;
        RECT 180.050 2.875 182.430 4.280 ;
        RECT 183.270 2.875 186.110 4.280 ;
        RECT 186.950 2.875 189.790 4.280 ;
        RECT 190.630 2.875 193.470 4.280 ;
        RECT 194.310 2.875 196.690 4.280 ;
        RECT 197.530 2.875 200.370 4.280 ;
        RECT 201.210 2.875 204.050 4.280 ;
        RECT 204.890 2.875 207.730 4.280 ;
        RECT 208.570 2.875 210.950 4.280 ;
        RECT 211.790 2.875 214.630 4.280 ;
        RECT 215.470 2.875 218.310 4.280 ;
        RECT 219.150 2.875 221.990 4.280 ;
        RECT 222.830 2.875 225.210 4.280 ;
        RECT 226.050 2.875 228.890 4.280 ;
        RECT 229.730 2.875 232.570 4.280 ;
        RECT 233.410 2.875 236.250 4.280 ;
        RECT 237.090 2.875 239.470 4.280 ;
        RECT 240.310 2.875 243.150 4.280 ;
        RECT 243.990 2.875 246.830 4.280 ;
        RECT 247.670 2.875 250.510 4.280 ;
        RECT 251.350 2.875 253.730 4.280 ;
        RECT 254.570 2.875 257.410 4.280 ;
        RECT 258.250 2.875 261.090 4.280 ;
        RECT 261.930 2.875 264.770 4.280 ;
        RECT 265.610 2.875 267.990 4.280 ;
        RECT 268.830 2.875 271.670 4.280 ;
        RECT 272.510 2.875 275.350 4.280 ;
        RECT 276.190 2.875 279.030 4.280 ;
        RECT 279.870 2.875 282.250 4.280 ;
        RECT 283.090 2.875 285.930 4.280 ;
        RECT 286.770 2.875 289.610 4.280 ;
        RECT 290.450 2.875 293.290 4.280 ;
        RECT 294.130 2.875 296.510 4.280 ;
        RECT 297.350 2.875 300.190 4.280 ;
        RECT 301.030 2.875 303.870 4.280 ;
        RECT 304.710 2.875 307.550 4.280 ;
        RECT 308.390 2.875 310.770 4.280 ;
        RECT 311.610 2.875 314.450 4.280 ;
        RECT 315.290 2.875 318.130 4.280 ;
        RECT 318.970 2.875 321.350 4.280 ;
        RECT 322.190 2.875 325.030 4.280 ;
        RECT 325.870 2.875 328.710 4.280 ;
        RECT 329.550 2.875 332.390 4.280 ;
        RECT 333.230 2.875 335.610 4.280 ;
        RECT 336.450 2.875 339.290 4.280 ;
        RECT 340.130 2.875 342.970 4.280 ;
        RECT 343.810 2.875 346.650 4.280 ;
        RECT 347.490 2.875 349.870 4.280 ;
        RECT 350.710 2.875 353.550 4.280 ;
        RECT 354.390 2.875 357.230 4.280 ;
        RECT 358.070 2.875 360.910 4.280 ;
        RECT 361.750 2.875 364.130 4.280 ;
        RECT 364.970 2.875 367.810 4.280 ;
        RECT 368.650 2.875 371.490 4.280 ;
        RECT 372.330 2.875 375.170 4.280 ;
        RECT 376.010 2.875 378.390 4.280 ;
        RECT 379.230 2.875 382.070 4.280 ;
        RECT 382.910 2.875 385.750 4.280 ;
        RECT 386.590 2.875 389.430 4.280 ;
        RECT 390.270 2.875 392.650 4.280 ;
        RECT 393.490 2.875 396.330 4.280 ;
        RECT 397.170 2.875 400.010 4.280 ;
        RECT 400.850 2.875 403.690 4.280 ;
        RECT 404.530 2.875 406.910 4.280 ;
        RECT 407.750 2.875 410.590 4.280 ;
        RECT 411.430 2.875 414.270 4.280 ;
        RECT 415.110 2.875 417.950 4.280 ;
        RECT 418.790 2.875 421.170 4.280 ;
        RECT 422.010 2.875 424.850 4.280 ;
        RECT 425.690 2.875 428.530 4.280 ;
        RECT 429.370 2.875 432.210 4.280 ;
        RECT 433.050 2.875 435.430 4.280 ;
        RECT 436.270 2.875 439.110 4.280 ;
        RECT 439.950 2.875 442.790 4.280 ;
        RECT 443.630 2.875 446.470 4.280 ;
        RECT 447.310 2.875 449.690 4.280 ;
        RECT 450.530 2.875 453.370 4.280 ;
        RECT 454.210 2.875 457.050 4.280 ;
        RECT 457.890 2.875 460.730 4.280 ;
        RECT 461.570 2.875 463.950 4.280 ;
        RECT 464.790 2.875 467.630 4.280 ;
        RECT 468.470 2.875 471.310 4.280 ;
        RECT 472.150 2.875 474.990 4.280 ;
        RECT 475.830 2.875 478.210 4.280 ;
        RECT 479.050 2.875 481.890 4.280 ;
        RECT 482.730 2.875 485.570 4.280 ;
        RECT 486.410 2.875 488.790 4.280 ;
        RECT 489.630 2.875 492.470 4.280 ;
        RECT 493.310 2.875 496.150 4.280 ;
        RECT 496.990 2.875 499.830 4.280 ;
        RECT 500.670 2.875 503.050 4.280 ;
        RECT 503.890 2.875 506.730 4.280 ;
        RECT 507.570 2.875 510.410 4.280 ;
        RECT 511.250 2.875 514.090 4.280 ;
        RECT 514.930 2.875 517.310 4.280 ;
        RECT 518.150 2.875 520.990 4.280 ;
        RECT 521.830 2.875 524.670 4.280 ;
        RECT 525.510 2.875 528.350 4.280 ;
        RECT 529.190 2.875 531.570 4.280 ;
        RECT 532.410 2.875 535.250 4.280 ;
        RECT 536.090 2.875 538.930 4.280 ;
        RECT 539.770 2.875 542.610 4.280 ;
        RECT 543.450 2.875 545.830 4.280 ;
        RECT 546.670 2.875 549.510 4.280 ;
        RECT 550.350 2.875 553.190 4.280 ;
        RECT 554.030 2.875 556.870 4.280 ;
        RECT 557.710 2.875 560.090 4.280 ;
        RECT 560.930 2.875 563.770 4.280 ;
        RECT 564.610 2.875 567.450 4.280 ;
        RECT 568.290 2.875 571.130 4.280 ;
        RECT 571.970 2.875 574.350 4.280 ;
        RECT 575.190 2.875 578.030 4.280 ;
        RECT 578.870 2.875 581.710 4.280 ;
        RECT 582.550 2.875 585.390 4.280 ;
        RECT 586.230 2.875 588.610 4.280 ;
        RECT 589.450 2.875 592.290 4.280 ;
        RECT 593.130 2.875 595.970 4.280 ;
        RECT 596.810 2.875 599.650 4.280 ;
        RECT 600.490 2.875 602.870 4.280 ;
        RECT 603.710 2.875 606.550 4.280 ;
        RECT 607.390 2.875 610.230 4.280 ;
        RECT 611.070 2.875 613.910 4.280 ;
        RECT 614.750 2.875 617.130 4.280 ;
        RECT 617.970 2.875 620.810 4.280 ;
        RECT 621.650 2.875 624.490 4.280 ;
        RECT 625.330 2.875 628.170 4.280 ;
        RECT 629.010 2.875 631.390 4.280 ;
        RECT 632.230 2.875 635.070 4.280 ;
        RECT 635.910 2.875 638.750 4.280 ;
        RECT 639.590 2.875 641.970 4.280 ;
        RECT 642.810 2.875 645.650 4.280 ;
        RECT 646.490 2.875 649.330 4.280 ;
        RECT 650.170 2.875 653.010 4.280 ;
        RECT 653.850 2.875 656.230 4.280 ;
        RECT 657.070 2.875 659.910 4.280 ;
        RECT 660.750 2.875 663.590 4.280 ;
        RECT 664.430 2.875 667.270 4.280 ;
        RECT 668.110 2.875 670.490 4.280 ;
        RECT 671.330 2.875 674.170 4.280 ;
        RECT 675.010 2.875 677.850 4.280 ;
        RECT 678.690 2.875 681.530 4.280 ;
        RECT 682.370 2.875 684.750 4.280 ;
        RECT 685.590 2.875 688.430 4.280 ;
        RECT 689.270 2.875 692.110 4.280 ;
        RECT 692.950 2.875 695.790 4.280 ;
        RECT 696.630 2.875 699.010 4.280 ;
        RECT 699.850 2.875 702.690 4.280 ;
        RECT 703.530 2.875 706.370 4.280 ;
        RECT 707.210 2.875 710.050 4.280 ;
        RECT 710.890 2.875 713.270 4.280 ;
        RECT 714.110 2.875 716.950 4.280 ;
        RECT 717.790 2.875 720.630 4.280 ;
        RECT 721.470 2.875 724.310 4.280 ;
        RECT 725.150 2.875 727.530 4.280 ;
        RECT 728.370 2.875 731.210 4.280 ;
        RECT 732.050 2.875 734.890 4.280 ;
        RECT 735.730 2.875 738.570 4.280 ;
        RECT 739.410 2.875 741.790 4.280 ;
        RECT 742.630 2.875 745.470 4.280 ;
        RECT 746.310 2.875 749.150 4.280 ;
        RECT 749.990 2.875 752.830 4.280 ;
        RECT 753.670 2.875 756.050 4.280 ;
        RECT 756.890 2.875 759.730 4.280 ;
        RECT 760.570 2.875 763.410 4.280 ;
        RECT 764.250 2.875 767.090 4.280 ;
        RECT 767.930 2.875 770.310 4.280 ;
        RECT 771.150 2.875 773.990 4.280 ;
        RECT 774.830 2.875 777.670 4.280 ;
        RECT 778.510 2.875 781.350 4.280 ;
        RECT 782.190 2.875 784.570 4.280 ;
        RECT 785.410 2.875 788.250 4.280 ;
        RECT 789.090 2.875 791.930 4.280 ;
        RECT 792.770 2.875 795.610 4.280 ;
        RECT 796.450 2.875 798.830 4.280 ;
        RECT 799.670 2.875 802.510 4.280 ;
        RECT 803.350 2.875 806.190 4.280 ;
        RECT 807.030 2.875 809.410 4.280 ;
        RECT 810.250 2.875 813.090 4.280 ;
        RECT 813.930 2.875 816.770 4.280 ;
        RECT 817.610 2.875 820.450 4.280 ;
        RECT 821.290 2.875 823.670 4.280 ;
        RECT 824.510 2.875 827.350 4.280 ;
        RECT 828.190 2.875 831.030 4.280 ;
        RECT 831.870 2.875 834.710 4.280 ;
        RECT 835.550 2.875 837.930 4.280 ;
        RECT 838.770 2.875 841.610 4.280 ;
        RECT 842.450 2.875 845.290 4.280 ;
        RECT 846.130 2.875 848.970 4.280 ;
        RECT 849.810 2.875 852.190 4.280 ;
        RECT 853.030 2.875 855.870 4.280 ;
        RECT 856.710 2.875 859.550 4.280 ;
        RECT 860.390 2.875 863.230 4.280 ;
        RECT 864.070 2.875 866.450 4.280 ;
        RECT 867.290 2.875 870.130 4.280 ;
        RECT 870.970 2.875 873.810 4.280 ;
        RECT 874.650 2.875 877.490 4.280 ;
        RECT 878.330 2.875 880.710 4.280 ;
        RECT 881.550 2.875 884.390 4.280 ;
        RECT 885.230 2.875 888.070 4.280 ;
        RECT 888.910 2.875 891.750 4.280 ;
        RECT 892.590 2.875 894.970 4.280 ;
        RECT 895.810 2.875 898.650 4.280 ;
        RECT 899.490 2.875 902.330 4.280 ;
        RECT 903.170 2.875 906.010 4.280 ;
        RECT 906.850 2.875 909.230 4.280 ;
        RECT 910.070 2.875 912.910 4.280 ;
        RECT 913.750 2.875 916.590 4.280 ;
        RECT 917.430 2.875 920.270 4.280 ;
        RECT 921.110 2.875 923.490 4.280 ;
        RECT 924.330 2.875 927.170 4.280 ;
        RECT 928.010 2.875 930.850 4.280 ;
        RECT 931.690 2.875 934.530 4.280 ;
        RECT 935.370 2.875 937.750 4.280 ;
        RECT 938.590 2.875 941.430 4.280 ;
        RECT 942.270 2.875 945.110 4.280 ;
        RECT 945.950 2.875 948.790 4.280 ;
        RECT 949.630 2.875 952.010 4.280 ;
        RECT 952.850 2.875 955.690 4.280 ;
        RECT 956.530 2.875 959.370 4.280 ;
        RECT 960.210 2.875 962.590 4.280 ;
        RECT 963.430 2.875 966.270 4.280 ;
        RECT 967.110 2.875 969.950 4.280 ;
        RECT 970.790 2.875 973.630 4.280 ;
        RECT 974.470 2.875 976.850 4.280 ;
        RECT 977.690 2.875 980.530 4.280 ;
        RECT 981.370 2.875 984.210 4.280 ;
        RECT 985.050 2.875 987.890 4.280 ;
        RECT 988.730 2.875 991.110 4.280 ;
        RECT 991.950 2.875 994.790 4.280 ;
        RECT 995.630 2.875 998.470 4.280 ;
        RECT 999.310 2.875 1002.150 4.280 ;
        RECT 1002.990 2.875 1005.370 4.280 ;
        RECT 1006.210 2.875 1009.050 4.280 ;
        RECT 1009.890 2.875 1012.730 4.280 ;
        RECT 1013.570 2.875 1016.410 4.280 ;
        RECT 1017.250 2.875 1019.630 4.280 ;
        RECT 1020.470 2.875 1023.310 4.280 ;
        RECT 1024.150 2.875 1026.990 4.280 ;
        RECT 1027.830 2.875 1030.670 4.280 ;
        RECT 1031.510 2.875 1033.890 4.280 ;
        RECT 1034.730 2.875 1037.570 4.280 ;
        RECT 1038.410 2.875 1041.250 4.280 ;
        RECT 1042.090 2.875 1044.930 4.280 ;
        RECT 1045.770 2.875 1048.150 4.280 ;
        RECT 1048.990 2.875 1051.830 4.280 ;
        RECT 1052.670 2.875 1055.510 4.280 ;
        RECT 1056.350 2.875 1059.190 4.280 ;
        RECT 1060.030 2.875 1062.410 4.280 ;
        RECT 1063.250 2.875 1066.090 4.280 ;
        RECT 1066.930 2.875 1069.770 4.280 ;
        RECT 1070.610 2.875 1073.450 4.280 ;
        RECT 1074.290 2.875 1076.670 4.280 ;
        RECT 1077.510 2.875 1080.350 4.280 ;
        RECT 1081.190 2.875 1084.030 4.280 ;
        RECT 1084.870 2.875 1087.710 4.280 ;
        RECT 1088.550 2.875 1090.930 4.280 ;
        RECT 1091.770 2.875 1094.610 4.280 ;
        RECT 1095.450 2.875 1098.290 4.280 ;
        RECT 1099.130 2.875 1101.970 4.280 ;
        RECT 1102.810 2.875 1105.190 4.280 ;
        RECT 1106.030 2.875 1108.870 4.280 ;
        RECT 1109.710 2.875 1112.550 4.280 ;
        RECT 1113.390 2.875 1116.230 4.280 ;
        RECT 1117.070 2.875 1119.450 4.280 ;
        RECT 1120.290 2.875 1123.130 4.280 ;
        RECT 1123.970 2.875 1126.810 4.280 ;
        RECT 1127.650 2.875 1130.030 4.280 ;
        RECT 1130.870 2.875 1133.710 4.280 ;
        RECT 1134.550 2.875 1137.390 4.280 ;
        RECT 1138.230 2.875 1141.070 4.280 ;
        RECT 1141.910 2.875 1144.290 4.280 ;
        RECT 1145.130 2.875 1147.970 4.280 ;
        RECT 1148.810 2.875 1151.650 4.280 ;
        RECT 1152.490 2.875 1155.330 4.280 ;
        RECT 1156.170 2.875 1158.550 4.280 ;
        RECT 1159.390 2.875 1162.230 4.280 ;
        RECT 1163.070 2.875 1165.910 4.280 ;
        RECT 1166.750 2.875 1169.590 4.280 ;
        RECT 1170.430 2.875 1172.810 4.280 ;
        RECT 1173.650 2.875 1176.490 4.280 ;
        RECT 1177.330 2.875 1180.170 4.280 ;
        RECT 1181.010 2.875 1183.850 4.280 ;
        RECT 1184.690 2.875 1187.070 4.280 ;
        RECT 1187.910 2.875 1190.750 4.280 ;
        RECT 1191.590 2.875 1194.430 4.280 ;
        RECT 1195.270 2.875 1198.110 4.280 ;
        RECT 1198.950 2.875 1201.330 4.280 ;
        RECT 1202.170 2.875 1205.010 4.280 ;
        RECT 1205.850 2.875 1208.690 4.280 ;
        RECT 1209.530 2.875 1212.370 4.280 ;
        RECT 1213.210 2.875 1215.590 4.280 ;
        RECT 1216.430 2.875 1219.270 4.280 ;
        RECT 1220.110 2.875 1222.950 4.280 ;
        RECT 1223.790 2.875 1226.630 4.280 ;
        RECT 1227.470 2.875 1229.850 4.280 ;
        RECT 1230.690 2.875 1233.530 4.280 ;
        RECT 1234.370 2.875 1237.210 4.280 ;
        RECT 1238.050 2.875 1240.890 4.280 ;
        RECT 1241.730 2.875 1244.110 4.280 ;
        RECT 1244.950 2.875 1247.790 4.280 ;
        RECT 1248.630 2.875 1251.470 4.280 ;
        RECT 1252.310 2.875 1255.150 4.280 ;
        RECT 1255.990 2.875 1258.370 4.280 ;
        RECT 1259.210 2.875 1262.050 4.280 ;
        RECT 1262.890 2.875 1265.730 4.280 ;
        RECT 1266.570 2.875 1269.410 4.280 ;
        RECT 1270.250 2.875 1272.630 4.280 ;
        RECT 1273.470 2.875 1276.310 4.280 ;
        RECT 1277.150 2.875 1279.990 4.280 ;
        RECT 1280.830 2.875 1283.210 4.280 ;
        RECT 1284.050 2.875 1286.890 4.280 ;
        RECT 1287.730 2.875 1290.570 4.280 ;
        RECT 1291.410 2.875 1294.250 4.280 ;
        RECT 1295.090 2.875 1297.470 4.280 ;
        RECT 1298.310 2.875 1301.150 4.280 ;
        RECT 1301.990 2.875 1304.830 4.280 ;
        RECT 1305.670 2.875 1308.510 4.280 ;
        RECT 1309.350 2.875 1311.730 4.280 ;
        RECT 1312.570 2.875 1315.410 4.280 ;
        RECT 1316.250 2.875 1319.090 4.280 ;
        RECT 1319.930 2.875 1322.770 4.280 ;
        RECT 1323.610 2.875 1325.990 4.280 ;
        RECT 1326.830 2.875 1329.670 4.280 ;
        RECT 1330.510 2.875 1333.350 4.280 ;
        RECT 1334.190 2.875 1337.030 4.280 ;
        RECT 1337.870 2.875 1340.250 4.280 ;
        RECT 1341.090 2.875 1343.930 4.280 ;
        RECT 1344.770 2.875 1347.610 4.280 ;
        RECT 1348.450 2.875 1351.290 4.280 ;
        RECT 1352.130 2.875 1354.510 4.280 ;
        RECT 1355.350 2.875 1358.190 4.280 ;
        RECT 1359.030 2.875 1361.870 4.280 ;
        RECT 1362.710 2.875 1365.550 4.280 ;
        RECT 1366.390 2.875 1368.770 4.280 ;
        RECT 1369.610 2.875 1372.450 4.280 ;
        RECT 1373.290 2.875 1376.130 4.280 ;
        RECT 1376.970 2.875 1379.810 4.280 ;
        RECT 1380.650 2.875 1383.030 4.280 ;
        RECT 1383.870 2.875 1386.710 4.280 ;
        RECT 1387.550 2.875 1390.390 4.280 ;
        RECT 1391.230 2.875 1394.070 4.280 ;
        RECT 1394.910 2.875 1397.290 4.280 ;
        RECT 1398.130 2.875 1400.970 4.280 ;
        RECT 1401.810 2.875 1404.650 4.280 ;
        RECT 1405.490 2.875 1408.330 4.280 ;
        RECT 1409.170 2.875 1411.550 4.280 ;
        RECT 1412.390 2.875 1415.230 4.280 ;
        RECT 1416.070 2.875 1418.910 4.280 ;
        RECT 1419.750 2.875 1422.590 4.280 ;
        RECT 1423.430 2.875 1425.810 4.280 ;
        RECT 1426.650 2.875 1429.490 4.280 ;
        RECT 1430.330 2.875 1433.170 4.280 ;
        RECT 1434.010 2.875 1436.850 4.280 ;
        RECT 1437.690 2.875 1440.070 4.280 ;
        RECT 1440.910 2.875 1443.750 4.280 ;
        RECT 1444.590 2.875 1447.430 4.280 ;
        RECT 1448.270 2.875 1450.650 4.280 ;
        RECT 1451.490 2.875 1454.330 4.280 ;
        RECT 1455.170 2.875 1458.010 4.280 ;
        RECT 1458.850 2.875 1461.690 4.280 ;
        RECT 1462.530 2.875 1464.910 4.280 ;
        RECT 1465.750 2.875 1468.590 4.280 ;
        RECT 1469.430 2.875 1472.270 4.280 ;
        RECT 1473.110 2.875 1475.950 4.280 ;
        RECT 1476.790 2.875 1479.170 4.280 ;
        RECT 1480.010 2.875 1482.850 4.280 ;
        RECT 1483.690 2.875 1486.530 4.280 ;
        RECT 1487.370 2.875 1490.210 4.280 ;
        RECT 1491.050 2.875 1493.430 4.280 ;
        RECT 1494.270 2.875 1497.110 4.280 ;
        RECT 1497.950 2.875 1500.790 4.280 ;
        RECT 1501.630 2.875 1504.470 4.280 ;
        RECT 1505.310 2.875 1507.690 4.280 ;
        RECT 1508.530 2.875 1511.370 4.280 ;
        RECT 1512.210 2.875 1515.050 4.280 ;
        RECT 1515.890 2.875 1518.730 4.280 ;
        RECT 1519.570 2.875 1521.950 4.280 ;
        RECT 1522.790 2.875 1525.630 4.280 ;
        RECT 1526.470 2.875 1529.310 4.280 ;
        RECT 1530.150 2.875 1532.990 4.280 ;
        RECT 1533.830 2.875 1536.210 4.280 ;
        RECT 1537.050 2.875 1539.890 4.280 ;
        RECT 1540.730 2.875 1543.570 4.280 ;
        RECT 1544.410 2.875 1547.250 4.280 ;
        RECT 1548.090 2.875 1550.470 4.280 ;
        RECT 1551.310 2.875 1554.150 4.280 ;
        RECT 1554.990 2.875 1557.830 4.280 ;
        RECT 1558.670 2.875 1561.510 4.280 ;
        RECT 1562.350 2.875 1564.730 4.280 ;
        RECT 1565.570 2.875 1568.410 4.280 ;
        RECT 1569.250 2.875 1572.090 4.280 ;
        RECT 1572.930 2.875 1575.770 4.280 ;
        RECT 1576.610 2.875 1578.990 4.280 ;
        RECT 1579.830 2.875 1582.670 4.280 ;
        RECT 1583.510 2.875 1586.350 4.280 ;
        RECT 1587.190 2.875 1590.030 4.280 ;
        RECT 1590.870 2.875 1593.250 4.280 ;
        RECT 1594.090 2.875 1596.930 4.280 ;
        RECT 1597.770 2.875 1600.610 4.280 ;
        RECT 1601.450 2.875 1603.830 4.280 ;
        RECT 1604.670 2.875 1607.510 4.280 ;
        RECT 1608.350 2.875 1611.190 4.280 ;
        RECT 1612.030 2.875 1614.870 4.280 ;
        RECT 1615.710 2.875 1618.090 4.280 ;
        RECT 1618.930 2.875 1621.770 4.280 ;
        RECT 1622.610 2.875 1625.450 4.280 ;
        RECT 1626.290 2.875 1629.130 4.280 ;
        RECT 1629.970 2.875 1632.350 4.280 ;
        RECT 1633.190 2.875 1636.030 4.280 ;
        RECT 1636.870 2.875 1639.710 4.280 ;
        RECT 1640.550 2.875 1643.390 4.280 ;
        RECT 1644.230 2.875 1646.610 4.280 ;
        RECT 1647.450 2.875 1650.290 4.280 ;
        RECT 1651.130 2.875 1653.970 4.280 ;
        RECT 1654.810 2.875 1657.650 4.280 ;
        RECT 1658.490 2.875 1660.870 4.280 ;
        RECT 1661.710 2.875 1664.550 4.280 ;
        RECT 1665.390 2.875 1668.230 4.280 ;
        RECT 1669.070 2.875 1671.910 4.280 ;
        RECT 1672.750 2.875 1675.130 4.280 ;
        RECT 1675.970 2.875 1678.810 4.280 ;
        RECT 1679.650 2.875 1682.490 4.280 ;
        RECT 1683.330 2.875 1686.170 4.280 ;
        RECT 1687.010 2.875 1689.390 4.280 ;
        RECT 1690.230 2.875 1693.070 4.280 ;
        RECT 1693.910 2.875 1696.750 4.280 ;
        RECT 1697.590 2.875 1700.430 4.280 ;
        RECT 1701.270 2.875 1703.650 4.280 ;
        RECT 1704.490 2.875 1707.330 4.280 ;
        RECT 1708.170 2.875 1711.010 4.280 ;
        RECT 1711.850 2.875 1714.690 4.280 ;
        RECT 1715.530 2.875 1717.910 4.280 ;
        RECT 1718.750 2.875 1721.590 4.280 ;
        RECT 1722.430 2.875 1725.270 4.280 ;
        RECT 1726.110 2.875 1728.950 4.280 ;
        RECT 1729.790 2.875 1732.170 4.280 ;
        RECT 1733.010 2.875 1735.850 4.280 ;
        RECT 1736.690 2.875 1739.530 4.280 ;
        RECT 1740.370 2.875 1743.210 4.280 ;
        RECT 1744.050 2.875 1746.430 4.280 ;
        RECT 1747.270 2.875 1750.110 4.280 ;
        RECT 1750.950 2.875 1753.790 4.280 ;
      LAYER met3 ;
        RECT 1.445 1764.960 1752.380 1766.465 ;
        RECT 4.400 1763.560 1752.380 1764.960 ;
        RECT 1.445 1758.840 1752.380 1763.560 ;
        RECT 4.400 1757.440 1752.380 1758.840 ;
        RECT 1.445 1752.720 1752.380 1757.440 ;
        RECT 4.400 1751.320 1752.380 1752.720 ;
        RECT 1.445 1747.960 1752.380 1751.320 ;
        RECT 1.445 1746.600 1751.980 1747.960 ;
        RECT 4.400 1746.560 1751.980 1746.600 ;
        RECT 4.400 1745.200 1752.380 1746.560 ;
        RECT 1.445 1740.480 1752.380 1745.200 ;
        RECT 4.400 1739.080 1752.380 1740.480 ;
        RECT 1.445 1734.360 1752.380 1739.080 ;
        RECT 4.400 1732.960 1752.380 1734.360 ;
        RECT 1.445 1728.240 1752.380 1732.960 ;
        RECT 4.400 1726.840 1752.380 1728.240 ;
        RECT 1.445 1722.120 1752.380 1726.840 ;
        RECT 4.400 1720.720 1752.380 1722.120 ;
        RECT 1.445 1716.000 1752.380 1720.720 ;
        RECT 4.400 1714.600 1752.380 1716.000 ;
        RECT 1.445 1709.880 1752.380 1714.600 ;
        RECT 4.400 1708.520 1752.380 1709.880 ;
        RECT 4.400 1708.480 1751.980 1708.520 ;
        RECT 1.445 1707.120 1751.980 1708.480 ;
        RECT 1.445 1703.760 1752.380 1707.120 ;
        RECT 4.400 1702.360 1752.380 1703.760 ;
        RECT 1.445 1697.640 1752.380 1702.360 ;
        RECT 4.400 1696.240 1752.380 1697.640 ;
        RECT 1.445 1691.520 1752.380 1696.240 ;
        RECT 4.400 1690.120 1752.380 1691.520 ;
        RECT 1.445 1685.400 1752.380 1690.120 ;
        RECT 4.400 1684.000 1752.380 1685.400 ;
        RECT 1.445 1679.280 1752.380 1684.000 ;
        RECT 4.400 1677.880 1752.380 1679.280 ;
        RECT 1.445 1673.160 1752.380 1677.880 ;
        RECT 4.400 1671.760 1752.380 1673.160 ;
        RECT 1.445 1669.080 1752.380 1671.760 ;
        RECT 1.445 1667.680 1751.980 1669.080 ;
        RECT 1.445 1667.040 1752.380 1667.680 ;
        RECT 4.400 1665.640 1752.380 1667.040 ;
        RECT 1.445 1660.920 1752.380 1665.640 ;
        RECT 4.400 1659.520 1752.380 1660.920 ;
        RECT 1.445 1654.800 1752.380 1659.520 ;
        RECT 4.400 1653.400 1752.380 1654.800 ;
        RECT 1.445 1648.680 1752.380 1653.400 ;
        RECT 4.400 1647.280 1752.380 1648.680 ;
        RECT 1.445 1642.560 1752.380 1647.280 ;
        RECT 4.400 1641.160 1752.380 1642.560 ;
        RECT 1.445 1636.440 1752.380 1641.160 ;
        RECT 4.400 1635.040 1752.380 1636.440 ;
        RECT 1.445 1630.320 1752.380 1635.040 ;
        RECT 4.400 1629.640 1752.380 1630.320 ;
        RECT 4.400 1628.920 1751.980 1629.640 ;
        RECT 1.445 1628.240 1751.980 1628.920 ;
        RECT 1.445 1624.200 1752.380 1628.240 ;
        RECT 4.400 1622.800 1752.380 1624.200 ;
        RECT 1.445 1618.080 1752.380 1622.800 ;
        RECT 4.400 1616.680 1752.380 1618.080 ;
        RECT 1.445 1611.960 1752.380 1616.680 ;
        RECT 4.400 1610.560 1752.380 1611.960 ;
        RECT 1.445 1606.520 1752.380 1610.560 ;
        RECT 4.400 1605.120 1752.380 1606.520 ;
        RECT 1.445 1600.400 1752.380 1605.120 ;
        RECT 4.400 1599.000 1752.380 1600.400 ;
        RECT 1.445 1594.280 1752.380 1599.000 ;
        RECT 4.400 1592.880 1752.380 1594.280 ;
        RECT 1.445 1590.880 1752.380 1592.880 ;
        RECT 1.445 1589.480 1751.980 1590.880 ;
        RECT 1.445 1588.160 1752.380 1589.480 ;
        RECT 4.400 1586.760 1752.380 1588.160 ;
        RECT 1.445 1582.040 1752.380 1586.760 ;
        RECT 4.400 1580.640 1752.380 1582.040 ;
        RECT 1.445 1575.920 1752.380 1580.640 ;
        RECT 4.400 1574.520 1752.380 1575.920 ;
        RECT 1.445 1569.800 1752.380 1574.520 ;
        RECT 4.400 1568.400 1752.380 1569.800 ;
        RECT 1.445 1563.680 1752.380 1568.400 ;
        RECT 4.400 1562.280 1752.380 1563.680 ;
        RECT 1.445 1557.560 1752.380 1562.280 ;
        RECT 4.400 1556.160 1752.380 1557.560 ;
        RECT 1.445 1551.440 1752.380 1556.160 ;
        RECT 4.400 1550.040 1751.980 1551.440 ;
        RECT 1.445 1545.320 1752.380 1550.040 ;
        RECT 4.400 1543.920 1752.380 1545.320 ;
        RECT 1.445 1539.200 1752.380 1543.920 ;
        RECT 4.400 1537.800 1752.380 1539.200 ;
        RECT 1.445 1533.080 1752.380 1537.800 ;
        RECT 4.400 1531.680 1752.380 1533.080 ;
        RECT 1.445 1526.960 1752.380 1531.680 ;
        RECT 4.400 1525.560 1752.380 1526.960 ;
        RECT 1.445 1520.840 1752.380 1525.560 ;
        RECT 4.400 1519.440 1752.380 1520.840 ;
        RECT 1.445 1514.720 1752.380 1519.440 ;
        RECT 4.400 1513.320 1752.380 1514.720 ;
        RECT 1.445 1512.000 1752.380 1513.320 ;
        RECT 1.445 1510.600 1751.980 1512.000 ;
        RECT 1.445 1508.600 1752.380 1510.600 ;
        RECT 4.400 1507.200 1752.380 1508.600 ;
        RECT 1.445 1502.480 1752.380 1507.200 ;
        RECT 4.400 1501.080 1752.380 1502.480 ;
        RECT 1.445 1496.360 1752.380 1501.080 ;
        RECT 4.400 1494.960 1752.380 1496.360 ;
        RECT 1.445 1490.240 1752.380 1494.960 ;
        RECT 4.400 1488.840 1752.380 1490.240 ;
        RECT 1.445 1484.120 1752.380 1488.840 ;
        RECT 4.400 1482.720 1752.380 1484.120 ;
        RECT 1.445 1478.000 1752.380 1482.720 ;
        RECT 4.400 1476.600 1752.380 1478.000 ;
        RECT 1.445 1472.560 1752.380 1476.600 ;
        RECT 1.445 1471.880 1751.980 1472.560 ;
        RECT 4.400 1471.160 1751.980 1471.880 ;
        RECT 4.400 1470.480 1752.380 1471.160 ;
        RECT 1.445 1465.760 1752.380 1470.480 ;
        RECT 4.400 1464.360 1752.380 1465.760 ;
        RECT 1.445 1459.640 1752.380 1464.360 ;
        RECT 4.400 1458.240 1752.380 1459.640 ;
        RECT 1.445 1453.520 1752.380 1458.240 ;
        RECT 4.400 1452.120 1752.380 1453.520 ;
        RECT 1.445 1448.080 1752.380 1452.120 ;
        RECT 4.400 1446.680 1752.380 1448.080 ;
        RECT 1.445 1441.960 1752.380 1446.680 ;
        RECT 4.400 1440.560 1752.380 1441.960 ;
        RECT 1.445 1435.840 1752.380 1440.560 ;
        RECT 4.400 1434.440 1752.380 1435.840 ;
        RECT 1.445 1433.800 1752.380 1434.440 ;
        RECT 1.445 1432.400 1751.980 1433.800 ;
        RECT 1.445 1429.720 1752.380 1432.400 ;
        RECT 4.400 1428.320 1752.380 1429.720 ;
        RECT 1.445 1423.600 1752.380 1428.320 ;
        RECT 4.400 1422.200 1752.380 1423.600 ;
        RECT 1.445 1417.480 1752.380 1422.200 ;
        RECT 4.400 1416.080 1752.380 1417.480 ;
        RECT 1.445 1411.360 1752.380 1416.080 ;
        RECT 4.400 1409.960 1752.380 1411.360 ;
        RECT 1.445 1405.240 1752.380 1409.960 ;
        RECT 4.400 1403.840 1752.380 1405.240 ;
        RECT 1.445 1399.120 1752.380 1403.840 ;
        RECT 4.400 1397.720 1752.380 1399.120 ;
        RECT 1.445 1394.360 1752.380 1397.720 ;
        RECT 1.445 1393.000 1751.980 1394.360 ;
        RECT 4.400 1392.960 1751.980 1393.000 ;
        RECT 4.400 1391.600 1752.380 1392.960 ;
        RECT 1.445 1386.880 1752.380 1391.600 ;
        RECT 4.400 1385.480 1752.380 1386.880 ;
        RECT 1.445 1380.760 1752.380 1385.480 ;
        RECT 4.400 1379.360 1752.380 1380.760 ;
        RECT 1.445 1374.640 1752.380 1379.360 ;
        RECT 4.400 1373.240 1752.380 1374.640 ;
        RECT 1.445 1368.520 1752.380 1373.240 ;
        RECT 4.400 1367.120 1752.380 1368.520 ;
        RECT 1.445 1362.400 1752.380 1367.120 ;
        RECT 4.400 1361.000 1752.380 1362.400 ;
        RECT 1.445 1356.280 1752.380 1361.000 ;
        RECT 4.400 1354.920 1752.380 1356.280 ;
        RECT 4.400 1354.880 1751.980 1354.920 ;
        RECT 1.445 1353.520 1751.980 1354.880 ;
        RECT 1.445 1350.160 1752.380 1353.520 ;
        RECT 4.400 1348.760 1752.380 1350.160 ;
        RECT 1.445 1344.040 1752.380 1348.760 ;
        RECT 4.400 1342.640 1752.380 1344.040 ;
        RECT 1.445 1337.920 1752.380 1342.640 ;
        RECT 4.400 1336.520 1752.380 1337.920 ;
        RECT 1.445 1331.800 1752.380 1336.520 ;
        RECT 4.400 1330.400 1752.380 1331.800 ;
        RECT 1.445 1325.680 1752.380 1330.400 ;
        RECT 4.400 1324.280 1752.380 1325.680 ;
        RECT 1.445 1319.560 1752.380 1324.280 ;
        RECT 4.400 1318.160 1752.380 1319.560 ;
        RECT 1.445 1315.480 1752.380 1318.160 ;
        RECT 1.445 1314.080 1751.980 1315.480 ;
        RECT 1.445 1313.440 1752.380 1314.080 ;
        RECT 4.400 1312.040 1752.380 1313.440 ;
        RECT 1.445 1307.320 1752.380 1312.040 ;
        RECT 4.400 1305.920 1752.380 1307.320 ;
        RECT 1.445 1301.200 1752.380 1305.920 ;
        RECT 4.400 1299.800 1752.380 1301.200 ;
        RECT 1.445 1295.080 1752.380 1299.800 ;
        RECT 4.400 1293.680 1752.380 1295.080 ;
        RECT 1.445 1288.960 1752.380 1293.680 ;
        RECT 4.400 1287.560 1752.380 1288.960 ;
        RECT 1.445 1283.520 1752.380 1287.560 ;
        RECT 4.400 1282.120 1752.380 1283.520 ;
        RECT 1.445 1277.400 1752.380 1282.120 ;
        RECT 4.400 1276.720 1752.380 1277.400 ;
        RECT 4.400 1276.000 1751.980 1276.720 ;
        RECT 1.445 1275.320 1751.980 1276.000 ;
        RECT 1.445 1271.280 1752.380 1275.320 ;
        RECT 4.400 1269.880 1752.380 1271.280 ;
        RECT 1.445 1265.160 1752.380 1269.880 ;
        RECT 4.400 1263.760 1752.380 1265.160 ;
        RECT 1.445 1259.040 1752.380 1263.760 ;
        RECT 4.400 1257.640 1752.380 1259.040 ;
        RECT 1.445 1252.920 1752.380 1257.640 ;
        RECT 4.400 1251.520 1752.380 1252.920 ;
        RECT 1.445 1246.800 1752.380 1251.520 ;
        RECT 4.400 1245.400 1752.380 1246.800 ;
        RECT 1.445 1240.680 1752.380 1245.400 ;
        RECT 4.400 1239.280 1752.380 1240.680 ;
        RECT 1.445 1237.280 1752.380 1239.280 ;
        RECT 1.445 1235.880 1751.980 1237.280 ;
        RECT 1.445 1234.560 1752.380 1235.880 ;
        RECT 4.400 1233.160 1752.380 1234.560 ;
        RECT 1.445 1228.440 1752.380 1233.160 ;
        RECT 4.400 1227.040 1752.380 1228.440 ;
        RECT 1.445 1222.320 1752.380 1227.040 ;
        RECT 4.400 1220.920 1752.380 1222.320 ;
        RECT 1.445 1216.200 1752.380 1220.920 ;
        RECT 4.400 1214.800 1752.380 1216.200 ;
        RECT 1.445 1210.080 1752.380 1214.800 ;
        RECT 4.400 1208.680 1752.380 1210.080 ;
        RECT 1.445 1203.960 1752.380 1208.680 ;
        RECT 4.400 1202.560 1752.380 1203.960 ;
        RECT 1.445 1197.840 1752.380 1202.560 ;
        RECT 4.400 1196.440 1751.980 1197.840 ;
        RECT 1.445 1191.720 1752.380 1196.440 ;
        RECT 4.400 1190.320 1752.380 1191.720 ;
        RECT 1.445 1185.600 1752.380 1190.320 ;
        RECT 4.400 1184.200 1752.380 1185.600 ;
        RECT 1.445 1179.480 1752.380 1184.200 ;
        RECT 4.400 1178.080 1752.380 1179.480 ;
        RECT 1.445 1173.360 1752.380 1178.080 ;
        RECT 4.400 1171.960 1752.380 1173.360 ;
        RECT 1.445 1167.240 1752.380 1171.960 ;
        RECT 4.400 1165.840 1752.380 1167.240 ;
        RECT 1.445 1161.120 1752.380 1165.840 ;
        RECT 4.400 1159.720 1752.380 1161.120 ;
        RECT 1.445 1158.400 1752.380 1159.720 ;
        RECT 1.445 1157.000 1751.980 1158.400 ;
        RECT 1.445 1155.000 1752.380 1157.000 ;
        RECT 4.400 1153.600 1752.380 1155.000 ;
        RECT 1.445 1148.880 1752.380 1153.600 ;
        RECT 4.400 1147.480 1752.380 1148.880 ;
        RECT 1.445 1142.760 1752.380 1147.480 ;
        RECT 4.400 1141.360 1752.380 1142.760 ;
        RECT 1.445 1136.640 1752.380 1141.360 ;
        RECT 4.400 1135.240 1752.380 1136.640 ;
        RECT 1.445 1130.520 1752.380 1135.240 ;
        RECT 4.400 1129.120 1752.380 1130.520 ;
        RECT 1.445 1125.080 1752.380 1129.120 ;
        RECT 4.400 1123.680 1752.380 1125.080 ;
        RECT 1.445 1119.640 1752.380 1123.680 ;
        RECT 1.445 1118.960 1751.980 1119.640 ;
        RECT 4.400 1118.240 1751.980 1118.960 ;
        RECT 4.400 1117.560 1752.380 1118.240 ;
        RECT 1.445 1112.840 1752.380 1117.560 ;
        RECT 4.400 1111.440 1752.380 1112.840 ;
        RECT 1.445 1106.720 1752.380 1111.440 ;
        RECT 4.400 1105.320 1752.380 1106.720 ;
        RECT 1.445 1100.600 1752.380 1105.320 ;
        RECT 4.400 1099.200 1752.380 1100.600 ;
        RECT 1.445 1094.480 1752.380 1099.200 ;
        RECT 4.400 1093.080 1752.380 1094.480 ;
        RECT 1.445 1088.360 1752.380 1093.080 ;
        RECT 4.400 1086.960 1752.380 1088.360 ;
        RECT 1.445 1082.240 1752.380 1086.960 ;
        RECT 4.400 1080.840 1752.380 1082.240 ;
        RECT 1.445 1080.200 1752.380 1080.840 ;
        RECT 1.445 1078.800 1751.980 1080.200 ;
        RECT 1.445 1076.120 1752.380 1078.800 ;
        RECT 4.400 1074.720 1752.380 1076.120 ;
        RECT 1.445 1070.000 1752.380 1074.720 ;
        RECT 4.400 1068.600 1752.380 1070.000 ;
        RECT 1.445 1063.880 1752.380 1068.600 ;
        RECT 4.400 1062.480 1752.380 1063.880 ;
        RECT 1.445 1057.760 1752.380 1062.480 ;
        RECT 4.400 1056.360 1752.380 1057.760 ;
        RECT 1.445 1051.640 1752.380 1056.360 ;
        RECT 4.400 1050.240 1752.380 1051.640 ;
        RECT 1.445 1045.520 1752.380 1050.240 ;
        RECT 4.400 1044.120 1752.380 1045.520 ;
        RECT 1.445 1040.760 1752.380 1044.120 ;
        RECT 1.445 1039.400 1751.980 1040.760 ;
        RECT 4.400 1039.360 1751.980 1039.400 ;
        RECT 4.400 1038.000 1752.380 1039.360 ;
        RECT 1.445 1033.280 1752.380 1038.000 ;
        RECT 4.400 1031.880 1752.380 1033.280 ;
        RECT 1.445 1027.160 1752.380 1031.880 ;
        RECT 4.400 1025.760 1752.380 1027.160 ;
        RECT 1.445 1021.040 1752.380 1025.760 ;
        RECT 4.400 1019.640 1752.380 1021.040 ;
        RECT 1.445 1014.920 1752.380 1019.640 ;
        RECT 4.400 1013.520 1752.380 1014.920 ;
        RECT 1.445 1008.800 1752.380 1013.520 ;
        RECT 4.400 1007.400 1752.380 1008.800 ;
        RECT 1.445 1002.680 1752.380 1007.400 ;
        RECT 4.400 1001.320 1752.380 1002.680 ;
        RECT 4.400 1001.280 1751.980 1001.320 ;
        RECT 1.445 999.920 1751.980 1001.280 ;
        RECT 1.445 996.560 1752.380 999.920 ;
        RECT 4.400 995.160 1752.380 996.560 ;
        RECT 1.445 990.440 1752.380 995.160 ;
        RECT 4.400 989.040 1752.380 990.440 ;
        RECT 1.445 984.320 1752.380 989.040 ;
        RECT 4.400 982.920 1752.380 984.320 ;
        RECT 1.445 978.200 1752.380 982.920 ;
        RECT 4.400 976.800 1752.380 978.200 ;
        RECT 1.445 972.080 1752.380 976.800 ;
        RECT 4.400 970.680 1752.380 972.080 ;
        RECT 1.445 966.640 1752.380 970.680 ;
        RECT 4.400 965.240 1752.380 966.640 ;
        RECT 1.445 962.560 1752.380 965.240 ;
        RECT 1.445 961.160 1751.980 962.560 ;
        RECT 1.445 960.520 1752.380 961.160 ;
        RECT 4.400 959.120 1752.380 960.520 ;
        RECT 1.445 954.400 1752.380 959.120 ;
        RECT 4.400 953.000 1752.380 954.400 ;
        RECT 1.445 948.280 1752.380 953.000 ;
        RECT 4.400 946.880 1752.380 948.280 ;
        RECT 1.445 942.160 1752.380 946.880 ;
        RECT 4.400 940.760 1752.380 942.160 ;
        RECT 1.445 936.040 1752.380 940.760 ;
        RECT 4.400 934.640 1752.380 936.040 ;
        RECT 1.445 929.920 1752.380 934.640 ;
        RECT 4.400 928.520 1752.380 929.920 ;
        RECT 1.445 923.800 1752.380 928.520 ;
        RECT 4.400 923.120 1752.380 923.800 ;
        RECT 4.400 922.400 1751.980 923.120 ;
        RECT 1.445 921.720 1751.980 922.400 ;
        RECT 1.445 917.680 1752.380 921.720 ;
        RECT 4.400 916.280 1752.380 917.680 ;
        RECT 1.445 911.560 1752.380 916.280 ;
        RECT 4.400 910.160 1752.380 911.560 ;
        RECT 1.445 905.440 1752.380 910.160 ;
        RECT 4.400 904.040 1752.380 905.440 ;
        RECT 1.445 899.320 1752.380 904.040 ;
        RECT 4.400 897.920 1752.380 899.320 ;
        RECT 1.445 893.200 1752.380 897.920 ;
        RECT 4.400 891.800 1752.380 893.200 ;
        RECT 1.445 887.080 1752.380 891.800 ;
        RECT 4.400 885.680 1752.380 887.080 ;
        RECT 1.445 883.680 1752.380 885.680 ;
        RECT 1.445 882.280 1751.980 883.680 ;
        RECT 1.445 880.960 1752.380 882.280 ;
        RECT 4.400 879.560 1752.380 880.960 ;
        RECT 1.445 874.840 1752.380 879.560 ;
        RECT 4.400 873.440 1752.380 874.840 ;
        RECT 1.445 868.720 1752.380 873.440 ;
        RECT 4.400 867.320 1752.380 868.720 ;
        RECT 1.445 862.600 1752.380 867.320 ;
        RECT 4.400 861.200 1752.380 862.600 ;
        RECT 1.445 856.480 1752.380 861.200 ;
        RECT 4.400 855.080 1752.380 856.480 ;
        RECT 1.445 850.360 1752.380 855.080 ;
        RECT 4.400 848.960 1752.380 850.360 ;
        RECT 1.445 844.240 1752.380 848.960 ;
        RECT 4.400 842.840 1751.980 844.240 ;
        RECT 1.445 838.120 1752.380 842.840 ;
        RECT 4.400 836.720 1752.380 838.120 ;
        RECT 1.445 832.000 1752.380 836.720 ;
        RECT 4.400 830.600 1752.380 832.000 ;
        RECT 1.445 825.880 1752.380 830.600 ;
        RECT 4.400 824.480 1752.380 825.880 ;
        RECT 1.445 819.760 1752.380 824.480 ;
        RECT 4.400 818.360 1752.380 819.760 ;
        RECT 1.445 813.640 1752.380 818.360 ;
        RECT 4.400 812.240 1752.380 813.640 ;
        RECT 1.445 807.520 1752.380 812.240 ;
        RECT 4.400 806.120 1752.380 807.520 ;
        RECT 1.445 805.480 1752.380 806.120 ;
        RECT 1.445 804.080 1751.980 805.480 ;
        RECT 1.445 802.080 1752.380 804.080 ;
        RECT 4.400 800.680 1752.380 802.080 ;
        RECT 1.445 795.960 1752.380 800.680 ;
        RECT 4.400 794.560 1752.380 795.960 ;
        RECT 1.445 789.840 1752.380 794.560 ;
        RECT 4.400 788.440 1752.380 789.840 ;
        RECT 1.445 783.720 1752.380 788.440 ;
        RECT 4.400 782.320 1752.380 783.720 ;
        RECT 1.445 777.600 1752.380 782.320 ;
        RECT 4.400 776.200 1752.380 777.600 ;
        RECT 1.445 771.480 1752.380 776.200 ;
        RECT 4.400 770.080 1752.380 771.480 ;
        RECT 1.445 766.040 1752.380 770.080 ;
        RECT 1.445 765.360 1751.980 766.040 ;
        RECT 4.400 764.640 1751.980 765.360 ;
        RECT 4.400 763.960 1752.380 764.640 ;
        RECT 1.445 759.240 1752.380 763.960 ;
        RECT 4.400 757.840 1752.380 759.240 ;
        RECT 1.445 753.120 1752.380 757.840 ;
        RECT 4.400 751.720 1752.380 753.120 ;
        RECT 1.445 747.000 1752.380 751.720 ;
        RECT 4.400 745.600 1752.380 747.000 ;
        RECT 1.445 740.880 1752.380 745.600 ;
        RECT 4.400 739.480 1752.380 740.880 ;
        RECT 1.445 734.760 1752.380 739.480 ;
        RECT 4.400 733.360 1752.380 734.760 ;
        RECT 1.445 728.640 1752.380 733.360 ;
        RECT 4.400 727.240 1752.380 728.640 ;
        RECT 1.445 726.600 1752.380 727.240 ;
        RECT 1.445 725.200 1751.980 726.600 ;
        RECT 1.445 722.520 1752.380 725.200 ;
        RECT 4.400 721.120 1752.380 722.520 ;
        RECT 1.445 716.400 1752.380 721.120 ;
        RECT 4.400 715.000 1752.380 716.400 ;
        RECT 1.445 710.280 1752.380 715.000 ;
        RECT 4.400 708.880 1752.380 710.280 ;
        RECT 1.445 704.160 1752.380 708.880 ;
        RECT 4.400 702.760 1752.380 704.160 ;
        RECT 1.445 698.040 1752.380 702.760 ;
        RECT 4.400 696.640 1752.380 698.040 ;
        RECT 1.445 691.920 1752.380 696.640 ;
        RECT 4.400 690.520 1752.380 691.920 ;
        RECT 1.445 687.160 1752.380 690.520 ;
        RECT 1.445 685.800 1751.980 687.160 ;
        RECT 4.400 685.760 1751.980 685.800 ;
        RECT 4.400 684.400 1752.380 685.760 ;
        RECT 1.445 679.680 1752.380 684.400 ;
        RECT 4.400 678.280 1752.380 679.680 ;
        RECT 1.445 673.560 1752.380 678.280 ;
        RECT 4.400 672.160 1752.380 673.560 ;
        RECT 1.445 667.440 1752.380 672.160 ;
        RECT 4.400 666.040 1752.380 667.440 ;
        RECT 1.445 661.320 1752.380 666.040 ;
        RECT 4.400 659.920 1752.380 661.320 ;
        RECT 1.445 655.200 1752.380 659.920 ;
        RECT 4.400 653.800 1752.380 655.200 ;
        RECT 1.445 649.080 1752.380 653.800 ;
        RECT 4.400 648.400 1752.380 649.080 ;
        RECT 4.400 647.680 1751.980 648.400 ;
        RECT 1.445 647.000 1751.980 647.680 ;
        RECT 1.445 643.640 1752.380 647.000 ;
        RECT 4.400 642.240 1752.380 643.640 ;
        RECT 1.445 637.520 1752.380 642.240 ;
        RECT 4.400 636.120 1752.380 637.520 ;
        RECT 1.445 631.400 1752.380 636.120 ;
        RECT 4.400 630.000 1752.380 631.400 ;
        RECT 1.445 625.280 1752.380 630.000 ;
        RECT 4.400 623.880 1752.380 625.280 ;
        RECT 1.445 619.160 1752.380 623.880 ;
        RECT 4.400 617.760 1752.380 619.160 ;
        RECT 1.445 613.040 1752.380 617.760 ;
        RECT 4.400 611.640 1752.380 613.040 ;
        RECT 1.445 608.960 1752.380 611.640 ;
        RECT 1.445 607.560 1751.980 608.960 ;
        RECT 1.445 606.920 1752.380 607.560 ;
        RECT 4.400 605.520 1752.380 606.920 ;
        RECT 1.445 600.800 1752.380 605.520 ;
        RECT 4.400 599.400 1752.380 600.800 ;
        RECT 1.445 594.680 1752.380 599.400 ;
        RECT 4.400 593.280 1752.380 594.680 ;
        RECT 1.445 588.560 1752.380 593.280 ;
        RECT 4.400 587.160 1752.380 588.560 ;
        RECT 1.445 582.440 1752.380 587.160 ;
        RECT 4.400 581.040 1752.380 582.440 ;
        RECT 1.445 576.320 1752.380 581.040 ;
        RECT 4.400 574.920 1752.380 576.320 ;
        RECT 1.445 570.200 1752.380 574.920 ;
        RECT 4.400 569.520 1752.380 570.200 ;
        RECT 4.400 568.800 1751.980 569.520 ;
        RECT 1.445 568.120 1751.980 568.800 ;
        RECT 1.445 564.080 1752.380 568.120 ;
        RECT 4.400 562.680 1752.380 564.080 ;
        RECT 1.445 557.960 1752.380 562.680 ;
        RECT 4.400 556.560 1752.380 557.960 ;
        RECT 1.445 551.840 1752.380 556.560 ;
        RECT 4.400 550.440 1752.380 551.840 ;
        RECT 1.445 545.720 1752.380 550.440 ;
        RECT 4.400 544.320 1752.380 545.720 ;
        RECT 1.445 539.600 1752.380 544.320 ;
        RECT 4.400 538.200 1752.380 539.600 ;
        RECT 1.445 533.480 1752.380 538.200 ;
        RECT 4.400 532.080 1752.380 533.480 ;
        RECT 1.445 530.080 1752.380 532.080 ;
        RECT 1.445 528.680 1751.980 530.080 ;
        RECT 1.445 527.360 1752.380 528.680 ;
        RECT 4.400 525.960 1752.380 527.360 ;
        RECT 1.445 521.240 1752.380 525.960 ;
        RECT 4.400 519.840 1752.380 521.240 ;
        RECT 1.445 515.120 1752.380 519.840 ;
        RECT 4.400 513.720 1752.380 515.120 ;
        RECT 1.445 509.000 1752.380 513.720 ;
        RECT 4.400 507.600 1752.380 509.000 ;
        RECT 1.445 502.880 1752.380 507.600 ;
        RECT 4.400 501.480 1752.380 502.880 ;
        RECT 1.445 496.760 1752.380 501.480 ;
        RECT 4.400 495.360 1752.380 496.760 ;
        RECT 1.445 491.320 1752.380 495.360 ;
        RECT 1.445 490.640 1751.980 491.320 ;
        RECT 4.400 489.920 1751.980 490.640 ;
        RECT 4.400 489.240 1752.380 489.920 ;
        RECT 1.445 485.200 1752.380 489.240 ;
        RECT 4.400 483.800 1752.380 485.200 ;
        RECT 1.445 479.080 1752.380 483.800 ;
        RECT 4.400 477.680 1752.380 479.080 ;
        RECT 1.445 472.960 1752.380 477.680 ;
        RECT 4.400 471.560 1752.380 472.960 ;
        RECT 1.445 466.840 1752.380 471.560 ;
        RECT 4.400 465.440 1752.380 466.840 ;
        RECT 1.445 460.720 1752.380 465.440 ;
        RECT 4.400 459.320 1752.380 460.720 ;
        RECT 1.445 454.600 1752.380 459.320 ;
        RECT 4.400 453.200 1752.380 454.600 ;
        RECT 1.445 451.880 1752.380 453.200 ;
        RECT 1.445 450.480 1751.980 451.880 ;
        RECT 1.445 448.480 1752.380 450.480 ;
        RECT 4.400 447.080 1752.380 448.480 ;
        RECT 1.445 442.360 1752.380 447.080 ;
        RECT 4.400 440.960 1752.380 442.360 ;
        RECT 1.445 436.240 1752.380 440.960 ;
        RECT 4.400 434.840 1752.380 436.240 ;
        RECT 1.445 430.120 1752.380 434.840 ;
        RECT 4.400 428.720 1752.380 430.120 ;
        RECT 1.445 424.000 1752.380 428.720 ;
        RECT 4.400 422.600 1752.380 424.000 ;
        RECT 1.445 417.880 1752.380 422.600 ;
        RECT 4.400 416.480 1752.380 417.880 ;
        RECT 1.445 412.440 1752.380 416.480 ;
        RECT 1.445 411.760 1751.980 412.440 ;
        RECT 4.400 411.040 1751.980 411.760 ;
        RECT 4.400 410.360 1752.380 411.040 ;
        RECT 1.445 405.640 1752.380 410.360 ;
        RECT 4.400 404.240 1752.380 405.640 ;
        RECT 1.445 399.520 1752.380 404.240 ;
        RECT 4.400 398.120 1752.380 399.520 ;
        RECT 1.445 393.400 1752.380 398.120 ;
        RECT 4.400 392.000 1752.380 393.400 ;
        RECT 1.445 387.280 1752.380 392.000 ;
        RECT 4.400 385.880 1752.380 387.280 ;
        RECT 1.445 381.160 1752.380 385.880 ;
        RECT 4.400 379.760 1752.380 381.160 ;
        RECT 1.445 375.040 1752.380 379.760 ;
        RECT 4.400 373.640 1752.380 375.040 ;
        RECT 1.445 373.000 1752.380 373.640 ;
        RECT 1.445 371.600 1751.980 373.000 ;
        RECT 1.445 368.920 1752.380 371.600 ;
        RECT 4.400 367.520 1752.380 368.920 ;
        RECT 1.445 362.800 1752.380 367.520 ;
        RECT 4.400 361.400 1752.380 362.800 ;
        RECT 1.445 356.680 1752.380 361.400 ;
        RECT 4.400 355.280 1752.380 356.680 ;
        RECT 1.445 350.560 1752.380 355.280 ;
        RECT 4.400 349.160 1752.380 350.560 ;
        RECT 1.445 344.440 1752.380 349.160 ;
        RECT 4.400 343.040 1752.380 344.440 ;
        RECT 1.445 338.320 1752.380 343.040 ;
        RECT 4.400 336.920 1752.380 338.320 ;
        RECT 1.445 334.240 1752.380 336.920 ;
        RECT 1.445 332.840 1751.980 334.240 ;
        RECT 1.445 332.200 1752.380 332.840 ;
        RECT 4.400 330.800 1752.380 332.200 ;
        RECT 1.445 326.080 1752.380 330.800 ;
        RECT 4.400 324.680 1752.380 326.080 ;
        RECT 1.445 320.640 1752.380 324.680 ;
        RECT 4.400 319.240 1752.380 320.640 ;
        RECT 1.445 314.520 1752.380 319.240 ;
        RECT 4.400 313.120 1752.380 314.520 ;
        RECT 1.445 308.400 1752.380 313.120 ;
        RECT 4.400 307.000 1752.380 308.400 ;
        RECT 1.445 302.280 1752.380 307.000 ;
        RECT 4.400 300.880 1752.380 302.280 ;
        RECT 1.445 296.160 1752.380 300.880 ;
        RECT 4.400 294.800 1752.380 296.160 ;
        RECT 4.400 294.760 1751.980 294.800 ;
        RECT 1.445 293.400 1751.980 294.760 ;
        RECT 1.445 290.040 1752.380 293.400 ;
        RECT 4.400 288.640 1752.380 290.040 ;
        RECT 1.445 283.920 1752.380 288.640 ;
        RECT 4.400 282.520 1752.380 283.920 ;
        RECT 1.445 277.800 1752.380 282.520 ;
        RECT 4.400 276.400 1752.380 277.800 ;
        RECT 1.445 271.680 1752.380 276.400 ;
        RECT 4.400 270.280 1752.380 271.680 ;
        RECT 1.445 265.560 1752.380 270.280 ;
        RECT 4.400 264.160 1752.380 265.560 ;
        RECT 1.445 259.440 1752.380 264.160 ;
        RECT 4.400 258.040 1752.380 259.440 ;
        RECT 1.445 255.360 1752.380 258.040 ;
        RECT 1.445 253.960 1751.980 255.360 ;
        RECT 1.445 253.320 1752.380 253.960 ;
        RECT 4.400 251.920 1752.380 253.320 ;
        RECT 1.445 247.200 1752.380 251.920 ;
        RECT 4.400 245.800 1752.380 247.200 ;
        RECT 1.445 241.080 1752.380 245.800 ;
        RECT 4.400 239.680 1752.380 241.080 ;
        RECT 1.445 234.960 1752.380 239.680 ;
        RECT 4.400 233.560 1752.380 234.960 ;
        RECT 1.445 228.840 1752.380 233.560 ;
        RECT 4.400 227.440 1752.380 228.840 ;
        RECT 1.445 222.720 1752.380 227.440 ;
        RECT 4.400 221.320 1752.380 222.720 ;
        RECT 1.445 216.600 1752.380 221.320 ;
        RECT 4.400 215.920 1752.380 216.600 ;
        RECT 4.400 215.200 1751.980 215.920 ;
        RECT 1.445 214.520 1751.980 215.200 ;
        RECT 1.445 210.480 1752.380 214.520 ;
        RECT 4.400 209.080 1752.380 210.480 ;
        RECT 1.445 204.360 1752.380 209.080 ;
        RECT 4.400 202.960 1752.380 204.360 ;
        RECT 1.445 198.240 1752.380 202.960 ;
        RECT 4.400 196.840 1752.380 198.240 ;
        RECT 1.445 192.120 1752.380 196.840 ;
        RECT 4.400 190.720 1752.380 192.120 ;
        RECT 1.445 186.000 1752.380 190.720 ;
        RECT 4.400 184.600 1752.380 186.000 ;
        RECT 1.445 179.880 1752.380 184.600 ;
        RECT 4.400 178.480 1752.380 179.880 ;
        RECT 1.445 177.160 1752.380 178.480 ;
        RECT 1.445 175.760 1751.980 177.160 ;
        RECT 1.445 173.760 1752.380 175.760 ;
        RECT 4.400 172.360 1752.380 173.760 ;
        RECT 1.445 167.640 1752.380 172.360 ;
        RECT 4.400 166.240 1752.380 167.640 ;
        RECT 1.445 162.200 1752.380 166.240 ;
        RECT 4.400 160.800 1752.380 162.200 ;
        RECT 1.445 156.080 1752.380 160.800 ;
        RECT 4.400 154.680 1752.380 156.080 ;
        RECT 1.445 149.960 1752.380 154.680 ;
        RECT 4.400 148.560 1752.380 149.960 ;
        RECT 1.445 143.840 1752.380 148.560 ;
        RECT 4.400 142.440 1752.380 143.840 ;
        RECT 1.445 137.720 1752.380 142.440 ;
        RECT 4.400 136.320 1751.980 137.720 ;
        RECT 1.445 131.600 1752.380 136.320 ;
        RECT 4.400 130.200 1752.380 131.600 ;
        RECT 1.445 125.480 1752.380 130.200 ;
        RECT 4.400 124.080 1752.380 125.480 ;
        RECT 1.445 119.360 1752.380 124.080 ;
        RECT 4.400 117.960 1752.380 119.360 ;
        RECT 1.445 113.240 1752.380 117.960 ;
        RECT 4.400 111.840 1752.380 113.240 ;
        RECT 1.445 107.120 1752.380 111.840 ;
        RECT 4.400 105.720 1752.380 107.120 ;
        RECT 1.445 101.000 1752.380 105.720 ;
        RECT 4.400 99.600 1752.380 101.000 ;
        RECT 1.445 98.280 1752.380 99.600 ;
        RECT 1.445 96.880 1751.980 98.280 ;
        RECT 1.445 94.880 1752.380 96.880 ;
        RECT 4.400 93.480 1752.380 94.880 ;
        RECT 1.445 88.760 1752.380 93.480 ;
        RECT 4.400 87.360 1752.380 88.760 ;
        RECT 1.445 82.640 1752.380 87.360 ;
        RECT 4.400 81.240 1752.380 82.640 ;
        RECT 1.445 76.520 1752.380 81.240 ;
        RECT 4.400 75.120 1752.380 76.520 ;
        RECT 1.445 70.400 1752.380 75.120 ;
        RECT 4.400 69.000 1752.380 70.400 ;
        RECT 1.445 64.280 1752.380 69.000 ;
        RECT 4.400 62.880 1752.380 64.280 ;
        RECT 1.445 58.840 1752.380 62.880 ;
        RECT 1.445 58.160 1751.980 58.840 ;
        RECT 4.400 57.440 1751.980 58.160 ;
        RECT 4.400 56.760 1752.380 57.440 ;
        RECT 1.445 52.040 1752.380 56.760 ;
        RECT 4.400 50.640 1752.380 52.040 ;
        RECT 1.445 45.920 1752.380 50.640 ;
        RECT 4.400 44.520 1752.380 45.920 ;
        RECT 1.445 39.800 1752.380 44.520 ;
        RECT 4.400 38.400 1752.380 39.800 ;
        RECT 1.445 33.680 1752.380 38.400 ;
        RECT 4.400 32.280 1752.380 33.680 ;
        RECT 1.445 27.560 1752.380 32.280 ;
        RECT 4.400 26.160 1752.380 27.560 ;
        RECT 1.445 21.440 1752.380 26.160 ;
        RECT 4.400 20.080 1752.380 21.440 ;
        RECT 4.400 20.040 1751.980 20.080 ;
        RECT 1.445 18.680 1751.980 20.040 ;
        RECT 1.445 15.320 1752.380 18.680 ;
        RECT 4.400 13.920 1752.380 15.320 ;
        RECT 1.445 9.200 1752.380 13.920 ;
        RECT 4.400 7.800 1752.380 9.200 ;
        RECT 1.445 3.760 1752.380 7.800 ;
        RECT 4.400 2.895 1752.380 3.760 ;
      LAYER met4 ;
        RECT 3.975 1755.040 1660.305 1766.465 ;
        RECT 3.975 11.735 20.640 1755.040 ;
        RECT 23.040 11.735 97.440 1755.040 ;
        RECT 99.840 11.735 174.240 1755.040 ;
        RECT 176.640 11.735 251.040 1755.040 ;
        RECT 253.440 11.735 327.840 1755.040 ;
        RECT 330.240 11.735 404.640 1755.040 ;
        RECT 407.040 11.735 481.440 1755.040 ;
        RECT 483.840 11.735 558.240 1755.040 ;
        RECT 560.640 11.735 635.040 1755.040 ;
        RECT 637.440 11.735 711.840 1755.040 ;
        RECT 714.240 11.735 788.640 1755.040 ;
        RECT 791.040 11.735 865.440 1755.040 ;
        RECT 867.840 11.735 942.240 1755.040 ;
        RECT 944.640 11.735 1019.040 1755.040 ;
        RECT 1021.440 11.735 1095.840 1755.040 ;
        RECT 1098.240 11.735 1172.640 1755.040 ;
        RECT 1175.040 11.735 1249.440 1755.040 ;
        RECT 1251.840 11.735 1326.240 1755.040 ;
        RECT 1328.640 11.735 1403.040 1755.040 ;
        RECT 1405.440 11.735 1479.840 1755.040 ;
        RECT 1482.240 11.735 1556.640 1755.040 ;
        RECT 1559.040 11.735 1633.440 1755.040 ;
        RECT 1635.840 11.735 1660.305 1755.040 ;
  END
END Marmot
END LIBRARY

