module user_project_wrapper (user_clock2,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \data_arrays_0_0_ext_ram_addr1[0] ;
 wire \data_arrays_0_0_ext_ram_addr1[1] ;
 wire \data_arrays_0_0_ext_ram_addr1[2] ;
 wire \data_arrays_0_0_ext_ram_addr1[3] ;
 wire \data_arrays_0_0_ext_ram_addr1[4] ;
 wire \data_arrays_0_0_ext_ram_addr1[5] ;
 wire \data_arrays_0_0_ext_ram_addr1[6] ;
 wire \data_arrays_0_0_ext_ram_addr1[7] ;
 wire \data_arrays_0_0_ext_ram_addr1[8] ;
 wire \data_arrays_0_0_ext_ram_addr[0] ;
 wire \data_arrays_0_0_ext_ram_addr[1] ;
 wire \data_arrays_0_0_ext_ram_addr[2] ;
 wire \data_arrays_0_0_ext_ram_addr[3] ;
 wire \data_arrays_0_0_ext_ram_addr[4] ;
 wire \data_arrays_0_0_ext_ram_addr[5] ;
 wire \data_arrays_0_0_ext_ram_addr[6] ;
 wire \data_arrays_0_0_ext_ram_addr[7] ;
 wire \data_arrays_0_0_ext_ram_addr[8] ;
 wire data_arrays_0_0_ext_ram_clk0;
 wire data_arrays_0_0_ext_ram_clk1;
 wire data_arrays_0_0_ext_ram_clk2;
 wire data_arrays_0_0_ext_ram_clk3;
 wire \data_arrays_0_0_ext_ram_csb1[0] ;
 wire \data_arrays_0_0_ext_ram_csb1[1] ;
 wire \data_arrays_0_0_ext_ram_csb1[2] ;
 wire \data_arrays_0_0_ext_ram_csb1[3] ;
 wire \data_arrays_0_0_ext_ram_csb1[4] ;
 wire \data_arrays_0_0_ext_ram_csb1[5] ;
 wire \data_arrays_0_0_ext_ram_csb1[6] ;
 wire \data_arrays_0_0_ext_ram_csb1[7] ;
 wire \data_arrays_0_0_ext_ram_csb[0] ;
 wire \data_arrays_0_0_ext_ram_csb[1] ;
 wire \data_arrays_0_0_ext_ram_csb[2] ;
 wire \data_arrays_0_0_ext_ram_csb[3] ;
 wire \data_arrays_0_0_ext_ram_rdata0[0] ;
 wire \data_arrays_0_0_ext_ram_rdata0[10] ;
 wire \data_arrays_0_0_ext_ram_rdata0[11] ;
 wire \data_arrays_0_0_ext_ram_rdata0[12] ;
 wire \data_arrays_0_0_ext_ram_rdata0[13] ;
 wire \data_arrays_0_0_ext_ram_rdata0[14] ;
 wire \data_arrays_0_0_ext_ram_rdata0[15] ;
 wire \data_arrays_0_0_ext_ram_rdata0[16] ;
 wire \data_arrays_0_0_ext_ram_rdata0[17] ;
 wire \data_arrays_0_0_ext_ram_rdata0[18] ;
 wire \data_arrays_0_0_ext_ram_rdata0[19] ;
 wire \data_arrays_0_0_ext_ram_rdata0[1] ;
 wire \data_arrays_0_0_ext_ram_rdata0[20] ;
 wire \data_arrays_0_0_ext_ram_rdata0[21] ;
 wire \data_arrays_0_0_ext_ram_rdata0[22] ;
 wire \data_arrays_0_0_ext_ram_rdata0[23] ;
 wire \data_arrays_0_0_ext_ram_rdata0[24] ;
 wire \data_arrays_0_0_ext_ram_rdata0[25] ;
 wire \data_arrays_0_0_ext_ram_rdata0[26] ;
 wire \data_arrays_0_0_ext_ram_rdata0[27] ;
 wire \data_arrays_0_0_ext_ram_rdata0[28] ;
 wire \data_arrays_0_0_ext_ram_rdata0[29] ;
 wire \data_arrays_0_0_ext_ram_rdata0[2] ;
 wire \data_arrays_0_0_ext_ram_rdata0[30] ;
 wire \data_arrays_0_0_ext_ram_rdata0[31] ;
 wire \data_arrays_0_0_ext_ram_rdata0[32] ;
 wire \data_arrays_0_0_ext_ram_rdata0[33] ;
 wire \data_arrays_0_0_ext_ram_rdata0[34] ;
 wire \data_arrays_0_0_ext_ram_rdata0[35] ;
 wire \data_arrays_0_0_ext_ram_rdata0[36] ;
 wire \data_arrays_0_0_ext_ram_rdata0[37] ;
 wire \data_arrays_0_0_ext_ram_rdata0[38] ;
 wire \data_arrays_0_0_ext_ram_rdata0[39] ;
 wire \data_arrays_0_0_ext_ram_rdata0[3] ;
 wire \data_arrays_0_0_ext_ram_rdata0[40] ;
 wire \data_arrays_0_0_ext_ram_rdata0[41] ;
 wire \data_arrays_0_0_ext_ram_rdata0[42] ;
 wire \data_arrays_0_0_ext_ram_rdata0[43] ;
 wire \data_arrays_0_0_ext_ram_rdata0[44] ;
 wire \data_arrays_0_0_ext_ram_rdata0[45] ;
 wire \data_arrays_0_0_ext_ram_rdata0[46] ;
 wire \data_arrays_0_0_ext_ram_rdata0[47] ;
 wire \data_arrays_0_0_ext_ram_rdata0[48] ;
 wire \data_arrays_0_0_ext_ram_rdata0[49] ;
 wire \data_arrays_0_0_ext_ram_rdata0[4] ;
 wire \data_arrays_0_0_ext_ram_rdata0[50] ;
 wire \data_arrays_0_0_ext_ram_rdata0[51] ;
 wire \data_arrays_0_0_ext_ram_rdata0[52] ;
 wire \data_arrays_0_0_ext_ram_rdata0[53] ;
 wire \data_arrays_0_0_ext_ram_rdata0[54] ;
 wire \data_arrays_0_0_ext_ram_rdata0[55] ;
 wire \data_arrays_0_0_ext_ram_rdata0[56] ;
 wire \data_arrays_0_0_ext_ram_rdata0[57] ;
 wire \data_arrays_0_0_ext_ram_rdata0[58] ;
 wire \data_arrays_0_0_ext_ram_rdata0[59] ;
 wire \data_arrays_0_0_ext_ram_rdata0[5] ;
 wire \data_arrays_0_0_ext_ram_rdata0[60] ;
 wire \data_arrays_0_0_ext_ram_rdata0[61] ;
 wire \data_arrays_0_0_ext_ram_rdata0[62] ;
 wire \data_arrays_0_0_ext_ram_rdata0[63] ;
 wire \data_arrays_0_0_ext_ram_rdata0[6] ;
 wire \data_arrays_0_0_ext_ram_rdata0[7] ;
 wire \data_arrays_0_0_ext_ram_rdata0[8] ;
 wire \data_arrays_0_0_ext_ram_rdata0[9] ;
 wire \data_arrays_0_0_ext_ram_rdata1[0] ;
 wire \data_arrays_0_0_ext_ram_rdata1[10] ;
 wire \data_arrays_0_0_ext_ram_rdata1[11] ;
 wire \data_arrays_0_0_ext_ram_rdata1[12] ;
 wire \data_arrays_0_0_ext_ram_rdata1[13] ;
 wire \data_arrays_0_0_ext_ram_rdata1[14] ;
 wire \data_arrays_0_0_ext_ram_rdata1[15] ;
 wire \data_arrays_0_0_ext_ram_rdata1[16] ;
 wire \data_arrays_0_0_ext_ram_rdata1[17] ;
 wire \data_arrays_0_0_ext_ram_rdata1[18] ;
 wire \data_arrays_0_0_ext_ram_rdata1[19] ;
 wire \data_arrays_0_0_ext_ram_rdata1[1] ;
 wire \data_arrays_0_0_ext_ram_rdata1[20] ;
 wire \data_arrays_0_0_ext_ram_rdata1[21] ;
 wire \data_arrays_0_0_ext_ram_rdata1[22] ;
 wire \data_arrays_0_0_ext_ram_rdata1[23] ;
 wire \data_arrays_0_0_ext_ram_rdata1[24] ;
 wire \data_arrays_0_0_ext_ram_rdata1[25] ;
 wire \data_arrays_0_0_ext_ram_rdata1[26] ;
 wire \data_arrays_0_0_ext_ram_rdata1[27] ;
 wire \data_arrays_0_0_ext_ram_rdata1[28] ;
 wire \data_arrays_0_0_ext_ram_rdata1[29] ;
 wire \data_arrays_0_0_ext_ram_rdata1[2] ;
 wire \data_arrays_0_0_ext_ram_rdata1[30] ;
 wire \data_arrays_0_0_ext_ram_rdata1[31] ;
 wire \data_arrays_0_0_ext_ram_rdata1[32] ;
 wire \data_arrays_0_0_ext_ram_rdata1[33] ;
 wire \data_arrays_0_0_ext_ram_rdata1[34] ;
 wire \data_arrays_0_0_ext_ram_rdata1[35] ;
 wire \data_arrays_0_0_ext_ram_rdata1[36] ;
 wire \data_arrays_0_0_ext_ram_rdata1[37] ;
 wire \data_arrays_0_0_ext_ram_rdata1[38] ;
 wire \data_arrays_0_0_ext_ram_rdata1[39] ;
 wire \data_arrays_0_0_ext_ram_rdata1[3] ;
 wire \data_arrays_0_0_ext_ram_rdata1[40] ;
 wire \data_arrays_0_0_ext_ram_rdata1[41] ;
 wire \data_arrays_0_0_ext_ram_rdata1[42] ;
 wire \data_arrays_0_0_ext_ram_rdata1[43] ;
 wire \data_arrays_0_0_ext_ram_rdata1[44] ;
 wire \data_arrays_0_0_ext_ram_rdata1[45] ;
 wire \data_arrays_0_0_ext_ram_rdata1[46] ;
 wire \data_arrays_0_0_ext_ram_rdata1[47] ;
 wire \data_arrays_0_0_ext_ram_rdata1[48] ;
 wire \data_arrays_0_0_ext_ram_rdata1[49] ;
 wire \data_arrays_0_0_ext_ram_rdata1[4] ;
 wire \data_arrays_0_0_ext_ram_rdata1[50] ;
 wire \data_arrays_0_0_ext_ram_rdata1[51] ;
 wire \data_arrays_0_0_ext_ram_rdata1[52] ;
 wire \data_arrays_0_0_ext_ram_rdata1[53] ;
 wire \data_arrays_0_0_ext_ram_rdata1[54] ;
 wire \data_arrays_0_0_ext_ram_rdata1[55] ;
 wire \data_arrays_0_0_ext_ram_rdata1[56] ;
 wire \data_arrays_0_0_ext_ram_rdata1[57] ;
 wire \data_arrays_0_0_ext_ram_rdata1[58] ;
 wire \data_arrays_0_0_ext_ram_rdata1[59] ;
 wire \data_arrays_0_0_ext_ram_rdata1[5] ;
 wire \data_arrays_0_0_ext_ram_rdata1[60] ;
 wire \data_arrays_0_0_ext_ram_rdata1[61] ;
 wire \data_arrays_0_0_ext_ram_rdata1[62] ;
 wire \data_arrays_0_0_ext_ram_rdata1[63] ;
 wire \data_arrays_0_0_ext_ram_rdata1[6] ;
 wire \data_arrays_0_0_ext_ram_rdata1[7] ;
 wire \data_arrays_0_0_ext_ram_rdata1[8] ;
 wire \data_arrays_0_0_ext_ram_rdata1[9] ;
 wire \data_arrays_0_0_ext_ram_rdata2[0] ;
 wire \data_arrays_0_0_ext_ram_rdata2[10] ;
 wire \data_arrays_0_0_ext_ram_rdata2[11] ;
 wire \data_arrays_0_0_ext_ram_rdata2[12] ;
 wire \data_arrays_0_0_ext_ram_rdata2[13] ;
 wire \data_arrays_0_0_ext_ram_rdata2[14] ;
 wire \data_arrays_0_0_ext_ram_rdata2[15] ;
 wire \data_arrays_0_0_ext_ram_rdata2[16] ;
 wire \data_arrays_0_0_ext_ram_rdata2[17] ;
 wire \data_arrays_0_0_ext_ram_rdata2[18] ;
 wire \data_arrays_0_0_ext_ram_rdata2[19] ;
 wire \data_arrays_0_0_ext_ram_rdata2[1] ;
 wire \data_arrays_0_0_ext_ram_rdata2[20] ;
 wire \data_arrays_0_0_ext_ram_rdata2[21] ;
 wire \data_arrays_0_0_ext_ram_rdata2[22] ;
 wire \data_arrays_0_0_ext_ram_rdata2[23] ;
 wire \data_arrays_0_0_ext_ram_rdata2[24] ;
 wire \data_arrays_0_0_ext_ram_rdata2[25] ;
 wire \data_arrays_0_0_ext_ram_rdata2[26] ;
 wire \data_arrays_0_0_ext_ram_rdata2[27] ;
 wire \data_arrays_0_0_ext_ram_rdata2[28] ;
 wire \data_arrays_0_0_ext_ram_rdata2[29] ;
 wire \data_arrays_0_0_ext_ram_rdata2[2] ;
 wire \data_arrays_0_0_ext_ram_rdata2[30] ;
 wire \data_arrays_0_0_ext_ram_rdata2[31] ;
 wire \data_arrays_0_0_ext_ram_rdata2[32] ;
 wire \data_arrays_0_0_ext_ram_rdata2[33] ;
 wire \data_arrays_0_0_ext_ram_rdata2[34] ;
 wire \data_arrays_0_0_ext_ram_rdata2[35] ;
 wire \data_arrays_0_0_ext_ram_rdata2[36] ;
 wire \data_arrays_0_0_ext_ram_rdata2[37] ;
 wire \data_arrays_0_0_ext_ram_rdata2[38] ;
 wire \data_arrays_0_0_ext_ram_rdata2[39] ;
 wire \data_arrays_0_0_ext_ram_rdata2[3] ;
 wire \data_arrays_0_0_ext_ram_rdata2[40] ;
 wire \data_arrays_0_0_ext_ram_rdata2[41] ;
 wire \data_arrays_0_0_ext_ram_rdata2[42] ;
 wire \data_arrays_0_0_ext_ram_rdata2[43] ;
 wire \data_arrays_0_0_ext_ram_rdata2[44] ;
 wire \data_arrays_0_0_ext_ram_rdata2[45] ;
 wire \data_arrays_0_0_ext_ram_rdata2[46] ;
 wire \data_arrays_0_0_ext_ram_rdata2[47] ;
 wire \data_arrays_0_0_ext_ram_rdata2[48] ;
 wire \data_arrays_0_0_ext_ram_rdata2[49] ;
 wire \data_arrays_0_0_ext_ram_rdata2[4] ;
 wire \data_arrays_0_0_ext_ram_rdata2[50] ;
 wire \data_arrays_0_0_ext_ram_rdata2[51] ;
 wire \data_arrays_0_0_ext_ram_rdata2[52] ;
 wire \data_arrays_0_0_ext_ram_rdata2[53] ;
 wire \data_arrays_0_0_ext_ram_rdata2[54] ;
 wire \data_arrays_0_0_ext_ram_rdata2[55] ;
 wire \data_arrays_0_0_ext_ram_rdata2[56] ;
 wire \data_arrays_0_0_ext_ram_rdata2[57] ;
 wire \data_arrays_0_0_ext_ram_rdata2[58] ;
 wire \data_arrays_0_0_ext_ram_rdata2[59] ;
 wire \data_arrays_0_0_ext_ram_rdata2[5] ;
 wire \data_arrays_0_0_ext_ram_rdata2[60] ;
 wire \data_arrays_0_0_ext_ram_rdata2[61] ;
 wire \data_arrays_0_0_ext_ram_rdata2[62] ;
 wire \data_arrays_0_0_ext_ram_rdata2[63] ;
 wire \data_arrays_0_0_ext_ram_rdata2[6] ;
 wire \data_arrays_0_0_ext_ram_rdata2[7] ;
 wire \data_arrays_0_0_ext_ram_rdata2[8] ;
 wire \data_arrays_0_0_ext_ram_rdata2[9] ;
 wire \data_arrays_0_0_ext_ram_rdata3[0] ;
 wire \data_arrays_0_0_ext_ram_rdata3[10] ;
 wire \data_arrays_0_0_ext_ram_rdata3[11] ;
 wire \data_arrays_0_0_ext_ram_rdata3[12] ;
 wire \data_arrays_0_0_ext_ram_rdata3[13] ;
 wire \data_arrays_0_0_ext_ram_rdata3[14] ;
 wire \data_arrays_0_0_ext_ram_rdata3[15] ;
 wire \data_arrays_0_0_ext_ram_rdata3[16] ;
 wire \data_arrays_0_0_ext_ram_rdata3[17] ;
 wire \data_arrays_0_0_ext_ram_rdata3[18] ;
 wire \data_arrays_0_0_ext_ram_rdata3[19] ;
 wire \data_arrays_0_0_ext_ram_rdata3[1] ;
 wire \data_arrays_0_0_ext_ram_rdata3[20] ;
 wire \data_arrays_0_0_ext_ram_rdata3[21] ;
 wire \data_arrays_0_0_ext_ram_rdata3[22] ;
 wire \data_arrays_0_0_ext_ram_rdata3[23] ;
 wire \data_arrays_0_0_ext_ram_rdata3[24] ;
 wire \data_arrays_0_0_ext_ram_rdata3[25] ;
 wire \data_arrays_0_0_ext_ram_rdata3[26] ;
 wire \data_arrays_0_0_ext_ram_rdata3[27] ;
 wire \data_arrays_0_0_ext_ram_rdata3[28] ;
 wire \data_arrays_0_0_ext_ram_rdata3[29] ;
 wire \data_arrays_0_0_ext_ram_rdata3[2] ;
 wire \data_arrays_0_0_ext_ram_rdata3[30] ;
 wire \data_arrays_0_0_ext_ram_rdata3[31] ;
 wire \data_arrays_0_0_ext_ram_rdata3[32] ;
 wire \data_arrays_0_0_ext_ram_rdata3[33] ;
 wire \data_arrays_0_0_ext_ram_rdata3[34] ;
 wire \data_arrays_0_0_ext_ram_rdata3[35] ;
 wire \data_arrays_0_0_ext_ram_rdata3[36] ;
 wire \data_arrays_0_0_ext_ram_rdata3[37] ;
 wire \data_arrays_0_0_ext_ram_rdata3[38] ;
 wire \data_arrays_0_0_ext_ram_rdata3[39] ;
 wire \data_arrays_0_0_ext_ram_rdata3[3] ;
 wire \data_arrays_0_0_ext_ram_rdata3[40] ;
 wire \data_arrays_0_0_ext_ram_rdata3[41] ;
 wire \data_arrays_0_0_ext_ram_rdata3[42] ;
 wire \data_arrays_0_0_ext_ram_rdata3[43] ;
 wire \data_arrays_0_0_ext_ram_rdata3[44] ;
 wire \data_arrays_0_0_ext_ram_rdata3[45] ;
 wire \data_arrays_0_0_ext_ram_rdata3[46] ;
 wire \data_arrays_0_0_ext_ram_rdata3[47] ;
 wire \data_arrays_0_0_ext_ram_rdata3[48] ;
 wire \data_arrays_0_0_ext_ram_rdata3[49] ;
 wire \data_arrays_0_0_ext_ram_rdata3[4] ;
 wire \data_arrays_0_0_ext_ram_rdata3[50] ;
 wire \data_arrays_0_0_ext_ram_rdata3[51] ;
 wire \data_arrays_0_0_ext_ram_rdata3[52] ;
 wire \data_arrays_0_0_ext_ram_rdata3[53] ;
 wire \data_arrays_0_0_ext_ram_rdata3[54] ;
 wire \data_arrays_0_0_ext_ram_rdata3[55] ;
 wire \data_arrays_0_0_ext_ram_rdata3[56] ;
 wire \data_arrays_0_0_ext_ram_rdata3[57] ;
 wire \data_arrays_0_0_ext_ram_rdata3[58] ;
 wire \data_arrays_0_0_ext_ram_rdata3[59] ;
 wire \data_arrays_0_0_ext_ram_rdata3[5] ;
 wire \data_arrays_0_0_ext_ram_rdata3[60] ;
 wire \data_arrays_0_0_ext_ram_rdata3[61] ;
 wire \data_arrays_0_0_ext_ram_rdata3[62] ;
 wire \data_arrays_0_0_ext_ram_rdata3[63] ;
 wire \data_arrays_0_0_ext_ram_rdata3[6] ;
 wire \data_arrays_0_0_ext_ram_rdata3[7] ;
 wire \data_arrays_0_0_ext_ram_rdata3[8] ;
 wire \data_arrays_0_0_ext_ram_rdata3[9] ;
 wire \data_arrays_0_0_ext_ram_wdata[0] ;
 wire \data_arrays_0_0_ext_ram_wdata[10] ;
 wire \data_arrays_0_0_ext_ram_wdata[11] ;
 wire \data_arrays_0_0_ext_ram_wdata[12] ;
 wire \data_arrays_0_0_ext_ram_wdata[13] ;
 wire \data_arrays_0_0_ext_ram_wdata[14] ;
 wire \data_arrays_0_0_ext_ram_wdata[15] ;
 wire \data_arrays_0_0_ext_ram_wdata[16] ;
 wire \data_arrays_0_0_ext_ram_wdata[17] ;
 wire \data_arrays_0_0_ext_ram_wdata[18] ;
 wire \data_arrays_0_0_ext_ram_wdata[19] ;
 wire \data_arrays_0_0_ext_ram_wdata[1] ;
 wire \data_arrays_0_0_ext_ram_wdata[20] ;
 wire \data_arrays_0_0_ext_ram_wdata[21] ;
 wire \data_arrays_0_0_ext_ram_wdata[22] ;
 wire \data_arrays_0_0_ext_ram_wdata[23] ;
 wire \data_arrays_0_0_ext_ram_wdata[24] ;
 wire \data_arrays_0_0_ext_ram_wdata[25] ;
 wire \data_arrays_0_0_ext_ram_wdata[26] ;
 wire \data_arrays_0_0_ext_ram_wdata[27] ;
 wire \data_arrays_0_0_ext_ram_wdata[28] ;
 wire \data_arrays_0_0_ext_ram_wdata[29] ;
 wire \data_arrays_0_0_ext_ram_wdata[2] ;
 wire \data_arrays_0_0_ext_ram_wdata[30] ;
 wire \data_arrays_0_0_ext_ram_wdata[31] ;
 wire \data_arrays_0_0_ext_ram_wdata[32] ;
 wire \data_arrays_0_0_ext_ram_wdata[33] ;
 wire \data_arrays_0_0_ext_ram_wdata[34] ;
 wire \data_arrays_0_0_ext_ram_wdata[35] ;
 wire \data_arrays_0_0_ext_ram_wdata[36] ;
 wire \data_arrays_0_0_ext_ram_wdata[37] ;
 wire \data_arrays_0_0_ext_ram_wdata[38] ;
 wire \data_arrays_0_0_ext_ram_wdata[39] ;
 wire \data_arrays_0_0_ext_ram_wdata[3] ;
 wire \data_arrays_0_0_ext_ram_wdata[40] ;
 wire \data_arrays_0_0_ext_ram_wdata[41] ;
 wire \data_arrays_0_0_ext_ram_wdata[42] ;
 wire \data_arrays_0_0_ext_ram_wdata[43] ;
 wire \data_arrays_0_0_ext_ram_wdata[44] ;
 wire \data_arrays_0_0_ext_ram_wdata[45] ;
 wire \data_arrays_0_0_ext_ram_wdata[46] ;
 wire \data_arrays_0_0_ext_ram_wdata[47] ;
 wire \data_arrays_0_0_ext_ram_wdata[48] ;
 wire \data_arrays_0_0_ext_ram_wdata[49] ;
 wire \data_arrays_0_0_ext_ram_wdata[4] ;
 wire \data_arrays_0_0_ext_ram_wdata[50] ;
 wire \data_arrays_0_0_ext_ram_wdata[51] ;
 wire \data_arrays_0_0_ext_ram_wdata[52] ;
 wire \data_arrays_0_0_ext_ram_wdata[53] ;
 wire \data_arrays_0_0_ext_ram_wdata[54] ;
 wire \data_arrays_0_0_ext_ram_wdata[55] ;
 wire \data_arrays_0_0_ext_ram_wdata[56] ;
 wire \data_arrays_0_0_ext_ram_wdata[57] ;
 wire \data_arrays_0_0_ext_ram_wdata[58] ;
 wire \data_arrays_0_0_ext_ram_wdata[59] ;
 wire \data_arrays_0_0_ext_ram_wdata[5] ;
 wire \data_arrays_0_0_ext_ram_wdata[60] ;
 wire \data_arrays_0_0_ext_ram_wdata[61] ;
 wire \data_arrays_0_0_ext_ram_wdata[62] ;
 wire \data_arrays_0_0_ext_ram_wdata[63] ;
 wire \data_arrays_0_0_ext_ram_wdata[6] ;
 wire \data_arrays_0_0_ext_ram_wdata[7] ;
 wire \data_arrays_0_0_ext_ram_wdata[8] ;
 wire \data_arrays_0_0_ext_ram_wdata[9] ;
 wire data_arrays_0_0_ext_ram_web;
 wire \data_arrays_0_0_ext_ram_wmask[0] ;
 wire \data_arrays_0_0_ext_ram_wmask[1] ;
 wire \ram_clk_delay_sel[0] ;
 wire \ram_clk_delay_sel[10] ;
 wire \ram_clk_delay_sel[11] ;
 wire \ram_clk_delay_sel[12] ;
 wire \ram_clk_delay_sel[13] ;
 wire \ram_clk_delay_sel[14] ;
 wire \ram_clk_delay_sel[15] ;
 wire \ram_clk_delay_sel[16] ;
 wire \ram_clk_delay_sel[17] ;
 wire \ram_clk_delay_sel[18] ;
 wire \ram_clk_delay_sel[19] ;
 wire \ram_clk_delay_sel[1] ;
 wire \ram_clk_delay_sel[20] ;
 wire \ram_clk_delay_sel[21] ;
 wire \ram_clk_delay_sel[22] ;
 wire \ram_clk_delay_sel[23] ;
 wire \ram_clk_delay_sel[24] ;
 wire \ram_clk_delay_sel[25] ;
 wire \ram_clk_delay_sel[26] ;
 wire \ram_clk_delay_sel[27] ;
 wire \ram_clk_delay_sel[28] ;
 wire \ram_clk_delay_sel[29] ;
 wire \ram_clk_delay_sel[2] ;
 wire \ram_clk_delay_sel[30] ;
 wire \ram_clk_delay_sel[31] ;
 wire \ram_clk_delay_sel[3] ;
 wire \ram_clk_delay_sel[4] ;
 wire \ram_clk_delay_sel[5] ;
 wire \ram_clk_delay_sel[6] ;
 wire \ram_clk_delay_sel[7] ;
 wire \ram_clk_delay_sel[8] ;
 wire \ram_clk_delay_sel[9] ;
 wire \tag_array_ext_ram_addr1[0] ;
 wire \tag_array_ext_ram_addr1[1] ;
 wire \tag_array_ext_ram_addr1[2] ;
 wire \tag_array_ext_ram_addr1[3] ;
 wire \tag_array_ext_ram_addr1[4] ;
 wire \tag_array_ext_ram_addr1[5] ;
 wire \tag_array_ext_ram_addr1[6] ;
 wire \tag_array_ext_ram_addr1[7] ;
 wire \tag_array_ext_ram_addr[0] ;
 wire \tag_array_ext_ram_addr[1] ;
 wire \tag_array_ext_ram_addr[2] ;
 wire \tag_array_ext_ram_addr[3] ;
 wire \tag_array_ext_ram_addr[4] ;
 wire \tag_array_ext_ram_addr[5] ;
 wire \tag_array_ext_ram_addr[6] ;
 wire \tag_array_ext_ram_addr[7] ;
 wire tag_array_ext_ram_clk;
 wire tag_array_ext_ram_csb;
 wire \tag_array_ext_ram_csb1[0] ;
 wire \tag_array_ext_ram_csb1[1] ;
 wire \tag_array_ext_ram_rdata0[0] ;
 wire \tag_array_ext_ram_rdata0[10] ;
 wire \tag_array_ext_ram_rdata0[11] ;
 wire \tag_array_ext_ram_rdata0[12] ;
 wire \tag_array_ext_ram_rdata0[13] ;
 wire \tag_array_ext_ram_rdata0[14] ;
 wire \tag_array_ext_ram_rdata0[15] ;
 wire \tag_array_ext_ram_rdata0[16] ;
 wire \tag_array_ext_ram_rdata0[17] ;
 wire \tag_array_ext_ram_rdata0[18] ;
 wire \tag_array_ext_ram_rdata0[19] ;
 wire \tag_array_ext_ram_rdata0[1] ;
 wire \tag_array_ext_ram_rdata0[20] ;
 wire \tag_array_ext_ram_rdata0[21] ;
 wire \tag_array_ext_ram_rdata0[22] ;
 wire \tag_array_ext_ram_rdata0[23] ;
 wire \tag_array_ext_ram_rdata0[24] ;
 wire \tag_array_ext_ram_rdata0[25] ;
 wire \tag_array_ext_ram_rdata0[26] ;
 wire \tag_array_ext_ram_rdata0[27] ;
 wire \tag_array_ext_ram_rdata0[28] ;
 wire \tag_array_ext_ram_rdata0[29] ;
 wire \tag_array_ext_ram_rdata0[2] ;
 wire \tag_array_ext_ram_rdata0[30] ;
 wire \tag_array_ext_ram_rdata0[31] ;
 wire \tag_array_ext_ram_rdata0[3] ;
 wire \tag_array_ext_ram_rdata0[4] ;
 wire \tag_array_ext_ram_rdata0[5] ;
 wire \tag_array_ext_ram_rdata0[6] ;
 wire \tag_array_ext_ram_rdata0[7] ;
 wire \tag_array_ext_ram_rdata0[8] ;
 wire \tag_array_ext_ram_rdata0[9] ;
 wire \tag_array_ext_ram_rdata1[0] ;
 wire \tag_array_ext_ram_rdata1[10] ;
 wire \tag_array_ext_ram_rdata1[11] ;
 wire \tag_array_ext_ram_rdata1[12] ;
 wire \tag_array_ext_ram_rdata1[13] ;
 wire \tag_array_ext_ram_rdata1[14] ;
 wire \tag_array_ext_ram_rdata1[15] ;
 wire \tag_array_ext_ram_rdata1[16] ;
 wire \tag_array_ext_ram_rdata1[17] ;
 wire \tag_array_ext_ram_rdata1[18] ;
 wire \tag_array_ext_ram_rdata1[19] ;
 wire \tag_array_ext_ram_rdata1[1] ;
 wire \tag_array_ext_ram_rdata1[20] ;
 wire \tag_array_ext_ram_rdata1[21] ;
 wire \tag_array_ext_ram_rdata1[22] ;
 wire \tag_array_ext_ram_rdata1[23] ;
 wire \tag_array_ext_ram_rdata1[24] ;
 wire \tag_array_ext_ram_rdata1[25] ;
 wire \tag_array_ext_ram_rdata1[26] ;
 wire \tag_array_ext_ram_rdata1[27] ;
 wire \tag_array_ext_ram_rdata1[28] ;
 wire \tag_array_ext_ram_rdata1[29] ;
 wire \tag_array_ext_ram_rdata1[2] ;
 wire \tag_array_ext_ram_rdata1[30] ;
 wire \tag_array_ext_ram_rdata1[31] ;
 wire \tag_array_ext_ram_rdata1[3] ;
 wire \tag_array_ext_ram_rdata1[4] ;
 wire \tag_array_ext_ram_rdata1[5] ;
 wire \tag_array_ext_ram_rdata1[6] ;
 wire \tag_array_ext_ram_rdata1[7] ;
 wire \tag_array_ext_ram_rdata1[8] ;
 wire \tag_array_ext_ram_rdata1[9] ;
 wire \tag_array_ext_ram_wdata[0] ;
 wire \tag_array_ext_ram_wdata[10] ;
 wire \tag_array_ext_ram_wdata[11] ;
 wire \tag_array_ext_ram_wdata[12] ;
 wire \tag_array_ext_ram_wdata[13] ;
 wire \tag_array_ext_ram_wdata[14] ;
 wire \tag_array_ext_ram_wdata[15] ;
 wire \tag_array_ext_ram_wdata[16] ;
 wire \tag_array_ext_ram_wdata[17] ;
 wire \tag_array_ext_ram_wdata[18] ;
 wire \tag_array_ext_ram_wdata[19] ;
 wire \tag_array_ext_ram_wdata[1] ;
 wire \tag_array_ext_ram_wdata[20] ;
 wire \tag_array_ext_ram_wdata[21] ;
 wire \tag_array_ext_ram_wdata[22] ;
 wire \tag_array_ext_ram_wdata[23] ;
 wire \tag_array_ext_ram_wdata[24] ;
 wire \tag_array_ext_ram_wdata[25] ;
 wire \tag_array_ext_ram_wdata[26] ;
 wire \tag_array_ext_ram_wdata[27] ;
 wire \tag_array_ext_ram_wdata[28] ;
 wire \tag_array_ext_ram_wdata[29] ;
 wire \tag_array_ext_ram_wdata[2] ;
 wire \tag_array_ext_ram_wdata[30] ;
 wire \tag_array_ext_ram_wdata[31] ;
 wire \tag_array_ext_ram_wdata[32] ;
 wire \tag_array_ext_ram_wdata[33] ;
 wire \tag_array_ext_ram_wdata[34] ;
 wire \tag_array_ext_ram_wdata[35] ;
 wire \tag_array_ext_ram_wdata[36] ;
 wire \tag_array_ext_ram_wdata[37] ;
 wire \tag_array_ext_ram_wdata[38] ;
 wire \tag_array_ext_ram_wdata[39] ;
 wire \tag_array_ext_ram_wdata[3] ;
 wire \tag_array_ext_ram_wdata[40] ;
 wire \tag_array_ext_ram_wdata[41] ;
 wire \tag_array_ext_ram_wdata[42] ;
 wire \tag_array_ext_ram_wdata[43] ;
 wire \tag_array_ext_ram_wdata[44] ;
 wire \tag_array_ext_ram_wdata[45] ;
 wire \tag_array_ext_ram_wdata[46] ;
 wire \tag_array_ext_ram_wdata[47] ;
 wire \tag_array_ext_ram_wdata[48] ;
 wire \tag_array_ext_ram_wdata[49] ;
 wire \tag_array_ext_ram_wdata[4] ;
 wire \tag_array_ext_ram_wdata[50] ;
 wire \tag_array_ext_ram_wdata[51] ;
 wire \tag_array_ext_ram_wdata[52] ;
 wire \tag_array_ext_ram_wdata[53] ;
 wire \tag_array_ext_ram_wdata[54] ;
 wire \tag_array_ext_ram_wdata[55] ;
 wire \tag_array_ext_ram_wdata[56] ;
 wire \tag_array_ext_ram_wdata[57] ;
 wire \tag_array_ext_ram_wdata[58] ;
 wire \tag_array_ext_ram_wdata[59] ;
 wire \tag_array_ext_ram_wdata[5] ;
 wire \tag_array_ext_ram_wdata[60] ;
 wire \tag_array_ext_ram_wdata[61] ;
 wire \tag_array_ext_ram_wdata[62] ;
 wire \tag_array_ext_ram_wdata[63] ;
 wire \tag_array_ext_ram_wdata[6] ;
 wire \tag_array_ext_ram_wdata[7] ;
 wire \tag_array_ext_ram_wdata[8] ;
 wire \tag_array_ext_ram_wdata[9] ;
 wire tag_array_ext_ram_web;
 wire \tag_array_ext_ram_wmask[0] ;
 wire \tag_array_ext_ram_wmask[1] ;

 Marmot Marmot (.data_arrays_0_0_ext_ram_web(data_arrays_0_0_ext_ram_web),
    .tag_array_ext_ram_csb(tag_array_ext_ram_csb),
    .tag_array_ext_ram_web(tag_array_ext_ram_web),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .data_arrays_0_0_ext_ram_addr({\data_arrays_0_0_ext_ram_addr[8] ,
    \data_arrays_0_0_ext_ram_addr[7] ,
    \data_arrays_0_0_ext_ram_addr[6] ,
    \data_arrays_0_0_ext_ram_addr[5] ,
    \data_arrays_0_0_ext_ram_addr[4] ,
    \data_arrays_0_0_ext_ram_addr[3] ,
    \data_arrays_0_0_ext_ram_addr[2] ,
    \data_arrays_0_0_ext_ram_addr[1] ,
    \data_arrays_0_0_ext_ram_addr[0] }),
    .data_arrays_0_0_ext_ram_addr1({\data_arrays_0_0_ext_ram_addr1[8] ,
    \data_arrays_0_0_ext_ram_addr1[7] ,
    \data_arrays_0_0_ext_ram_addr1[6] ,
    \data_arrays_0_0_ext_ram_addr1[5] ,
    \data_arrays_0_0_ext_ram_addr1[4] ,
    \data_arrays_0_0_ext_ram_addr1[3] ,
    \data_arrays_0_0_ext_ram_addr1[2] ,
    \data_arrays_0_0_ext_ram_addr1[1] ,
    \data_arrays_0_0_ext_ram_addr1[0] }),
    .data_arrays_0_0_ext_ram_csb({\data_arrays_0_0_ext_ram_csb[3] ,
    \data_arrays_0_0_ext_ram_csb[2] ,
    \data_arrays_0_0_ext_ram_csb[1] ,
    \data_arrays_0_0_ext_ram_csb[0] }),
    .data_arrays_0_0_ext_ram_csb1({\data_arrays_0_0_ext_ram_csb1[7] ,
    \data_arrays_0_0_ext_ram_csb1[6] ,
    \data_arrays_0_0_ext_ram_csb1[5] ,
    \data_arrays_0_0_ext_ram_csb1[4] ,
    \data_arrays_0_0_ext_ram_csb1[3] ,
    \data_arrays_0_0_ext_ram_csb1[2] ,
    \data_arrays_0_0_ext_ram_csb1[1] ,
    \data_arrays_0_0_ext_ram_csb1[0] }),
    .data_arrays_0_0_ext_ram_rdata0({\data_arrays_0_0_ext_ram_rdata0[63] ,
    \data_arrays_0_0_ext_ram_rdata0[62] ,
    \data_arrays_0_0_ext_ram_rdata0[61] ,
    \data_arrays_0_0_ext_ram_rdata0[60] ,
    \data_arrays_0_0_ext_ram_rdata0[59] ,
    \data_arrays_0_0_ext_ram_rdata0[58] ,
    \data_arrays_0_0_ext_ram_rdata0[57] ,
    \data_arrays_0_0_ext_ram_rdata0[56] ,
    \data_arrays_0_0_ext_ram_rdata0[55] ,
    \data_arrays_0_0_ext_ram_rdata0[54] ,
    \data_arrays_0_0_ext_ram_rdata0[53] ,
    \data_arrays_0_0_ext_ram_rdata0[52] ,
    \data_arrays_0_0_ext_ram_rdata0[51] ,
    \data_arrays_0_0_ext_ram_rdata0[50] ,
    \data_arrays_0_0_ext_ram_rdata0[49] ,
    \data_arrays_0_0_ext_ram_rdata0[48] ,
    \data_arrays_0_0_ext_ram_rdata0[47] ,
    \data_arrays_0_0_ext_ram_rdata0[46] ,
    \data_arrays_0_0_ext_ram_rdata0[45] ,
    \data_arrays_0_0_ext_ram_rdata0[44] ,
    \data_arrays_0_0_ext_ram_rdata0[43] ,
    \data_arrays_0_0_ext_ram_rdata0[42] ,
    \data_arrays_0_0_ext_ram_rdata0[41] ,
    \data_arrays_0_0_ext_ram_rdata0[40] ,
    \data_arrays_0_0_ext_ram_rdata0[39] ,
    \data_arrays_0_0_ext_ram_rdata0[38] ,
    \data_arrays_0_0_ext_ram_rdata0[37] ,
    \data_arrays_0_0_ext_ram_rdata0[36] ,
    \data_arrays_0_0_ext_ram_rdata0[35] ,
    \data_arrays_0_0_ext_ram_rdata0[34] ,
    \data_arrays_0_0_ext_ram_rdata0[33] ,
    \data_arrays_0_0_ext_ram_rdata0[32] ,
    \data_arrays_0_0_ext_ram_rdata0[31] ,
    \data_arrays_0_0_ext_ram_rdata0[30] ,
    \data_arrays_0_0_ext_ram_rdata0[29] ,
    \data_arrays_0_0_ext_ram_rdata0[28] ,
    \data_arrays_0_0_ext_ram_rdata0[27] ,
    \data_arrays_0_0_ext_ram_rdata0[26] ,
    \data_arrays_0_0_ext_ram_rdata0[25] ,
    \data_arrays_0_0_ext_ram_rdata0[24] ,
    \data_arrays_0_0_ext_ram_rdata0[23] ,
    \data_arrays_0_0_ext_ram_rdata0[22] ,
    \data_arrays_0_0_ext_ram_rdata0[21] ,
    \data_arrays_0_0_ext_ram_rdata0[20] ,
    \data_arrays_0_0_ext_ram_rdata0[19] ,
    \data_arrays_0_0_ext_ram_rdata0[18] ,
    \data_arrays_0_0_ext_ram_rdata0[17] ,
    \data_arrays_0_0_ext_ram_rdata0[16] ,
    \data_arrays_0_0_ext_ram_rdata0[15] ,
    \data_arrays_0_0_ext_ram_rdata0[14] ,
    \data_arrays_0_0_ext_ram_rdata0[13] ,
    \data_arrays_0_0_ext_ram_rdata0[12] ,
    \data_arrays_0_0_ext_ram_rdata0[11] ,
    \data_arrays_0_0_ext_ram_rdata0[10] ,
    \data_arrays_0_0_ext_ram_rdata0[9] ,
    \data_arrays_0_0_ext_ram_rdata0[8] ,
    \data_arrays_0_0_ext_ram_rdata0[7] ,
    \data_arrays_0_0_ext_ram_rdata0[6] ,
    \data_arrays_0_0_ext_ram_rdata0[5] ,
    \data_arrays_0_0_ext_ram_rdata0[4] ,
    \data_arrays_0_0_ext_ram_rdata0[3] ,
    \data_arrays_0_0_ext_ram_rdata0[2] ,
    \data_arrays_0_0_ext_ram_rdata0[1] ,
    \data_arrays_0_0_ext_ram_rdata0[0] }),
    .data_arrays_0_0_ext_ram_rdata1({\data_arrays_0_0_ext_ram_rdata1[63] ,
    \data_arrays_0_0_ext_ram_rdata1[62] ,
    \data_arrays_0_0_ext_ram_rdata1[61] ,
    \data_arrays_0_0_ext_ram_rdata1[60] ,
    \data_arrays_0_0_ext_ram_rdata1[59] ,
    \data_arrays_0_0_ext_ram_rdata1[58] ,
    \data_arrays_0_0_ext_ram_rdata1[57] ,
    \data_arrays_0_0_ext_ram_rdata1[56] ,
    \data_arrays_0_0_ext_ram_rdata1[55] ,
    \data_arrays_0_0_ext_ram_rdata1[54] ,
    \data_arrays_0_0_ext_ram_rdata1[53] ,
    \data_arrays_0_0_ext_ram_rdata1[52] ,
    \data_arrays_0_0_ext_ram_rdata1[51] ,
    \data_arrays_0_0_ext_ram_rdata1[50] ,
    \data_arrays_0_0_ext_ram_rdata1[49] ,
    \data_arrays_0_0_ext_ram_rdata1[48] ,
    \data_arrays_0_0_ext_ram_rdata1[47] ,
    \data_arrays_0_0_ext_ram_rdata1[46] ,
    \data_arrays_0_0_ext_ram_rdata1[45] ,
    \data_arrays_0_0_ext_ram_rdata1[44] ,
    \data_arrays_0_0_ext_ram_rdata1[43] ,
    \data_arrays_0_0_ext_ram_rdata1[42] ,
    \data_arrays_0_0_ext_ram_rdata1[41] ,
    \data_arrays_0_0_ext_ram_rdata1[40] ,
    \data_arrays_0_0_ext_ram_rdata1[39] ,
    \data_arrays_0_0_ext_ram_rdata1[38] ,
    \data_arrays_0_0_ext_ram_rdata1[37] ,
    \data_arrays_0_0_ext_ram_rdata1[36] ,
    \data_arrays_0_0_ext_ram_rdata1[35] ,
    \data_arrays_0_0_ext_ram_rdata1[34] ,
    \data_arrays_0_0_ext_ram_rdata1[33] ,
    \data_arrays_0_0_ext_ram_rdata1[32] ,
    \data_arrays_0_0_ext_ram_rdata1[31] ,
    \data_arrays_0_0_ext_ram_rdata1[30] ,
    \data_arrays_0_0_ext_ram_rdata1[29] ,
    \data_arrays_0_0_ext_ram_rdata1[28] ,
    \data_arrays_0_0_ext_ram_rdata1[27] ,
    \data_arrays_0_0_ext_ram_rdata1[26] ,
    \data_arrays_0_0_ext_ram_rdata1[25] ,
    \data_arrays_0_0_ext_ram_rdata1[24] ,
    \data_arrays_0_0_ext_ram_rdata1[23] ,
    \data_arrays_0_0_ext_ram_rdata1[22] ,
    \data_arrays_0_0_ext_ram_rdata1[21] ,
    \data_arrays_0_0_ext_ram_rdata1[20] ,
    \data_arrays_0_0_ext_ram_rdata1[19] ,
    \data_arrays_0_0_ext_ram_rdata1[18] ,
    \data_arrays_0_0_ext_ram_rdata1[17] ,
    \data_arrays_0_0_ext_ram_rdata1[16] ,
    \data_arrays_0_0_ext_ram_rdata1[15] ,
    \data_arrays_0_0_ext_ram_rdata1[14] ,
    \data_arrays_0_0_ext_ram_rdata1[13] ,
    \data_arrays_0_0_ext_ram_rdata1[12] ,
    \data_arrays_0_0_ext_ram_rdata1[11] ,
    \data_arrays_0_0_ext_ram_rdata1[10] ,
    \data_arrays_0_0_ext_ram_rdata1[9] ,
    \data_arrays_0_0_ext_ram_rdata1[8] ,
    \data_arrays_0_0_ext_ram_rdata1[7] ,
    \data_arrays_0_0_ext_ram_rdata1[6] ,
    \data_arrays_0_0_ext_ram_rdata1[5] ,
    \data_arrays_0_0_ext_ram_rdata1[4] ,
    \data_arrays_0_0_ext_ram_rdata1[3] ,
    \data_arrays_0_0_ext_ram_rdata1[2] ,
    \data_arrays_0_0_ext_ram_rdata1[1] ,
    \data_arrays_0_0_ext_ram_rdata1[0] }),
    .data_arrays_0_0_ext_ram_rdata2({\data_arrays_0_0_ext_ram_rdata2[63] ,
    \data_arrays_0_0_ext_ram_rdata2[62] ,
    \data_arrays_0_0_ext_ram_rdata2[61] ,
    \data_arrays_0_0_ext_ram_rdata2[60] ,
    \data_arrays_0_0_ext_ram_rdata2[59] ,
    \data_arrays_0_0_ext_ram_rdata2[58] ,
    \data_arrays_0_0_ext_ram_rdata2[57] ,
    \data_arrays_0_0_ext_ram_rdata2[56] ,
    \data_arrays_0_0_ext_ram_rdata2[55] ,
    \data_arrays_0_0_ext_ram_rdata2[54] ,
    \data_arrays_0_0_ext_ram_rdata2[53] ,
    \data_arrays_0_0_ext_ram_rdata2[52] ,
    \data_arrays_0_0_ext_ram_rdata2[51] ,
    \data_arrays_0_0_ext_ram_rdata2[50] ,
    \data_arrays_0_0_ext_ram_rdata2[49] ,
    \data_arrays_0_0_ext_ram_rdata2[48] ,
    \data_arrays_0_0_ext_ram_rdata2[47] ,
    \data_arrays_0_0_ext_ram_rdata2[46] ,
    \data_arrays_0_0_ext_ram_rdata2[45] ,
    \data_arrays_0_0_ext_ram_rdata2[44] ,
    \data_arrays_0_0_ext_ram_rdata2[43] ,
    \data_arrays_0_0_ext_ram_rdata2[42] ,
    \data_arrays_0_0_ext_ram_rdata2[41] ,
    \data_arrays_0_0_ext_ram_rdata2[40] ,
    \data_arrays_0_0_ext_ram_rdata2[39] ,
    \data_arrays_0_0_ext_ram_rdata2[38] ,
    \data_arrays_0_0_ext_ram_rdata2[37] ,
    \data_arrays_0_0_ext_ram_rdata2[36] ,
    \data_arrays_0_0_ext_ram_rdata2[35] ,
    \data_arrays_0_0_ext_ram_rdata2[34] ,
    \data_arrays_0_0_ext_ram_rdata2[33] ,
    \data_arrays_0_0_ext_ram_rdata2[32] ,
    \data_arrays_0_0_ext_ram_rdata2[31] ,
    \data_arrays_0_0_ext_ram_rdata2[30] ,
    \data_arrays_0_0_ext_ram_rdata2[29] ,
    \data_arrays_0_0_ext_ram_rdata2[28] ,
    \data_arrays_0_0_ext_ram_rdata2[27] ,
    \data_arrays_0_0_ext_ram_rdata2[26] ,
    \data_arrays_0_0_ext_ram_rdata2[25] ,
    \data_arrays_0_0_ext_ram_rdata2[24] ,
    \data_arrays_0_0_ext_ram_rdata2[23] ,
    \data_arrays_0_0_ext_ram_rdata2[22] ,
    \data_arrays_0_0_ext_ram_rdata2[21] ,
    \data_arrays_0_0_ext_ram_rdata2[20] ,
    \data_arrays_0_0_ext_ram_rdata2[19] ,
    \data_arrays_0_0_ext_ram_rdata2[18] ,
    \data_arrays_0_0_ext_ram_rdata2[17] ,
    \data_arrays_0_0_ext_ram_rdata2[16] ,
    \data_arrays_0_0_ext_ram_rdata2[15] ,
    \data_arrays_0_0_ext_ram_rdata2[14] ,
    \data_arrays_0_0_ext_ram_rdata2[13] ,
    \data_arrays_0_0_ext_ram_rdata2[12] ,
    \data_arrays_0_0_ext_ram_rdata2[11] ,
    \data_arrays_0_0_ext_ram_rdata2[10] ,
    \data_arrays_0_0_ext_ram_rdata2[9] ,
    \data_arrays_0_0_ext_ram_rdata2[8] ,
    \data_arrays_0_0_ext_ram_rdata2[7] ,
    \data_arrays_0_0_ext_ram_rdata2[6] ,
    \data_arrays_0_0_ext_ram_rdata2[5] ,
    \data_arrays_0_0_ext_ram_rdata2[4] ,
    \data_arrays_0_0_ext_ram_rdata2[3] ,
    \data_arrays_0_0_ext_ram_rdata2[2] ,
    \data_arrays_0_0_ext_ram_rdata2[1] ,
    \data_arrays_0_0_ext_ram_rdata2[0] }),
    .data_arrays_0_0_ext_ram_rdata3({\data_arrays_0_0_ext_ram_rdata3[63] ,
    \data_arrays_0_0_ext_ram_rdata3[62] ,
    \data_arrays_0_0_ext_ram_rdata3[61] ,
    \data_arrays_0_0_ext_ram_rdata3[60] ,
    \data_arrays_0_0_ext_ram_rdata3[59] ,
    \data_arrays_0_0_ext_ram_rdata3[58] ,
    \data_arrays_0_0_ext_ram_rdata3[57] ,
    \data_arrays_0_0_ext_ram_rdata3[56] ,
    \data_arrays_0_0_ext_ram_rdata3[55] ,
    \data_arrays_0_0_ext_ram_rdata3[54] ,
    \data_arrays_0_0_ext_ram_rdata3[53] ,
    \data_arrays_0_0_ext_ram_rdata3[52] ,
    \data_arrays_0_0_ext_ram_rdata3[51] ,
    \data_arrays_0_0_ext_ram_rdata3[50] ,
    \data_arrays_0_0_ext_ram_rdata3[49] ,
    \data_arrays_0_0_ext_ram_rdata3[48] ,
    \data_arrays_0_0_ext_ram_rdata3[47] ,
    \data_arrays_0_0_ext_ram_rdata3[46] ,
    \data_arrays_0_0_ext_ram_rdata3[45] ,
    \data_arrays_0_0_ext_ram_rdata3[44] ,
    \data_arrays_0_0_ext_ram_rdata3[43] ,
    \data_arrays_0_0_ext_ram_rdata3[42] ,
    \data_arrays_0_0_ext_ram_rdata3[41] ,
    \data_arrays_0_0_ext_ram_rdata3[40] ,
    \data_arrays_0_0_ext_ram_rdata3[39] ,
    \data_arrays_0_0_ext_ram_rdata3[38] ,
    \data_arrays_0_0_ext_ram_rdata3[37] ,
    \data_arrays_0_0_ext_ram_rdata3[36] ,
    \data_arrays_0_0_ext_ram_rdata3[35] ,
    \data_arrays_0_0_ext_ram_rdata3[34] ,
    \data_arrays_0_0_ext_ram_rdata3[33] ,
    \data_arrays_0_0_ext_ram_rdata3[32] ,
    \data_arrays_0_0_ext_ram_rdata3[31] ,
    \data_arrays_0_0_ext_ram_rdata3[30] ,
    \data_arrays_0_0_ext_ram_rdata3[29] ,
    \data_arrays_0_0_ext_ram_rdata3[28] ,
    \data_arrays_0_0_ext_ram_rdata3[27] ,
    \data_arrays_0_0_ext_ram_rdata3[26] ,
    \data_arrays_0_0_ext_ram_rdata3[25] ,
    \data_arrays_0_0_ext_ram_rdata3[24] ,
    \data_arrays_0_0_ext_ram_rdata3[23] ,
    \data_arrays_0_0_ext_ram_rdata3[22] ,
    \data_arrays_0_0_ext_ram_rdata3[21] ,
    \data_arrays_0_0_ext_ram_rdata3[20] ,
    \data_arrays_0_0_ext_ram_rdata3[19] ,
    \data_arrays_0_0_ext_ram_rdata3[18] ,
    \data_arrays_0_0_ext_ram_rdata3[17] ,
    \data_arrays_0_0_ext_ram_rdata3[16] ,
    \data_arrays_0_0_ext_ram_rdata3[15] ,
    \data_arrays_0_0_ext_ram_rdata3[14] ,
    \data_arrays_0_0_ext_ram_rdata3[13] ,
    \data_arrays_0_0_ext_ram_rdata3[12] ,
    \data_arrays_0_0_ext_ram_rdata3[11] ,
    \data_arrays_0_0_ext_ram_rdata3[10] ,
    \data_arrays_0_0_ext_ram_rdata3[9] ,
    \data_arrays_0_0_ext_ram_rdata3[8] ,
    \data_arrays_0_0_ext_ram_rdata3[7] ,
    \data_arrays_0_0_ext_ram_rdata3[6] ,
    \data_arrays_0_0_ext_ram_rdata3[5] ,
    \data_arrays_0_0_ext_ram_rdata3[4] ,
    \data_arrays_0_0_ext_ram_rdata3[3] ,
    \data_arrays_0_0_ext_ram_rdata3[2] ,
    \data_arrays_0_0_ext_ram_rdata3[1] ,
    \data_arrays_0_0_ext_ram_rdata3[0] }),
    .data_arrays_0_0_ext_ram_wdata({\data_arrays_0_0_ext_ram_wdata[63] ,
    \data_arrays_0_0_ext_ram_wdata[62] ,
    \data_arrays_0_0_ext_ram_wdata[61] ,
    \data_arrays_0_0_ext_ram_wdata[60] ,
    \data_arrays_0_0_ext_ram_wdata[59] ,
    \data_arrays_0_0_ext_ram_wdata[58] ,
    \data_arrays_0_0_ext_ram_wdata[57] ,
    \data_arrays_0_0_ext_ram_wdata[56] ,
    \data_arrays_0_0_ext_ram_wdata[55] ,
    \data_arrays_0_0_ext_ram_wdata[54] ,
    \data_arrays_0_0_ext_ram_wdata[53] ,
    \data_arrays_0_0_ext_ram_wdata[52] ,
    \data_arrays_0_0_ext_ram_wdata[51] ,
    \data_arrays_0_0_ext_ram_wdata[50] ,
    \data_arrays_0_0_ext_ram_wdata[49] ,
    \data_arrays_0_0_ext_ram_wdata[48] ,
    \data_arrays_0_0_ext_ram_wdata[47] ,
    \data_arrays_0_0_ext_ram_wdata[46] ,
    \data_arrays_0_0_ext_ram_wdata[45] ,
    \data_arrays_0_0_ext_ram_wdata[44] ,
    \data_arrays_0_0_ext_ram_wdata[43] ,
    \data_arrays_0_0_ext_ram_wdata[42] ,
    \data_arrays_0_0_ext_ram_wdata[41] ,
    \data_arrays_0_0_ext_ram_wdata[40] ,
    \data_arrays_0_0_ext_ram_wdata[39] ,
    \data_arrays_0_0_ext_ram_wdata[38] ,
    \data_arrays_0_0_ext_ram_wdata[37] ,
    \data_arrays_0_0_ext_ram_wdata[36] ,
    \data_arrays_0_0_ext_ram_wdata[35] ,
    \data_arrays_0_0_ext_ram_wdata[34] ,
    \data_arrays_0_0_ext_ram_wdata[33] ,
    \data_arrays_0_0_ext_ram_wdata[32] ,
    \data_arrays_0_0_ext_ram_wdata[31] ,
    \data_arrays_0_0_ext_ram_wdata[30] ,
    \data_arrays_0_0_ext_ram_wdata[29] ,
    \data_arrays_0_0_ext_ram_wdata[28] ,
    \data_arrays_0_0_ext_ram_wdata[27] ,
    \data_arrays_0_0_ext_ram_wdata[26] ,
    \data_arrays_0_0_ext_ram_wdata[25] ,
    \data_arrays_0_0_ext_ram_wdata[24] ,
    \data_arrays_0_0_ext_ram_wdata[23] ,
    \data_arrays_0_0_ext_ram_wdata[22] ,
    \data_arrays_0_0_ext_ram_wdata[21] ,
    \data_arrays_0_0_ext_ram_wdata[20] ,
    \data_arrays_0_0_ext_ram_wdata[19] ,
    \data_arrays_0_0_ext_ram_wdata[18] ,
    \data_arrays_0_0_ext_ram_wdata[17] ,
    \data_arrays_0_0_ext_ram_wdata[16] ,
    \data_arrays_0_0_ext_ram_wdata[15] ,
    \data_arrays_0_0_ext_ram_wdata[14] ,
    \data_arrays_0_0_ext_ram_wdata[13] ,
    \data_arrays_0_0_ext_ram_wdata[12] ,
    \data_arrays_0_0_ext_ram_wdata[11] ,
    \data_arrays_0_0_ext_ram_wdata[10] ,
    \data_arrays_0_0_ext_ram_wdata[9] ,
    \data_arrays_0_0_ext_ram_wdata[8] ,
    \data_arrays_0_0_ext_ram_wdata[7] ,
    \data_arrays_0_0_ext_ram_wdata[6] ,
    \data_arrays_0_0_ext_ram_wdata[5] ,
    \data_arrays_0_0_ext_ram_wdata[4] ,
    \data_arrays_0_0_ext_ram_wdata[3] ,
    \data_arrays_0_0_ext_ram_wdata[2] ,
    \data_arrays_0_0_ext_ram_wdata[1] ,
    \data_arrays_0_0_ext_ram_wdata[0] }),
    .data_arrays_0_0_ext_ram_wmask({\data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[0] }),
    .io_in({io_in[37],
    io_in[36],
    io_in[35],
    io_in[34],
    io_in[33],
    io_in[32],
    io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21],
    io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6],
    io_in[5],
    io_in[4],
    io_in[3],
    io_in[2],
    io_in[1],
    io_in[0]}),
    .io_oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .io_out({io_out[37],
    io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8],
    io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .irq({user_irq[2],
    user_irq[1],
    user_irq[0]}),
    .la_data_in({la_data_in[127],
    la_data_in[126],
    la_data_in[125],
    la_data_in[124],
    la_data_in[123],
    la_data_in[122],
    la_data_in[121],
    la_data_in[120],
    la_data_in[119],
    la_data_in[118],
    la_data_in[117],
    la_data_in[116],
    la_data_in[115],
    la_data_in[114],
    la_data_in[113],
    la_data_in[112],
    la_data_in[111],
    la_data_in[110],
    la_data_in[109],
    la_data_in[108],
    la_data_in[107],
    la_data_in[106],
    la_data_in[105],
    la_data_in[104],
    la_data_in[103],
    la_data_in[102],
    la_data_in[101],
    la_data_in[100],
    la_data_in[99],
    la_data_in[98],
    la_data_in[97],
    la_data_in[96],
    la_data_in[95],
    la_data_in[94],
    la_data_in[93],
    la_data_in[92],
    la_data_in[91],
    la_data_in[90],
    la_data_in[89],
    la_data_in[88],
    la_data_in[87],
    la_data_in[86],
    la_data_in[85],
    la_data_in[84],
    la_data_in[83],
    la_data_in[82],
    la_data_in[81],
    la_data_in[80],
    la_data_in[79],
    la_data_in[78],
    la_data_in[77],
    la_data_in[76],
    la_data_in[75],
    la_data_in[74],
    la_data_in[73],
    la_data_in[72],
    la_data_in[71],
    la_data_in[70],
    la_data_in[69],
    la_data_in[68],
    la_data_in[67],
    la_data_in[66],
    la_data_in[65],
    la_data_in[64],
    la_data_in[63],
    la_data_in[62],
    la_data_in[61],
    la_data_in[60],
    la_data_in[59],
    la_data_in[58],
    la_data_in[57],
    la_data_in[56],
    la_data_in[55],
    la_data_in[54],
    la_data_in[53],
    la_data_in[52],
    la_data_in[51],
    la_data_in[50],
    la_data_in[49],
    la_data_in[48],
    la_data_in[47],
    la_data_in[46],
    la_data_in[45],
    la_data_in[44],
    la_data_in[43],
    la_data_in[42],
    la_data_in[41],
    la_data_in[40],
    la_data_in[39],
    la_data_in[38],
    la_data_in[37],
    la_data_in[36],
    la_data_in[35],
    la_data_in[34],
    la_data_in[33],
    la_data_in[32],
    la_data_in[31],
    la_data_in[30],
    la_data_in[29],
    la_data_in[28],
    la_data_in[27],
    la_data_in[26],
    la_data_in[25],
    la_data_in[24],
    la_data_in[23],
    la_data_in[22],
    la_data_in[21],
    la_data_in[20],
    la_data_in[19],
    la_data_in[18],
    la_data_in[17],
    la_data_in[16],
    la_data_in[15],
    la_data_in[14],
    la_data_in[13],
    la_data_in[12],
    la_data_in[11],
    la_data_in[10],
    la_data_in[9],
    la_data_in[8],
    la_data_in[7],
    la_data_in[6],
    la_data_in[5],
    la_data_in[4],
    la_data_in[3],
    la_data_in[2],
    la_data_in[1],
    la_data_in[0]}),
    .la_data_out({la_data_out[127],
    la_data_out[126],
    la_data_out[125],
    la_data_out[124],
    la_data_out[123],
    la_data_out[122],
    la_data_out[121],
    la_data_out[120],
    la_data_out[119],
    la_data_out[118],
    la_data_out[117],
    la_data_out[116],
    la_data_out[115],
    la_data_out[114],
    la_data_out[113],
    la_data_out[112],
    la_data_out[111],
    la_data_out[110],
    la_data_out[109],
    la_data_out[108],
    la_data_out[107],
    la_data_out[106],
    la_data_out[105],
    la_data_out[104],
    la_data_out[103],
    la_data_out[102],
    la_data_out[101],
    la_data_out[100],
    la_data_out[99],
    la_data_out[98],
    la_data_out[97],
    la_data_out[96],
    la_data_out[95],
    la_data_out[94],
    la_data_out[93],
    la_data_out[92],
    la_data_out[91],
    la_data_out[90],
    la_data_out[89],
    la_data_out[88],
    la_data_out[87],
    la_data_out[86],
    la_data_out[85],
    la_data_out[84],
    la_data_out[83],
    la_data_out[82],
    la_data_out[81],
    la_data_out[80],
    la_data_out[79],
    la_data_out[78],
    la_data_out[77],
    la_data_out[76],
    la_data_out[75],
    la_data_out[74],
    la_data_out[73],
    la_data_out[72],
    la_data_out[71],
    la_data_out[70],
    la_data_out[69],
    la_data_out[68],
    la_data_out[67],
    la_data_out[66],
    la_data_out[65],
    la_data_out[64],
    la_data_out[63],
    la_data_out[62],
    la_data_out[61],
    la_data_out[60],
    la_data_out[59],
    la_data_out[58],
    la_data_out[57],
    la_data_out[56],
    la_data_out[55],
    la_data_out[54],
    la_data_out[53],
    la_data_out[52],
    la_data_out[51],
    la_data_out[50],
    la_data_out[49],
    la_data_out[48],
    la_data_out[47],
    la_data_out[46],
    la_data_out[45],
    la_data_out[44],
    la_data_out[43],
    la_data_out[42],
    la_data_out[41],
    la_data_out[40],
    la_data_out[39],
    la_data_out[38],
    la_data_out[37],
    la_data_out[36],
    la_data_out[35],
    la_data_out[34],
    la_data_out[33],
    la_data_out[32],
    la_data_out[31],
    la_data_out[30],
    la_data_out[29],
    la_data_out[28],
    la_data_out[27],
    la_data_out[26],
    la_data_out[25],
    la_data_out[24],
    la_data_out[23],
    la_data_out[22],
    la_data_out[21],
    la_data_out[20],
    la_data_out[19],
    la_data_out[18],
    la_data_out[17],
    la_data_out[16],
    la_data_out[15],
    la_data_out[14],
    la_data_out[13],
    la_data_out[12],
    la_data_out[11],
    la_data_out[10],
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0]}),
    .la_oenb({la_oenb[127],
    la_oenb[126],
    la_oenb[125],
    la_oenb[124],
    la_oenb[123],
    la_oenb[122],
    la_oenb[121],
    la_oenb[120],
    la_oenb[119],
    la_oenb[118],
    la_oenb[117],
    la_oenb[116],
    la_oenb[115],
    la_oenb[114],
    la_oenb[113],
    la_oenb[112],
    la_oenb[111],
    la_oenb[110],
    la_oenb[109],
    la_oenb[108],
    la_oenb[107],
    la_oenb[106],
    la_oenb[105],
    la_oenb[104],
    la_oenb[103],
    la_oenb[102],
    la_oenb[101],
    la_oenb[100],
    la_oenb[99],
    la_oenb[98],
    la_oenb[97],
    la_oenb[96],
    la_oenb[95],
    la_oenb[94],
    la_oenb[93],
    la_oenb[92],
    la_oenb[91],
    la_oenb[90],
    la_oenb[89],
    la_oenb[88],
    la_oenb[87],
    la_oenb[86],
    la_oenb[85],
    la_oenb[84],
    la_oenb[83],
    la_oenb[82],
    la_oenb[81],
    la_oenb[80],
    la_oenb[79],
    la_oenb[78],
    la_oenb[77],
    la_oenb[76],
    la_oenb[75],
    la_oenb[74],
    la_oenb[73],
    la_oenb[72],
    la_oenb[71],
    la_oenb[70],
    la_oenb[69],
    la_oenb[68],
    la_oenb[67],
    la_oenb[66],
    la_oenb[65],
    la_oenb[64],
    la_oenb[63],
    la_oenb[62],
    la_oenb[61],
    la_oenb[60],
    la_oenb[59],
    la_oenb[58],
    la_oenb[57],
    la_oenb[56],
    la_oenb[55],
    la_oenb[54],
    la_oenb[53],
    la_oenb[52],
    la_oenb[51],
    la_oenb[50],
    la_oenb[49],
    la_oenb[48],
    la_oenb[47],
    la_oenb[46],
    la_oenb[45],
    la_oenb[44],
    la_oenb[43],
    la_oenb[42],
    la_oenb[41],
    la_oenb[40],
    la_oenb[39],
    la_oenb[38],
    la_oenb[37],
    la_oenb[36],
    la_oenb[35],
    la_oenb[34],
    la_oenb[33],
    la_oenb[32],
    la_oenb[31],
    la_oenb[30],
    la_oenb[29],
    la_oenb[28],
    la_oenb[27],
    la_oenb[26],
    la_oenb[25],
    la_oenb[24],
    la_oenb[23],
    la_oenb[22],
    la_oenb[21],
    la_oenb[20],
    la_oenb[19],
    la_oenb[18],
    la_oenb[17],
    la_oenb[16],
    la_oenb[15],
    la_oenb[14],
    la_oenb[13],
    la_oenb[12],
    la_oenb[11],
    la_oenb[10],
    la_oenb[9],
    la_oenb[8],
    la_oenb[7],
    la_oenb[6],
    la_oenb[5],
    la_oenb[4],
    la_oenb[3],
    la_oenb[2],
    la_oenb[1],
    la_oenb[0]}),
    .ram_clk_delay_sel({\ram_clk_delay_sel[31] ,
    \ram_clk_delay_sel[30] ,
    \ram_clk_delay_sel[29] ,
    \ram_clk_delay_sel[28] ,
    \ram_clk_delay_sel[27] ,
    \ram_clk_delay_sel[26] ,
    \ram_clk_delay_sel[25] ,
    \ram_clk_delay_sel[24] ,
    \ram_clk_delay_sel[23] ,
    \ram_clk_delay_sel[22] ,
    \ram_clk_delay_sel[21] ,
    \ram_clk_delay_sel[20] ,
    \ram_clk_delay_sel[19] ,
    \ram_clk_delay_sel[18] ,
    \ram_clk_delay_sel[17] ,
    \ram_clk_delay_sel[16] ,
    \ram_clk_delay_sel[15] ,
    \ram_clk_delay_sel[14] ,
    \ram_clk_delay_sel[13] ,
    \ram_clk_delay_sel[12] ,
    \ram_clk_delay_sel[11] ,
    \ram_clk_delay_sel[10] ,
    \ram_clk_delay_sel[9] ,
    \ram_clk_delay_sel[8] ,
    \ram_clk_delay_sel[7] ,
    \ram_clk_delay_sel[6] ,
    \ram_clk_delay_sel[5] ,
    \ram_clk_delay_sel[4] ,
    \ram_clk_delay_sel[3] ,
    \ram_clk_delay_sel[2] ,
    \ram_clk_delay_sel[1] ,
    \ram_clk_delay_sel[0] }),
    .tag_array_ext_ram_addr({\tag_array_ext_ram_addr[7] ,
    \tag_array_ext_ram_addr[6] ,
    \tag_array_ext_ram_addr[5] ,
    \tag_array_ext_ram_addr[4] ,
    \tag_array_ext_ram_addr[3] ,
    \tag_array_ext_ram_addr[2] ,
    \tag_array_ext_ram_addr[1] ,
    \tag_array_ext_ram_addr[0] }),
    .tag_array_ext_ram_addr1({\tag_array_ext_ram_addr1[7] ,
    \tag_array_ext_ram_addr1[6] ,
    \tag_array_ext_ram_addr1[5] ,
    \tag_array_ext_ram_addr1[4] ,
    \tag_array_ext_ram_addr1[3] ,
    \tag_array_ext_ram_addr1[2] ,
    \tag_array_ext_ram_addr1[1] ,
    \tag_array_ext_ram_addr1[0] }),
    .tag_array_ext_ram_csb1({\tag_array_ext_ram_csb1[1] ,
    \tag_array_ext_ram_csb1[0] }),
    .tag_array_ext_ram_rdata0({\tag_array_ext_ram_rdata0[31] ,
    \tag_array_ext_ram_rdata0[30] ,
    \tag_array_ext_ram_rdata0[29] ,
    \tag_array_ext_ram_rdata0[28] ,
    \tag_array_ext_ram_rdata0[27] ,
    \tag_array_ext_ram_rdata0[26] ,
    \tag_array_ext_ram_rdata0[25] ,
    \tag_array_ext_ram_rdata0[24] ,
    \tag_array_ext_ram_rdata0[23] ,
    \tag_array_ext_ram_rdata0[22] ,
    \tag_array_ext_ram_rdata0[21] ,
    \tag_array_ext_ram_rdata0[20] ,
    \tag_array_ext_ram_rdata0[19] ,
    \tag_array_ext_ram_rdata0[18] ,
    \tag_array_ext_ram_rdata0[17] ,
    \tag_array_ext_ram_rdata0[16] ,
    \tag_array_ext_ram_rdata0[15] ,
    \tag_array_ext_ram_rdata0[14] ,
    \tag_array_ext_ram_rdata0[13] ,
    \tag_array_ext_ram_rdata0[12] ,
    \tag_array_ext_ram_rdata0[11] ,
    \tag_array_ext_ram_rdata0[10] ,
    \tag_array_ext_ram_rdata0[9] ,
    \tag_array_ext_ram_rdata0[8] ,
    \tag_array_ext_ram_rdata0[7] ,
    \tag_array_ext_ram_rdata0[6] ,
    \tag_array_ext_ram_rdata0[5] ,
    \tag_array_ext_ram_rdata0[4] ,
    \tag_array_ext_ram_rdata0[3] ,
    \tag_array_ext_ram_rdata0[2] ,
    \tag_array_ext_ram_rdata0[1] ,
    \tag_array_ext_ram_rdata0[0] }),
    .tag_array_ext_ram_rdata1({\tag_array_ext_ram_rdata1[31] ,
    \tag_array_ext_ram_rdata1[30] ,
    \tag_array_ext_ram_rdata1[29] ,
    \tag_array_ext_ram_rdata1[28] ,
    \tag_array_ext_ram_rdata1[27] ,
    \tag_array_ext_ram_rdata1[26] ,
    \tag_array_ext_ram_rdata1[25] ,
    \tag_array_ext_ram_rdata1[24] ,
    \tag_array_ext_ram_rdata1[23] ,
    \tag_array_ext_ram_rdata1[22] ,
    \tag_array_ext_ram_rdata1[21] ,
    \tag_array_ext_ram_rdata1[20] ,
    \tag_array_ext_ram_rdata1[19] ,
    \tag_array_ext_ram_rdata1[18] ,
    \tag_array_ext_ram_rdata1[17] ,
    \tag_array_ext_ram_rdata1[16] ,
    \tag_array_ext_ram_rdata1[15] ,
    \tag_array_ext_ram_rdata1[14] ,
    \tag_array_ext_ram_rdata1[13] ,
    \tag_array_ext_ram_rdata1[12] ,
    \tag_array_ext_ram_rdata1[11] ,
    \tag_array_ext_ram_rdata1[10] ,
    \tag_array_ext_ram_rdata1[9] ,
    \tag_array_ext_ram_rdata1[8] ,
    \tag_array_ext_ram_rdata1[7] ,
    \tag_array_ext_ram_rdata1[6] ,
    \tag_array_ext_ram_rdata1[5] ,
    \tag_array_ext_ram_rdata1[4] ,
    \tag_array_ext_ram_rdata1[3] ,
    \tag_array_ext_ram_rdata1[2] ,
    \tag_array_ext_ram_rdata1[1] ,
    \tag_array_ext_ram_rdata1[0] }),
    .tag_array_ext_ram_wdata({\tag_array_ext_ram_wdata[63] ,
    \tag_array_ext_ram_wdata[62] ,
    \tag_array_ext_ram_wdata[61] ,
    \tag_array_ext_ram_wdata[60] ,
    \tag_array_ext_ram_wdata[59] ,
    \tag_array_ext_ram_wdata[58] ,
    \tag_array_ext_ram_wdata[57] ,
    \tag_array_ext_ram_wdata[56] ,
    \tag_array_ext_ram_wdata[55] ,
    \tag_array_ext_ram_wdata[54] ,
    \tag_array_ext_ram_wdata[53] ,
    \tag_array_ext_ram_wdata[52] ,
    \tag_array_ext_ram_wdata[51] ,
    \tag_array_ext_ram_wdata[50] ,
    \tag_array_ext_ram_wdata[49] ,
    \tag_array_ext_ram_wdata[48] ,
    \tag_array_ext_ram_wdata[47] ,
    \tag_array_ext_ram_wdata[46] ,
    \tag_array_ext_ram_wdata[45] ,
    \tag_array_ext_ram_wdata[44] ,
    \tag_array_ext_ram_wdata[43] ,
    \tag_array_ext_ram_wdata[42] ,
    \tag_array_ext_ram_wdata[41] ,
    \tag_array_ext_ram_wdata[40] ,
    \tag_array_ext_ram_wdata[39] ,
    \tag_array_ext_ram_wdata[38] ,
    \tag_array_ext_ram_wdata[37] ,
    \tag_array_ext_ram_wdata[36] ,
    \tag_array_ext_ram_wdata[35] ,
    \tag_array_ext_ram_wdata[34] ,
    \tag_array_ext_ram_wdata[33] ,
    \tag_array_ext_ram_wdata[32] ,
    \tag_array_ext_ram_wdata[31] ,
    \tag_array_ext_ram_wdata[30] ,
    \tag_array_ext_ram_wdata[29] ,
    \tag_array_ext_ram_wdata[28] ,
    \tag_array_ext_ram_wdata[27] ,
    \tag_array_ext_ram_wdata[26] ,
    \tag_array_ext_ram_wdata[25] ,
    \tag_array_ext_ram_wdata[24] ,
    \tag_array_ext_ram_wdata[23] ,
    \tag_array_ext_ram_wdata[22] ,
    \tag_array_ext_ram_wdata[21] ,
    \tag_array_ext_ram_wdata[20] ,
    \tag_array_ext_ram_wdata[19] ,
    \tag_array_ext_ram_wdata[18] ,
    \tag_array_ext_ram_wdata[17] ,
    \tag_array_ext_ram_wdata[16] ,
    \tag_array_ext_ram_wdata[15] ,
    \tag_array_ext_ram_wdata[14] ,
    \tag_array_ext_ram_wdata[13] ,
    \tag_array_ext_ram_wdata[12] ,
    \tag_array_ext_ram_wdata[11] ,
    \tag_array_ext_ram_wdata[10] ,
    \tag_array_ext_ram_wdata[9] ,
    \tag_array_ext_ram_wdata[8] ,
    \tag_array_ext_ram_wdata[7] ,
    \tag_array_ext_ram_wdata[6] ,
    \tag_array_ext_ram_wdata[5] ,
    \tag_array_ext_ram_wdata[4] ,
    \tag_array_ext_ram_wdata[3] ,
    \tag_array_ext_ram_wdata[2] ,
    \tag_array_ext_ram_wdata[1] ,
    \tag_array_ext_ram_wdata[0] }),
    .tag_array_ext_ram_wmask({\tag_array_ext_ram_wmask[1] ,
    \tag_array_ext_ram_wmask[0] }),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 sky130_sram_2kbyte_1rw1r_32x512_8 data_arrays_0_0_ext_ram0h (.csb0(\data_arrays_0_0_ext_ram_csb[0] ),
    .csb1(\data_arrays_0_0_ext_ram_csb1[0] ),
    .web0(data_arrays_0_0_ext_ram_web),
    .clk0(data_arrays_0_0_ext_ram_clk0),
    .clk1(data_arrays_0_0_ext_ram_clk0),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\data_arrays_0_0_ext_ram_addr[8] ,
    \data_arrays_0_0_ext_ram_addr[7] ,
    \data_arrays_0_0_ext_ram_addr[6] ,
    \data_arrays_0_0_ext_ram_addr[5] ,
    \data_arrays_0_0_ext_ram_addr[4] ,
    \data_arrays_0_0_ext_ram_addr[3] ,
    \data_arrays_0_0_ext_ram_addr[2] ,
    \data_arrays_0_0_ext_ram_addr[1] ,
    \data_arrays_0_0_ext_ram_addr[0] }),
    .addr1({\data_arrays_0_0_ext_ram_addr1[8] ,
    \data_arrays_0_0_ext_ram_addr1[7] ,
    \data_arrays_0_0_ext_ram_addr1[6] ,
    \data_arrays_0_0_ext_ram_addr1[5] ,
    \data_arrays_0_0_ext_ram_addr1[4] ,
    \data_arrays_0_0_ext_ram_addr1[3] ,
    \data_arrays_0_0_ext_ram_addr1[2] ,
    \data_arrays_0_0_ext_ram_addr1[1] ,
    \data_arrays_0_0_ext_ram_addr1[0] }),
    .din0({\data_arrays_0_0_ext_ram_wdata[63] ,
    \data_arrays_0_0_ext_ram_wdata[62] ,
    \data_arrays_0_0_ext_ram_wdata[61] ,
    \data_arrays_0_0_ext_ram_wdata[60] ,
    \data_arrays_0_0_ext_ram_wdata[59] ,
    \data_arrays_0_0_ext_ram_wdata[58] ,
    \data_arrays_0_0_ext_ram_wdata[57] ,
    \data_arrays_0_0_ext_ram_wdata[56] ,
    \data_arrays_0_0_ext_ram_wdata[55] ,
    \data_arrays_0_0_ext_ram_wdata[54] ,
    \data_arrays_0_0_ext_ram_wdata[53] ,
    \data_arrays_0_0_ext_ram_wdata[52] ,
    \data_arrays_0_0_ext_ram_wdata[51] ,
    \data_arrays_0_0_ext_ram_wdata[50] ,
    \data_arrays_0_0_ext_ram_wdata[49] ,
    \data_arrays_0_0_ext_ram_wdata[48] ,
    \data_arrays_0_0_ext_ram_wdata[47] ,
    \data_arrays_0_0_ext_ram_wdata[46] ,
    \data_arrays_0_0_ext_ram_wdata[45] ,
    \data_arrays_0_0_ext_ram_wdata[44] ,
    \data_arrays_0_0_ext_ram_wdata[43] ,
    \data_arrays_0_0_ext_ram_wdata[42] ,
    \data_arrays_0_0_ext_ram_wdata[41] ,
    \data_arrays_0_0_ext_ram_wdata[40] ,
    \data_arrays_0_0_ext_ram_wdata[39] ,
    \data_arrays_0_0_ext_ram_wdata[38] ,
    \data_arrays_0_0_ext_ram_wdata[37] ,
    \data_arrays_0_0_ext_ram_wdata[36] ,
    \data_arrays_0_0_ext_ram_wdata[35] ,
    \data_arrays_0_0_ext_ram_wdata[34] ,
    \data_arrays_0_0_ext_ram_wdata[33] ,
    \data_arrays_0_0_ext_ram_wdata[32] }),
    .dout0({\data_arrays_0_0_ext_ram_rdata0[63] ,
    \data_arrays_0_0_ext_ram_rdata0[62] ,
    \data_arrays_0_0_ext_ram_rdata0[61] ,
    \data_arrays_0_0_ext_ram_rdata0[60] ,
    \data_arrays_0_0_ext_ram_rdata0[59] ,
    \data_arrays_0_0_ext_ram_rdata0[58] ,
    \data_arrays_0_0_ext_ram_rdata0[57] ,
    \data_arrays_0_0_ext_ram_rdata0[56] ,
    \data_arrays_0_0_ext_ram_rdata0[55] ,
    \data_arrays_0_0_ext_ram_rdata0[54] ,
    \data_arrays_0_0_ext_ram_rdata0[53] ,
    \data_arrays_0_0_ext_ram_rdata0[52] ,
    \data_arrays_0_0_ext_ram_rdata0[51] ,
    \data_arrays_0_0_ext_ram_rdata0[50] ,
    \data_arrays_0_0_ext_ram_rdata0[49] ,
    \data_arrays_0_0_ext_ram_rdata0[48] ,
    \data_arrays_0_0_ext_ram_rdata0[47] ,
    \data_arrays_0_0_ext_ram_rdata0[46] ,
    \data_arrays_0_0_ext_ram_rdata0[45] ,
    \data_arrays_0_0_ext_ram_rdata0[44] ,
    \data_arrays_0_0_ext_ram_rdata0[43] ,
    \data_arrays_0_0_ext_ram_rdata0[42] ,
    \data_arrays_0_0_ext_ram_rdata0[41] ,
    \data_arrays_0_0_ext_ram_rdata0[40] ,
    \data_arrays_0_0_ext_ram_rdata0[39] ,
    \data_arrays_0_0_ext_ram_rdata0[38] ,
    \data_arrays_0_0_ext_ram_rdata0[37] ,
    \data_arrays_0_0_ext_ram_rdata0[36] ,
    \data_arrays_0_0_ext_ram_rdata0[35] ,
    \data_arrays_0_0_ext_ram_rdata0[34] ,
    \data_arrays_0_0_ext_ram_rdata0[33] ,
    \data_arrays_0_0_ext_ram_rdata0[32] }),
    .dout1({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .wmask0({\data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 data_arrays_0_0_ext_ram0l (.csb0(\data_arrays_0_0_ext_ram_csb[0] ),
    .csb1(\data_arrays_0_0_ext_ram_csb1[1] ),
    .web0(data_arrays_0_0_ext_ram_web),
    .clk0(data_arrays_0_0_ext_ram_clk0),
    .clk1(data_arrays_0_0_ext_ram_clk0),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\data_arrays_0_0_ext_ram_addr[8] ,
    \data_arrays_0_0_ext_ram_addr[7] ,
    \data_arrays_0_0_ext_ram_addr[6] ,
    \data_arrays_0_0_ext_ram_addr[5] ,
    \data_arrays_0_0_ext_ram_addr[4] ,
    \data_arrays_0_0_ext_ram_addr[3] ,
    \data_arrays_0_0_ext_ram_addr[2] ,
    \data_arrays_0_0_ext_ram_addr[1] ,
    \data_arrays_0_0_ext_ram_addr[0] }),
    .addr1({\data_arrays_0_0_ext_ram_addr1[8] ,
    \data_arrays_0_0_ext_ram_addr1[7] ,
    \data_arrays_0_0_ext_ram_addr1[6] ,
    \data_arrays_0_0_ext_ram_addr1[5] ,
    \data_arrays_0_0_ext_ram_addr1[4] ,
    \data_arrays_0_0_ext_ram_addr1[3] ,
    \data_arrays_0_0_ext_ram_addr1[2] ,
    \data_arrays_0_0_ext_ram_addr1[1] ,
    \data_arrays_0_0_ext_ram_addr1[0] }),
    .din0({\data_arrays_0_0_ext_ram_wdata[31] ,
    \data_arrays_0_0_ext_ram_wdata[30] ,
    \data_arrays_0_0_ext_ram_wdata[29] ,
    \data_arrays_0_0_ext_ram_wdata[28] ,
    \data_arrays_0_0_ext_ram_wdata[27] ,
    \data_arrays_0_0_ext_ram_wdata[26] ,
    \data_arrays_0_0_ext_ram_wdata[25] ,
    \data_arrays_0_0_ext_ram_wdata[24] ,
    \data_arrays_0_0_ext_ram_wdata[23] ,
    \data_arrays_0_0_ext_ram_wdata[22] ,
    \data_arrays_0_0_ext_ram_wdata[21] ,
    \data_arrays_0_0_ext_ram_wdata[20] ,
    \data_arrays_0_0_ext_ram_wdata[19] ,
    \data_arrays_0_0_ext_ram_wdata[18] ,
    \data_arrays_0_0_ext_ram_wdata[17] ,
    \data_arrays_0_0_ext_ram_wdata[16] ,
    \data_arrays_0_0_ext_ram_wdata[15] ,
    \data_arrays_0_0_ext_ram_wdata[14] ,
    \data_arrays_0_0_ext_ram_wdata[13] ,
    \data_arrays_0_0_ext_ram_wdata[12] ,
    \data_arrays_0_0_ext_ram_wdata[11] ,
    \data_arrays_0_0_ext_ram_wdata[10] ,
    \data_arrays_0_0_ext_ram_wdata[9] ,
    \data_arrays_0_0_ext_ram_wdata[8] ,
    \data_arrays_0_0_ext_ram_wdata[7] ,
    \data_arrays_0_0_ext_ram_wdata[6] ,
    \data_arrays_0_0_ext_ram_wdata[5] ,
    \data_arrays_0_0_ext_ram_wdata[4] ,
    \data_arrays_0_0_ext_ram_wdata[3] ,
    \data_arrays_0_0_ext_ram_wdata[2] ,
    \data_arrays_0_0_ext_ram_wdata[1] ,
    \data_arrays_0_0_ext_ram_wdata[0] }),
    .dout0({\data_arrays_0_0_ext_ram_rdata0[31] ,
    \data_arrays_0_0_ext_ram_rdata0[30] ,
    \data_arrays_0_0_ext_ram_rdata0[29] ,
    \data_arrays_0_0_ext_ram_rdata0[28] ,
    \data_arrays_0_0_ext_ram_rdata0[27] ,
    \data_arrays_0_0_ext_ram_rdata0[26] ,
    \data_arrays_0_0_ext_ram_rdata0[25] ,
    \data_arrays_0_0_ext_ram_rdata0[24] ,
    \data_arrays_0_0_ext_ram_rdata0[23] ,
    \data_arrays_0_0_ext_ram_rdata0[22] ,
    \data_arrays_0_0_ext_ram_rdata0[21] ,
    \data_arrays_0_0_ext_ram_rdata0[20] ,
    \data_arrays_0_0_ext_ram_rdata0[19] ,
    \data_arrays_0_0_ext_ram_rdata0[18] ,
    \data_arrays_0_0_ext_ram_rdata0[17] ,
    \data_arrays_0_0_ext_ram_rdata0[16] ,
    \data_arrays_0_0_ext_ram_rdata0[15] ,
    \data_arrays_0_0_ext_ram_rdata0[14] ,
    \data_arrays_0_0_ext_ram_rdata0[13] ,
    \data_arrays_0_0_ext_ram_rdata0[12] ,
    \data_arrays_0_0_ext_ram_rdata0[11] ,
    \data_arrays_0_0_ext_ram_rdata0[10] ,
    \data_arrays_0_0_ext_ram_rdata0[9] ,
    \data_arrays_0_0_ext_ram_rdata0[8] ,
    \data_arrays_0_0_ext_ram_rdata0[7] ,
    \data_arrays_0_0_ext_ram_rdata0[6] ,
    \data_arrays_0_0_ext_ram_rdata0[5] ,
    \data_arrays_0_0_ext_ram_rdata0[4] ,
    \data_arrays_0_0_ext_ram_rdata0[3] ,
    \data_arrays_0_0_ext_ram_rdata0[2] ,
    \data_arrays_0_0_ext_ram_rdata0[1] ,
    \data_arrays_0_0_ext_ram_rdata0[0] }),
    .dout1({_NC33,
    _NC34,
    _NC35,
    _NC36,
    _NC37,
    _NC38,
    _NC39,
    _NC40,
    _NC41,
    _NC42,
    _NC43,
    _NC44,
    _NC45,
    _NC46,
    _NC47,
    _NC48,
    _NC49,
    _NC50,
    _NC51,
    _NC52,
    _NC53,
    _NC54,
    _NC55,
    _NC56,
    _NC57,
    _NC58,
    _NC59,
    _NC60,
    _NC61,
    _NC62,
    _NC63,
    _NC64}),
    .wmask0({\data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 data_arrays_0_0_ext_ram1h (.csb0(\data_arrays_0_0_ext_ram_csb[1] ),
    .csb1(\data_arrays_0_0_ext_ram_csb1[2] ),
    .web0(data_arrays_0_0_ext_ram_web),
    .clk0(data_arrays_0_0_ext_ram_clk1),
    .clk1(data_arrays_0_0_ext_ram_clk1),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\data_arrays_0_0_ext_ram_addr[8] ,
    \data_arrays_0_0_ext_ram_addr[7] ,
    \data_arrays_0_0_ext_ram_addr[6] ,
    \data_arrays_0_0_ext_ram_addr[5] ,
    \data_arrays_0_0_ext_ram_addr[4] ,
    \data_arrays_0_0_ext_ram_addr[3] ,
    \data_arrays_0_0_ext_ram_addr[2] ,
    \data_arrays_0_0_ext_ram_addr[1] ,
    \data_arrays_0_0_ext_ram_addr[0] }),
    .addr1({\data_arrays_0_0_ext_ram_addr1[8] ,
    \data_arrays_0_0_ext_ram_addr1[7] ,
    \data_arrays_0_0_ext_ram_addr1[6] ,
    \data_arrays_0_0_ext_ram_addr1[5] ,
    \data_arrays_0_0_ext_ram_addr1[4] ,
    \data_arrays_0_0_ext_ram_addr1[3] ,
    \data_arrays_0_0_ext_ram_addr1[2] ,
    \data_arrays_0_0_ext_ram_addr1[1] ,
    \data_arrays_0_0_ext_ram_addr1[0] }),
    .din0({\data_arrays_0_0_ext_ram_wdata[63] ,
    \data_arrays_0_0_ext_ram_wdata[62] ,
    \data_arrays_0_0_ext_ram_wdata[61] ,
    \data_arrays_0_0_ext_ram_wdata[60] ,
    \data_arrays_0_0_ext_ram_wdata[59] ,
    \data_arrays_0_0_ext_ram_wdata[58] ,
    \data_arrays_0_0_ext_ram_wdata[57] ,
    \data_arrays_0_0_ext_ram_wdata[56] ,
    \data_arrays_0_0_ext_ram_wdata[55] ,
    \data_arrays_0_0_ext_ram_wdata[54] ,
    \data_arrays_0_0_ext_ram_wdata[53] ,
    \data_arrays_0_0_ext_ram_wdata[52] ,
    \data_arrays_0_0_ext_ram_wdata[51] ,
    \data_arrays_0_0_ext_ram_wdata[50] ,
    \data_arrays_0_0_ext_ram_wdata[49] ,
    \data_arrays_0_0_ext_ram_wdata[48] ,
    \data_arrays_0_0_ext_ram_wdata[47] ,
    \data_arrays_0_0_ext_ram_wdata[46] ,
    \data_arrays_0_0_ext_ram_wdata[45] ,
    \data_arrays_0_0_ext_ram_wdata[44] ,
    \data_arrays_0_0_ext_ram_wdata[43] ,
    \data_arrays_0_0_ext_ram_wdata[42] ,
    \data_arrays_0_0_ext_ram_wdata[41] ,
    \data_arrays_0_0_ext_ram_wdata[40] ,
    \data_arrays_0_0_ext_ram_wdata[39] ,
    \data_arrays_0_0_ext_ram_wdata[38] ,
    \data_arrays_0_0_ext_ram_wdata[37] ,
    \data_arrays_0_0_ext_ram_wdata[36] ,
    \data_arrays_0_0_ext_ram_wdata[35] ,
    \data_arrays_0_0_ext_ram_wdata[34] ,
    \data_arrays_0_0_ext_ram_wdata[33] ,
    \data_arrays_0_0_ext_ram_wdata[32] }),
    .dout0({\data_arrays_0_0_ext_ram_rdata1[63] ,
    \data_arrays_0_0_ext_ram_rdata1[62] ,
    \data_arrays_0_0_ext_ram_rdata1[61] ,
    \data_arrays_0_0_ext_ram_rdata1[60] ,
    \data_arrays_0_0_ext_ram_rdata1[59] ,
    \data_arrays_0_0_ext_ram_rdata1[58] ,
    \data_arrays_0_0_ext_ram_rdata1[57] ,
    \data_arrays_0_0_ext_ram_rdata1[56] ,
    \data_arrays_0_0_ext_ram_rdata1[55] ,
    \data_arrays_0_0_ext_ram_rdata1[54] ,
    \data_arrays_0_0_ext_ram_rdata1[53] ,
    \data_arrays_0_0_ext_ram_rdata1[52] ,
    \data_arrays_0_0_ext_ram_rdata1[51] ,
    \data_arrays_0_0_ext_ram_rdata1[50] ,
    \data_arrays_0_0_ext_ram_rdata1[49] ,
    \data_arrays_0_0_ext_ram_rdata1[48] ,
    \data_arrays_0_0_ext_ram_rdata1[47] ,
    \data_arrays_0_0_ext_ram_rdata1[46] ,
    \data_arrays_0_0_ext_ram_rdata1[45] ,
    \data_arrays_0_0_ext_ram_rdata1[44] ,
    \data_arrays_0_0_ext_ram_rdata1[43] ,
    \data_arrays_0_0_ext_ram_rdata1[42] ,
    \data_arrays_0_0_ext_ram_rdata1[41] ,
    \data_arrays_0_0_ext_ram_rdata1[40] ,
    \data_arrays_0_0_ext_ram_rdata1[39] ,
    \data_arrays_0_0_ext_ram_rdata1[38] ,
    \data_arrays_0_0_ext_ram_rdata1[37] ,
    \data_arrays_0_0_ext_ram_rdata1[36] ,
    \data_arrays_0_0_ext_ram_rdata1[35] ,
    \data_arrays_0_0_ext_ram_rdata1[34] ,
    \data_arrays_0_0_ext_ram_rdata1[33] ,
    \data_arrays_0_0_ext_ram_rdata1[32] }),
    .dout1({_NC65,
    _NC66,
    _NC67,
    _NC68,
    _NC69,
    _NC70,
    _NC71,
    _NC72,
    _NC73,
    _NC74,
    _NC75,
    _NC76,
    _NC77,
    _NC78,
    _NC79,
    _NC80,
    _NC81,
    _NC82,
    _NC83,
    _NC84,
    _NC85,
    _NC86,
    _NC87,
    _NC88,
    _NC89,
    _NC90,
    _NC91,
    _NC92,
    _NC93,
    _NC94,
    _NC95,
    _NC96}),
    .wmask0({\data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 data_arrays_0_0_ext_ram1l (.csb0(\data_arrays_0_0_ext_ram_csb[1] ),
    .csb1(\data_arrays_0_0_ext_ram_csb1[3] ),
    .web0(data_arrays_0_0_ext_ram_web),
    .clk0(data_arrays_0_0_ext_ram_clk1),
    .clk1(data_arrays_0_0_ext_ram_clk1),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\data_arrays_0_0_ext_ram_addr[8] ,
    \data_arrays_0_0_ext_ram_addr[7] ,
    \data_arrays_0_0_ext_ram_addr[6] ,
    \data_arrays_0_0_ext_ram_addr[5] ,
    \data_arrays_0_0_ext_ram_addr[4] ,
    \data_arrays_0_0_ext_ram_addr[3] ,
    \data_arrays_0_0_ext_ram_addr[2] ,
    \data_arrays_0_0_ext_ram_addr[1] ,
    \data_arrays_0_0_ext_ram_addr[0] }),
    .addr1({\data_arrays_0_0_ext_ram_addr1[8] ,
    \data_arrays_0_0_ext_ram_addr1[7] ,
    \data_arrays_0_0_ext_ram_addr1[6] ,
    \data_arrays_0_0_ext_ram_addr1[5] ,
    \data_arrays_0_0_ext_ram_addr1[4] ,
    \data_arrays_0_0_ext_ram_addr1[3] ,
    \data_arrays_0_0_ext_ram_addr1[2] ,
    \data_arrays_0_0_ext_ram_addr1[1] ,
    \data_arrays_0_0_ext_ram_addr1[0] }),
    .din0({\data_arrays_0_0_ext_ram_wdata[31] ,
    \data_arrays_0_0_ext_ram_wdata[30] ,
    \data_arrays_0_0_ext_ram_wdata[29] ,
    \data_arrays_0_0_ext_ram_wdata[28] ,
    \data_arrays_0_0_ext_ram_wdata[27] ,
    \data_arrays_0_0_ext_ram_wdata[26] ,
    \data_arrays_0_0_ext_ram_wdata[25] ,
    \data_arrays_0_0_ext_ram_wdata[24] ,
    \data_arrays_0_0_ext_ram_wdata[23] ,
    \data_arrays_0_0_ext_ram_wdata[22] ,
    \data_arrays_0_0_ext_ram_wdata[21] ,
    \data_arrays_0_0_ext_ram_wdata[20] ,
    \data_arrays_0_0_ext_ram_wdata[19] ,
    \data_arrays_0_0_ext_ram_wdata[18] ,
    \data_arrays_0_0_ext_ram_wdata[17] ,
    \data_arrays_0_0_ext_ram_wdata[16] ,
    \data_arrays_0_0_ext_ram_wdata[15] ,
    \data_arrays_0_0_ext_ram_wdata[14] ,
    \data_arrays_0_0_ext_ram_wdata[13] ,
    \data_arrays_0_0_ext_ram_wdata[12] ,
    \data_arrays_0_0_ext_ram_wdata[11] ,
    \data_arrays_0_0_ext_ram_wdata[10] ,
    \data_arrays_0_0_ext_ram_wdata[9] ,
    \data_arrays_0_0_ext_ram_wdata[8] ,
    \data_arrays_0_0_ext_ram_wdata[7] ,
    \data_arrays_0_0_ext_ram_wdata[6] ,
    \data_arrays_0_0_ext_ram_wdata[5] ,
    \data_arrays_0_0_ext_ram_wdata[4] ,
    \data_arrays_0_0_ext_ram_wdata[3] ,
    \data_arrays_0_0_ext_ram_wdata[2] ,
    \data_arrays_0_0_ext_ram_wdata[1] ,
    \data_arrays_0_0_ext_ram_wdata[0] }),
    .dout0({\data_arrays_0_0_ext_ram_rdata1[31] ,
    \data_arrays_0_0_ext_ram_rdata1[30] ,
    \data_arrays_0_0_ext_ram_rdata1[29] ,
    \data_arrays_0_0_ext_ram_rdata1[28] ,
    \data_arrays_0_0_ext_ram_rdata1[27] ,
    \data_arrays_0_0_ext_ram_rdata1[26] ,
    \data_arrays_0_0_ext_ram_rdata1[25] ,
    \data_arrays_0_0_ext_ram_rdata1[24] ,
    \data_arrays_0_0_ext_ram_rdata1[23] ,
    \data_arrays_0_0_ext_ram_rdata1[22] ,
    \data_arrays_0_0_ext_ram_rdata1[21] ,
    \data_arrays_0_0_ext_ram_rdata1[20] ,
    \data_arrays_0_0_ext_ram_rdata1[19] ,
    \data_arrays_0_0_ext_ram_rdata1[18] ,
    \data_arrays_0_0_ext_ram_rdata1[17] ,
    \data_arrays_0_0_ext_ram_rdata1[16] ,
    \data_arrays_0_0_ext_ram_rdata1[15] ,
    \data_arrays_0_0_ext_ram_rdata1[14] ,
    \data_arrays_0_0_ext_ram_rdata1[13] ,
    \data_arrays_0_0_ext_ram_rdata1[12] ,
    \data_arrays_0_0_ext_ram_rdata1[11] ,
    \data_arrays_0_0_ext_ram_rdata1[10] ,
    \data_arrays_0_0_ext_ram_rdata1[9] ,
    \data_arrays_0_0_ext_ram_rdata1[8] ,
    \data_arrays_0_0_ext_ram_rdata1[7] ,
    \data_arrays_0_0_ext_ram_rdata1[6] ,
    \data_arrays_0_0_ext_ram_rdata1[5] ,
    \data_arrays_0_0_ext_ram_rdata1[4] ,
    \data_arrays_0_0_ext_ram_rdata1[3] ,
    \data_arrays_0_0_ext_ram_rdata1[2] ,
    \data_arrays_0_0_ext_ram_rdata1[1] ,
    \data_arrays_0_0_ext_ram_rdata1[0] }),
    .dout1({_NC97,
    _NC98,
    _NC99,
    _NC100,
    _NC101,
    _NC102,
    _NC103,
    _NC104,
    _NC105,
    _NC106,
    _NC107,
    _NC108,
    _NC109,
    _NC110,
    _NC111,
    _NC112,
    _NC113,
    _NC114,
    _NC115,
    _NC116,
    _NC117,
    _NC118,
    _NC119,
    _NC120,
    _NC121,
    _NC122,
    _NC123,
    _NC124,
    _NC125,
    _NC126,
    _NC127,
    _NC128}),
    .wmask0({\data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 data_arrays_0_0_ext_ram2h (.csb0(\data_arrays_0_0_ext_ram_csb[2] ),
    .csb1(\data_arrays_0_0_ext_ram_csb1[4] ),
    .web0(data_arrays_0_0_ext_ram_web),
    .clk0(data_arrays_0_0_ext_ram_clk2),
    .clk1(data_arrays_0_0_ext_ram_clk2),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\data_arrays_0_0_ext_ram_addr[8] ,
    \data_arrays_0_0_ext_ram_addr[7] ,
    \data_arrays_0_0_ext_ram_addr[6] ,
    \data_arrays_0_0_ext_ram_addr[5] ,
    \data_arrays_0_0_ext_ram_addr[4] ,
    \data_arrays_0_0_ext_ram_addr[3] ,
    \data_arrays_0_0_ext_ram_addr[2] ,
    \data_arrays_0_0_ext_ram_addr[1] ,
    \data_arrays_0_0_ext_ram_addr[0] }),
    .addr1({\data_arrays_0_0_ext_ram_addr1[8] ,
    \data_arrays_0_0_ext_ram_addr1[7] ,
    \data_arrays_0_0_ext_ram_addr1[6] ,
    \data_arrays_0_0_ext_ram_addr1[5] ,
    \data_arrays_0_0_ext_ram_addr1[4] ,
    \data_arrays_0_0_ext_ram_addr1[3] ,
    \data_arrays_0_0_ext_ram_addr1[2] ,
    \data_arrays_0_0_ext_ram_addr1[1] ,
    \data_arrays_0_0_ext_ram_addr1[0] }),
    .din0({\data_arrays_0_0_ext_ram_wdata[63] ,
    \data_arrays_0_0_ext_ram_wdata[62] ,
    \data_arrays_0_0_ext_ram_wdata[61] ,
    \data_arrays_0_0_ext_ram_wdata[60] ,
    \data_arrays_0_0_ext_ram_wdata[59] ,
    \data_arrays_0_0_ext_ram_wdata[58] ,
    \data_arrays_0_0_ext_ram_wdata[57] ,
    \data_arrays_0_0_ext_ram_wdata[56] ,
    \data_arrays_0_0_ext_ram_wdata[55] ,
    \data_arrays_0_0_ext_ram_wdata[54] ,
    \data_arrays_0_0_ext_ram_wdata[53] ,
    \data_arrays_0_0_ext_ram_wdata[52] ,
    \data_arrays_0_0_ext_ram_wdata[51] ,
    \data_arrays_0_0_ext_ram_wdata[50] ,
    \data_arrays_0_0_ext_ram_wdata[49] ,
    \data_arrays_0_0_ext_ram_wdata[48] ,
    \data_arrays_0_0_ext_ram_wdata[47] ,
    \data_arrays_0_0_ext_ram_wdata[46] ,
    \data_arrays_0_0_ext_ram_wdata[45] ,
    \data_arrays_0_0_ext_ram_wdata[44] ,
    \data_arrays_0_0_ext_ram_wdata[43] ,
    \data_arrays_0_0_ext_ram_wdata[42] ,
    \data_arrays_0_0_ext_ram_wdata[41] ,
    \data_arrays_0_0_ext_ram_wdata[40] ,
    \data_arrays_0_0_ext_ram_wdata[39] ,
    \data_arrays_0_0_ext_ram_wdata[38] ,
    \data_arrays_0_0_ext_ram_wdata[37] ,
    \data_arrays_0_0_ext_ram_wdata[36] ,
    \data_arrays_0_0_ext_ram_wdata[35] ,
    \data_arrays_0_0_ext_ram_wdata[34] ,
    \data_arrays_0_0_ext_ram_wdata[33] ,
    \data_arrays_0_0_ext_ram_wdata[32] }),
    .dout0({\data_arrays_0_0_ext_ram_rdata2[63] ,
    \data_arrays_0_0_ext_ram_rdata2[62] ,
    \data_arrays_0_0_ext_ram_rdata2[61] ,
    \data_arrays_0_0_ext_ram_rdata2[60] ,
    \data_arrays_0_0_ext_ram_rdata2[59] ,
    \data_arrays_0_0_ext_ram_rdata2[58] ,
    \data_arrays_0_0_ext_ram_rdata2[57] ,
    \data_arrays_0_0_ext_ram_rdata2[56] ,
    \data_arrays_0_0_ext_ram_rdata2[55] ,
    \data_arrays_0_0_ext_ram_rdata2[54] ,
    \data_arrays_0_0_ext_ram_rdata2[53] ,
    \data_arrays_0_0_ext_ram_rdata2[52] ,
    \data_arrays_0_0_ext_ram_rdata2[51] ,
    \data_arrays_0_0_ext_ram_rdata2[50] ,
    \data_arrays_0_0_ext_ram_rdata2[49] ,
    \data_arrays_0_0_ext_ram_rdata2[48] ,
    \data_arrays_0_0_ext_ram_rdata2[47] ,
    \data_arrays_0_0_ext_ram_rdata2[46] ,
    \data_arrays_0_0_ext_ram_rdata2[45] ,
    \data_arrays_0_0_ext_ram_rdata2[44] ,
    \data_arrays_0_0_ext_ram_rdata2[43] ,
    \data_arrays_0_0_ext_ram_rdata2[42] ,
    \data_arrays_0_0_ext_ram_rdata2[41] ,
    \data_arrays_0_0_ext_ram_rdata2[40] ,
    \data_arrays_0_0_ext_ram_rdata2[39] ,
    \data_arrays_0_0_ext_ram_rdata2[38] ,
    \data_arrays_0_0_ext_ram_rdata2[37] ,
    \data_arrays_0_0_ext_ram_rdata2[36] ,
    \data_arrays_0_0_ext_ram_rdata2[35] ,
    \data_arrays_0_0_ext_ram_rdata2[34] ,
    \data_arrays_0_0_ext_ram_rdata2[33] ,
    \data_arrays_0_0_ext_ram_rdata2[32] }),
    .dout1({_NC129,
    _NC130,
    _NC131,
    _NC132,
    _NC133,
    _NC134,
    _NC135,
    _NC136,
    _NC137,
    _NC138,
    _NC139,
    _NC140,
    _NC141,
    _NC142,
    _NC143,
    _NC144,
    _NC145,
    _NC146,
    _NC147,
    _NC148,
    _NC149,
    _NC150,
    _NC151,
    _NC152,
    _NC153,
    _NC154,
    _NC155,
    _NC156,
    _NC157,
    _NC158,
    _NC159,
    _NC160}),
    .wmask0({\data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 data_arrays_0_0_ext_ram2l (.csb0(\data_arrays_0_0_ext_ram_csb[2] ),
    .csb1(\data_arrays_0_0_ext_ram_csb1[5] ),
    .web0(data_arrays_0_0_ext_ram_web),
    .clk0(data_arrays_0_0_ext_ram_clk2),
    .clk1(data_arrays_0_0_ext_ram_clk2),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\data_arrays_0_0_ext_ram_addr[8] ,
    \data_arrays_0_0_ext_ram_addr[7] ,
    \data_arrays_0_0_ext_ram_addr[6] ,
    \data_arrays_0_0_ext_ram_addr[5] ,
    \data_arrays_0_0_ext_ram_addr[4] ,
    \data_arrays_0_0_ext_ram_addr[3] ,
    \data_arrays_0_0_ext_ram_addr[2] ,
    \data_arrays_0_0_ext_ram_addr[1] ,
    \data_arrays_0_0_ext_ram_addr[0] }),
    .addr1({\data_arrays_0_0_ext_ram_addr1[8] ,
    \data_arrays_0_0_ext_ram_addr1[7] ,
    \data_arrays_0_0_ext_ram_addr1[6] ,
    \data_arrays_0_0_ext_ram_addr1[5] ,
    \data_arrays_0_0_ext_ram_addr1[4] ,
    \data_arrays_0_0_ext_ram_addr1[3] ,
    \data_arrays_0_0_ext_ram_addr1[2] ,
    \data_arrays_0_0_ext_ram_addr1[1] ,
    \data_arrays_0_0_ext_ram_addr1[0] }),
    .din0({\data_arrays_0_0_ext_ram_wdata[31] ,
    \data_arrays_0_0_ext_ram_wdata[30] ,
    \data_arrays_0_0_ext_ram_wdata[29] ,
    \data_arrays_0_0_ext_ram_wdata[28] ,
    \data_arrays_0_0_ext_ram_wdata[27] ,
    \data_arrays_0_0_ext_ram_wdata[26] ,
    \data_arrays_0_0_ext_ram_wdata[25] ,
    \data_arrays_0_0_ext_ram_wdata[24] ,
    \data_arrays_0_0_ext_ram_wdata[23] ,
    \data_arrays_0_0_ext_ram_wdata[22] ,
    \data_arrays_0_0_ext_ram_wdata[21] ,
    \data_arrays_0_0_ext_ram_wdata[20] ,
    \data_arrays_0_0_ext_ram_wdata[19] ,
    \data_arrays_0_0_ext_ram_wdata[18] ,
    \data_arrays_0_0_ext_ram_wdata[17] ,
    \data_arrays_0_0_ext_ram_wdata[16] ,
    \data_arrays_0_0_ext_ram_wdata[15] ,
    \data_arrays_0_0_ext_ram_wdata[14] ,
    \data_arrays_0_0_ext_ram_wdata[13] ,
    \data_arrays_0_0_ext_ram_wdata[12] ,
    \data_arrays_0_0_ext_ram_wdata[11] ,
    \data_arrays_0_0_ext_ram_wdata[10] ,
    \data_arrays_0_0_ext_ram_wdata[9] ,
    \data_arrays_0_0_ext_ram_wdata[8] ,
    \data_arrays_0_0_ext_ram_wdata[7] ,
    \data_arrays_0_0_ext_ram_wdata[6] ,
    \data_arrays_0_0_ext_ram_wdata[5] ,
    \data_arrays_0_0_ext_ram_wdata[4] ,
    \data_arrays_0_0_ext_ram_wdata[3] ,
    \data_arrays_0_0_ext_ram_wdata[2] ,
    \data_arrays_0_0_ext_ram_wdata[1] ,
    \data_arrays_0_0_ext_ram_wdata[0] }),
    .dout0({\data_arrays_0_0_ext_ram_rdata2[31] ,
    \data_arrays_0_0_ext_ram_rdata2[30] ,
    \data_arrays_0_0_ext_ram_rdata2[29] ,
    \data_arrays_0_0_ext_ram_rdata2[28] ,
    \data_arrays_0_0_ext_ram_rdata2[27] ,
    \data_arrays_0_0_ext_ram_rdata2[26] ,
    \data_arrays_0_0_ext_ram_rdata2[25] ,
    \data_arrays_0_0_ext_ram_rdata2[24] ,
    \data_arrays_0_0_ext_ram_rdata2[23] ,
    \data_arrays_0_0_ext_ram_rdata2[22] ,
    \data_arrays_0_0_ext_ram_rdata2[21] ,
    \data_arrays_0_0_ext_ram_rdata2[20] ,
    \data_arrays_0_0_ext_ram_rdata2[19] ,
    \data_arrays_0_0_ext_ram_rdata2[18] ,
    \data_arrays_0_0_ext_ram_rdata2[17] ,
    \data_arrays_0_0_ext_ram_rdata2[16] ,
    \data_arrays_0_0_ext_ram_rdata2[15] ,
    \data_arrays_0_0_ext_ram_rdata2[14] ,
    \data_arrays_0_0_ext_ram_rdata2[13] ,
    \data_arrays_0_0_ext_ram_rdata2[12] ,
    \data_arrays_0_0_ext_ram_rdata2[11] ,
    \data_arrays_0_0_ext_ram_rdata2[10] ,
    \data_arrays_0_0_ext_ram_rdata2[9] ,
    \data_arrays_0_0_ext_ram_rdata2[8] ,
    \data_arrays_0_0_ext_ram_rdata2[7] ,
    \data_arrays_0_0_ext_ram_rdata2[6] ,
    \data_arrays_0_0_ext_ram_rdata2[5] ,
    \data_arrays_0_0_ext_ram_rdata2[4] ,
    \data_arrays_0_0_ext_ram_rdata2[3] ,
    \data_arrays_0_0_ext_ram_rdata2[2] ,
    \data_arrays_0_0_ext_ram_rdata2[1] ,
    \data_arrays_0_0_ext_ram_rdata2[0] }),
    .dout1({_NC161,
    _NC162,
    _NC163,
    _NC164,
    _NC165,
    _NC166,
    _NC167,
    _NC168,
    _NC169,
    _NC170,
    _NC171,
    _NC172,
    _NC173,
    _NC174,
    _NC175,
    _NC176,
    _NC177,
    _NC178,
    _NC179,
    _NC180,
    _NC181,
    _NC182,
    _NC183,
    _NC184,
    _NC185,
    _NC186,
    _NC187,
    _NC188,
    _NC189,
    _NC190,
    _NC191,
    _NC192}),
    .wmask0({\data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 data_arrays_0_0_ext_ram3h (.csb0(\data_arrays_0_0_ext_ram_csb[3] ),
    .csb1(\data_arrays_0_0_ext_ram_csb1[6] ),
    .web0(data_arrays_0_0_ext_ram_web),
    .clk0(data_arrays_0_0_ext_ram_clk3),
    .clk1(data_arrays_0_0_ext_ram_clk3),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\data_arrays_0_0_ext_ram_addr[8] ,
    \data_arrays_0_0_ext_ram_addr[7] ,
    \data_arrays_0_0_ext_ram_addr[6] ,
    \data_arrays_0_0_ext_ram_addr[5] ,
    \data_arrays_0_0_ext_ram_addr[4] ,
    \data_arrays_0_0_ext_ram_addr[3] ,
    \data_arrays_0_0_ext_ram_addr[2] ,
    \data_arrays_0_0_ext_ram_addr[1] ,
    \data_arrays_0_0_ext_ram_addr[0] }),
    .addr1({\data_arrays_0_0_ext_ram_addr1[8] ,
    \data_arrays_0_0_ext_ram_addr1[7] ,
    \data_arrays_0_0_ext_ram_addr1[6] ,
    \data_arrays_0_0_ext_ram_addr1[5] ,
    \data_arrays_0_0_ext_ram_addr1[4] ,
    \data_arrays_0_0_ext_ram_addr1[3] ,
    \data_arrays_0_0_ext_ram_addr1[2] ,
    \data_arrays_0_0_ext_ram_addr1[1] ,
    \data_arrays_0_0_ext_ram_addr1[0] }),
    .din0({\data_arrays_0_0_ext_ram_wdata[63] ,
    \data_arrays_0_0_ext_ram_wdata[62] ,
    \data_arrays_0_0_ext_ram_wdata[61] ,
    \data_arrays_0_0_ext_ram_wdata[60] ,
    \data_arrays_0_0_ext_ram_wdata[59] ,
    \data_arrays_0_0_ext_ram_wdata[58] ,
    \data_arrays_0_0_ext_ram_wdata[57] ,
    \data_arrays_0_0_ext_ram_wdata[56] ,
    \data_arrays_0_0_ext_ram_wdata[55] ,
    \data_arrays_0_0_ext_ram_wdata[54] ,
    \data_arrays_0_0_ext_ram_wdata[53] ,
    \data_arrays_0_0_ext_ram_wdata[52] ,
    \data_arrays_0_0_ext_ram_wdata[51] ,
    \data_arrays_0_0_ext_ram_wdata[50] ,
    \data_arrays_0_0_ext_ram_wdata[49] ,
    \data_arrays_0_0_ext_ram_wdata[48] ,
    \data_arrays_0_0_ext_ram_wdata[47] ,
    \data_arrays_0_0_ext_ram_wdata[46] ,
    \data_arrays_0_0_ext_ram_wdata[45] ,
    \data_arrays_0_0_ext_ram_wdata[44] ,
    \data_arrays_0_0_ext_ram_wdata[43] ,
    \data_arrays_0_0_ext_ram_wdata[42] ,
    \data_arrays_0_0_ext_ram_wdata[41] ,
    \data_arrays_0_0_ext_ram_wdata[40] ,
    \data_arrays_0_0_ext_ram_wdata[39] ,
    \data_arrays_0_0_ext_ram_wdata[38] ,
    \data_arrays_0_0_ext_ram_wdata[37] ,
    \data_arrays_0_0_ext_ram_wdata[36] ,
    \data_arrays_0_0_ext_ram_wdata[35] ,
    \data_arrays_0_0_ext_ram_wdata[34] ,
    \data_arrays_0_0_ext_ram_wdata[33] ,
    \data_arrays_0_0_ext_ram_wdata[32] }),
    .dout0({\data_arrays_0_0_ext_ram_rdata3[63] ,
    \data_arrays_0_0_ext_ram_rdata3[62] ,
    \data_arrays_0_0_ext_ram_rdata3[61] ,
    \data_arrays_0_0_ext_ram_rdata3[60] ,
    \data_arrays_0_0_ext_ram_rdata3[59] ,
    \data_arrays_0_0_ext_ram_rdata3[58] ,
    \data_arrays_0_0_ext_ram_rdata3[57] ,
    \data_arrays_0_0_ext_ram_rdata3[56] ,
    \data_arrays_0_0_ext_ram_rdata3[55] ,
    \data_arrays_0_0_ext_ram_rdata3[54] ,
    \data_arrays_0_0_ext_ram_rdata3[53] ,
    \data_arrays_0_0_ext_ram_rdata3[52] ,
    \data_arrays_0_0_ext_ram_rdata3[51] ,
    \data_arrays_0_0_ext_ram_rdata3[50] ,
    \data_arrays_0_0_ext_ram_rdata3[49] ,
    \data_arrays_0_0_ext_ram_rdata3[48] ,
    \data_arrays_0_0_ext_ram_rdata3[47] ,
    \data_arrays_0_0_ext_ram_rdata3[46] ,
    \data_arrays_0_0_ext_ram_rdata3[45] ,
    \data_arrays_0_0_ext_ram_rdata3[44] ,
    \data_arrays_0_0_ext_ram_rdata3[43] ,
    \data_arrays_0_0_ext_ram_rdata3[42] ,
    \data_arrays_0_0_ext_ram_rdata3[41] ,
    \data_arrays_0_0_ext_ram_rdata3[40] ,
    \data_arrays_0_0_ext_ram_rdata3[39] ,
    \data_arrays_0_0_ext_ram_rdata3[38] ,
    \data_arrays_0_0_ext_ram_rdata3[37] ,
    \data_arrays_0_0_ext_ram_rdata3[36] ,
    \data_arrays_0_0_ext_ram_rdata3[35] ,
    \data_arrays_0_0_ext_ram_rdata3[34] ,
    \data_arrays_0_0_ext_ram_rdata3[33] ,
    \data_arrays_0_0_ext_ram_rdata3[32] }),
    .dout1({_NC193,
    _NC194,
    _NC195,
    _NC196,
    _NC197,
    _NC198,
    _NC199,
    _NC200,
    _NC201,
    _NC202,
    _NC203,
    _NC204,
    _NC205,
    _NC206,
    _NC207,
    _NC208,
    _NC209,
    _NC210,
    _NC211,
    _NC212,
    _NC213,
    _NC214,
    _NC215,
    _NC216,
    _NC217,
    _NC218,
    _NC219,
    _NC220,
    _NC221,
    _NC222,
    _NC223,
    _NC224}),
    .wmask0({\data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] ,
    \data_arrays_0_0_ext_ram_wmask[1] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 data_arrays_0_0_ext_ram3l (.csb0(\data_arrays_0_0_ext_ram_csb[3] ),
    .csb1(\data_arrays_0_0_ext_ram_csb1[7] ),
    .web0(data_arrays_0_0_ext_ram_web),
    .clk0(data_arrays_0_0_ext_ram_clk3),
    .clk1(data_arrays_0_0_ext_ram_clk3),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\data_arrays_0_0_ext_ram_addr[8] ,
    \data_arrays_0_0_ext_ram_addr[7] ,
    \data_arrays_0_0_ext_ram_addr[6] ,
    \data_arrays_0_0_ext_ram_addr[5] ,
    \data_arrays_0_0_ext_ram_addr[4] ,
    \data_arrays_0_0_ext_ram_addr[3] ,
    \data_arrays_0_0_ext_ram_addr[2] ,
    \data_arrays_0_0_ext_ram_addr[1] ,
    \data_arrays_0_0_ext_ram_addr[0] }),
    .addr1({\data_arrays_0_0_ext_ram_addr1[8] ,
    \data_arrays_0_0_ext_ram_addr1[7] ,
    \data_arrays_0_0_ext_ram_addr1[6] ,
    \data_arrays_0_0_ext_ram_addr1[5] ,
    \data_arrays_0_0_ext_ram_addr1[4] ,
    \data_arrays_0_0_ext_ram_addr1[3] ,
    \data_arrays_0_0_ext_ram_addr1[2] ,
    \data_arrays_0_0_ext_ram_addr1[1] ,
    \data_arrays_0_0_ext_ram_addr1[0] }),
    .din0({\data_arrays_0_0_ext_ram_wdata[31] ,
    \data_arrays_0_0_ext_ram_wdata[30] ,
    \data_arrays_0_0_ext_ram_wdata[29] ,
    \data_arrays_0_0_ext_ram_wdata[28] ,
    \data_arrays_0_0_ext_ram_wdata[27] ,
    \data_arrays_0_0_ext_ram_wdata[26] ,
    \data_arrays_0_0_ext_ram_wdata[25] ,
    \data_arrays_0_0_ext_ram_wdata[24] ,
    \data_arrays_0_0_ext_ram_wdata[23] ,
    \data_arrays_0_0_ext_ram_wdata[22] ,
    \data_arrays_0_0_ext_ram_wdata[21] ,
    \data_arrays_0_0_ext_ram_wdata[20] ,
    \data_arrays_0_0_ext_ram_wdata[19] ,
    \data_arrays_0_0_ext_ram_wdata[18] ,
    \data_arrays_0_0_ext_ram_wdata[17] ,
    \data_arrays_0_0_ext_ram_wdata[16] ,
    \data_arrays_0_0_ext_ram_wdata[15] ,
    \data_arrays_0_0_ext_ram_wdata[14] ,
    \data_arrays_0_0_ext_ram_wdata[13] ,
    \data_arrays_0_0_ext_ram_wdata[12] ,
    \data_arrays_0_0_ext_ram_wdata[11] ,
    \data_arrays_0_0_ext_ram_wdata[10] ,
    \data_arrays_0_0_ext_ram_wdata[9] ,
    \data_arrays_0_0_ext_ram_wdata[8] ,
    \data_arrays_0_0_ext_ram_wdata[7] ,
    \data_arrays_0_0_ext_ram_wdata[6] ,
    \data_arrays_0_0_ext_ram_wdata[5] ,
    \data_arrays_0_0_ext_ram_wdata[4] ,
    \data_arrays_0_0_ext_ram_wdata[3] ,
    \data_arrays_0_0_ext_ram_wdata[2] ,
    \data_arrays_0_0_ext_ram_wdata[1] ,
    \data_arrays_0_0_ext_ram_wdata[0] }),
    .dout0({\data_arrays_0_0_ext_ram_rdata3[31] ,
    \data_arrays_0_0_ext_ram_rdata3[30] ,
    \data_arrays_0_0_ext_ram_rdata3[29] ,
    \data_arrays_0_0_ext_ram_rdata3[28] ,
    \data_arrays_0_0_ext_ram_rdata3[27] ,
    \data_arrays_0_0_ext_ram_rdata3[26] ,
    \data_arrays_0_0_ext_ram_rdata3[25] ,
    \data_arrays_0_0_ext_ram_rdata3[24] ,
    \data_arrays_0_0_ext_ram_rdata3[23] ,
    \data_arrays_0_0_ext_ram_rdata3[22] ,
    \data_arrays_0_0_ext_ram_rdata3[21] ,
    \data_arrays_0_0_ext_ram_rdata3[20] ,
    \data_arrays_0_0_ext_ram_rdata3[19] ,
    \data_arrays_0_0_ext_ram_rdata3[18] ,
    \data_arrays_0_0_ext_ram_rdata3[17] ,
    \data_arrays_0_0_ext_ram_rdata3[16] ,
    \data_arrays_0_0_ext_ram_rdata3[15] ,
    \data_arrays_0_0_ext_ram_rdata3[14] ,
    \data_arrays_0_0_ext_ram_rdata3[13] ,
    \data_arrays_0_0_ext_ram_rdata3[12] ,
    \data_arrays_0_0_ext_ram_rdata3[11] ,
    \data_arrays_0_0_ext_ram_rdata3[10] ,
    \data_arrays_0_0_ext_ram_rdata3[9] ,
    \data_arrays_0_0_ext_ram_rdata3[8] ,
    \data_arrays_0_0_ext_ram_rdata3[7] ,
    \data_arrays_0_0_ext_ram_rdata3[6] ,
    \data_arrays_0_0_ext_ram_rdata3[5] ,
    \data_arrays_0_0_ext_ram_rdata3[4] ,
    \data_arrays_0_0_ext_ram_rdata3[3] ,
    \data_arrays_0_0_ext_ram_rdata3[2] ,
    \data_arrays_0_0_ext_ram_rdata3[1] ,
    \data_arrays_0_0_ext_ram_rdata3[0] }),
    .dout1({_NC225,
    _NC226,
    _NC227,
    _NC228,
    _NC229,
    _NC230,
    _NC231,
    _NC232,
    _NC233,
    _NC234,
    _NC235,
    _NC236,
    _NC237,
    _NC238,
    _NC239,
    _NC240,
    _NC241,
    _NC242,
    _NC243,
    _NC244,
    _NC245,
    _NC246,
    _NC247,
    _NC248,
    _NC249,
    _NC250,
    _NC251,
    _NC252,
    _NC253,
    _NC254,
    _NC255,
    _NC256}),
    .wmask0({\data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] ,
    \data_arrays_0_0_ext_ram_wmask[0] }));
 sky130_sram_1kbyte_1rw1r_32x256_8 tag_array_ext_ram0h (.csb0(tag_array_ext_ram_csb),
    .csb1(\tag_array_ext_ram_csb1[1] ),
    .web0(tag_array_ext_ram_web),
    .clk0(tag_array_ext_ram_clk),
    .clk1(tag_array_ext_ram_clk),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\tag_array_ext_ram_addr[7] ,
    \tag_array_ext_ram_addr[6] ,
    \tag_array_ext_ram_addr[5] ,
    \tag_array_ext_ram_addr[4] ,
    \tag_array_ext_ram_addr[3] ,
    \tag_array_ext_ram_addr[2] ,
    \tag_array_ext_ram_addr[1] ,
    \tag_array_ext_ram_addr[0] }),
    .addr1({\tag_array_ext_ram_addr1[7] ,
    \tag_array_ext_ram_addr1[6] ,
    \tag_array_ext_ram_addr1[5] ,
    \tag_array_ext_ram_addr1[4] ,
    \tag_array_ext_ram_addr1[3] ,
    \tag_array_ext_ram_addr1[2] ,
    \tag_array_ext_ram_addr1[1] ,
    \tag_array_ext_ram_addr1[0] }),
    .din0({\tag_array_ext_ram_wdata[63] ,
    \tag_array_ext_ram_wdata[62] ,
    \tag_array_ext_ram_wdata[61] ,
    \tag_array_ext_ram_wdata[60] ,
    \tag_array_ext_ram_wdata[59] ,
    \tag_array_ext_ram_wdata[58] ,
    \tag_array_ext_ram_wdata[57] ,
    \tag_array_ext_ram_wdata[56] ,
    \tag_array_ext_ram_wdata[55] ,
    \tag_array_ext_ram_wdata[54] ,
    \tag_array_ext_ram_wdata[53] ,
    \tag_array_ext_ram_wdata[52] ,
    \tag_array_ext_ram_wdata[51] ,
    \tag_array_ext_ram_wdata[50] ,
    \tag_array_ext_ram_wdata[49] ,
    \tag_array_ext_ram_wdata[48] ,
    \tag_array_ext_ram_wdata[47] ,
    \tag_array_ext_ram_wdata[46] ,
    \tag_array_ext_ram_wdata[45] ,
    \tag_array_ext_ram_wdata[44] ,
    \tag_array_ext_ram_wdata[43] ,
    \tag_array_ext_ram_wdata[42] ,
    \tag_array_ext_ram_wdata[41] ,
    \tag_array_ext_ram_wdata[40] ,
    \tag_array_ext_ram_wdata[39] ,
    \tag_array_ext_ram_wdata[38] ,
    \tag_array_ext_ram_wdata[37] ,
    \tag_array_ext_ram_wdata[36] ,
    \tag_array_ext_ram_wdata[35] ,
    \tag_array_ext_ram_wdata[34] ,
    \tag_array_ext_ram_wdata[33] ,
    \tag_array_ext_ram_wdata[32] }),
    .dout0({\tag_array_ext_ram_rdata1[31] ,
    \tag_array_ext_ram_rdata1[30] ,
    \tag_array_ext_ram_rdata1[29] ,
    \tag_array_ext_ram_rdata1[28] ,
    \tag_array_ext_ram_rdata1[27] ,
    \tag_array_ext_ram_rdata1[26] ,
    \tag_array_ext_ram_rdata1[25] ,
    \tag_array_ext_ram_rdata1[24] ,
    \tag_array_ext_ram_rdata1[23] ,
    \tag_array_ext_ram_rdata1[22] ,
    \tag_array_ext_ram_rdata1[21] ,
    \tag_array_ext_ram_rdata1[20] ,
    \tag_array_ext_ram_rdata1[19] ,
    \tag_array_ext_ram_rdata1[18] ,
    \tag_array_ext_ram_rdata1[17] ,
    \tag_array_ext_ram_rdata1[16] ,
    \tag_array_ext_ram_rdata1[15] ,
    \tag_array_ext_ram_rdata1[14] ,
    \tag_array_ext_ram_rdata1[13] ,
    \tag_array_ext_ram_rdata1[12] ,
    \tag_array_ext_ram_rdata1[11] ,
    \tag_array_ext_ram_rdata1[10] ,
    \tag_array_ext_ram_rdata1[9] ,
    \tag_array_ext_ram_rdata1[8] ,
    \tag_array_ext_ram_rdata1[7] ,
    \tag_array_ext_ram_rdata1[6] ,
    \tag_array_ext_ram_rdata1[5] ,
    \tag_array_ext_ram_rdata1[4] ,
    \tag_array_ext_ram_rdata1[3] ,
    \tag_array_ext_ram_rdata1[2] ,
    \tag_array_ext_ram_rdata1[1] ,
    \tag_array_ext_ram_rdata1[0] }),
    .dout1({_NC257,
    _NC258,
    _NC259,
    _NC260,
    _NC261,
    _NC262,
    _NC263,
    _NC264,
    _NC265,
    _NC266,
    _NC267,
    _NC268,
    _NC269,
    _NC270,
    _NC271,
    _NC272,
    _NC273,
    _NC274,
    _NC275,
    _NC276,
    _NC277,
    _NC278,
    _NC279,
    _NC280,
    _NC281,
    _NC282,
    _NC283,
    _NC284,
    _NC285,
    _NC286,
    _NC287,
    _NC288}),
    .wmask0({\tag_array_ext_ram_wmask[1] ,
    \tag_array_ext_ram_wmask[1] ,
    \tag_array_ext_ram_wmask[1] ,
    \tag_array_ext_ram_wmask[1] }));
 sky130_sram_1kbyte_1rw1r_32x256_8 tag_array_ext_ram0l (.csb0(tag_array_ext_ram_csb),
    .csb1(\tag_array_ext_ram_csb1[0] ),
    .web0(tag_array_ext_ram_web),
    .clk0(tag_array_ext_ram_clk),
    .clk1(tag_array_ext_ram_clk),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\tag_array_ext_ram_addr[7] ,
    \tag_array_ext_ram_addr[6] ,
    \tag_array_ext_ram_addr[5] ,
    \tag_array_ext_ram_addr[4] ,
    \tag_array_ext_ram_addr[3] ,
    \tag_array_ext_ram_addr[2] ,
    \tag_array_ext_ram_addr[1] ,
    \tag_array_ext_ram_addr[0] }),
    .addr1({\tag_array_ext_ram_addr1[7] ,
    \tag_array_ext_ram_addr1[6] ,
    \tag_array_ext_ram_addr1[5] ,
    \tag_array_ext_ram_addr1[4] ,
    \tag_array_ext_ram_addr1[3] ,
    \tag_array_ext_ram_addr1[2] ,
    \tag_array_ext_ram_addr1[1] ,
    \tag_array_ext_ram_addr1[0] }),
    .din0({\tag_array_ext_ram_wdata[31] ,
    \tag_array_ext_ram_wdata[30] ,
    \tag_array_ext_ram_wdata[29] ,
    \tag_array_ext_ram_wdata[28] ,
    \tag_array_ext_ram_wdata[27] ,
    \tag_array_ext_ram_wdata[26] ,
    \tag_array_ext_ram_wdata[25] ,
    \tag_array_ext_ram_wdata[24] ,
    \tag_array_ext_ram_wdata[23] ,
    \tag_array_ext_ram_wdata[22] ,
    \tag_array_ext_ram_wdata[21] ,
    \tag_array_ext_ram_wdata[20] ,
    \tag_array_ext_ram_wdata[19] ,
    \tag_array_ext_ram_wdata[18] ,
    \tag_array_ext_ram_wdata[17] ,
    \tag_array_ext_ram_wdata[16] ,
    \tag_array_ext_ram_wdata[15] ,
    \tag_array_ext_ram_wdata[14] ,
    \tag_array_ext_ram_wdata[13] ,
    \tag_array_ext_ram_wdata[12] ,
    \tag_array_ext_ram_wdata[11] ,
    \tag_array_ext_ram_wdata[10] ,
    \tag_array_ext_ram_wdata[9] ,
    \tag_array_ext_ram_wdata[8] ,
    \tag_array_ext_ram_wdata[7] ,
    \tag_array_ext_ram_wdata[6] ,
    \tag_array_ext_ram_wdata[5] ,
    \tag_array_ext_ram_wdata[4] ,
    \tag_array_ext_ram_wdata[3] ,
    \tag_array_ext_ram_wdata[2] ,
    \tag_array_ext_ram_wdata[1] ,
    \tag_array_ext_ram_wdata[0] }),
    .dout0({\tag_array_ext_ram_rdata0[31] ,
    \tag_array_ext_ram_rdata0[30] ,
    \tag_array_ext_ram_rdata0[29] ,
    \tag_array_ext_ram_rdata0[28] ,
    \tag_array_ext_ram_rdata0[27] ,
    \tag_array_ext_ram_rdata0[26] ,
    \tag_array_ext_ram_rdata0[25] ,
    \tag_array_ext_ram_rdata0[24] ,
    \tag_array_ext_ram_rdata0[23] ,
    \tag_array_ext_ram_rdata0[22] ,
    \tag_array_ext_ram_rdata0[21] ,
    \tag_array_ext_ram_rdata0[20] ,
    \tag_array_ext_ram_rdata0[19] ,
    \tag_array_ext_ram_rdata0[18] ,
    \tag_array_ext_ram_rdata0[17] ,
    \tag_array_ext_ram_rdata0[16] ,
    \tag_array_ext_ram_rdata0[15] ,
    \tag_array_ext_ram_rdata0[14] ,
    \tag_array_ext_ram_rdata0[13] ,
    \tag_array_ext_ram_rdata0[12] ,
    \tag_array_ext_ram_rdata0[11] ,
    \tag_array_ext_ram_rdata0[10] ,
    \tag_array_ext_ram_rdata0[9] ,
    \tag_array_ext_ram_rdata0[8] ,
    \tag_array_ext_ram_rdata0[7] ,
    \tag_array_ext_ram_rdata0[6] ,
    \tag_array_ext_ram_rdata0[5] ,
    \tag_array_ext_ram_rdata0[4] ,
    \tag_array_ext_ram_rdata0[3] ,
    \tag_array_ext_ram_rdata0[2] ,
    \tag_array_ext_ram_rdata0[1] ,
    \tag_array_ext_ram_rdata0[0] }),
    .dout1({_NC289,
    _NC290,
    _NC291,
    _NC292,
    _NC293,
    _NC294,
    _NC295,
    _NC296,
    _NC297,
    _NC298,
    _NC299,
    _NC300,
    _NC301,
    _NC302,
    _NC303,
    _NC304,
    _NC305,
    _NC306,
    _NC307,
    _NC308,
    _NC309,
    _NC310,
    _NC311,
    _NC312,
    _NC313,
    _NC314,
    _NC315,
    _NC316,
    _NC317,
    _NC318,
    _NC319,
    _NC320}),
    .wmask0({\tag_array_ext_ram_wmask[0] ,
    \tag_array_ext_ram_wmask[0] ,
    \tag_array_ext_ram_wmask[0] ,
    \tag_array_ext_ram_wmask[0] }));
 clk_skew_adjust u_clk_skew_adjust_0 (.clk_in(wb_clk_i),
    .clk_out(tag_array_ext_ram_clk),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\ram_clk_delay_sel[4] ,
    \ram_clk_delay_sel[3] ,
    \ram_clk_delay_sel[2] ,
    \ram_clk_delay_sel[1] ,
    \ram_clk_delay_sel[0] }));
 clk_skew_adjust u_clk_skew_adjust_1 (.clk_in(wb_clk_i),
    .clk_out(data_arrays_0_0_ext_ram_clk0),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\ram_clk_delay_sel[9] ,
    \ram_clk_delay_sel[8] ,
    \ram_clk_delay_sel[7] ,
    \ram_clk_delay_sel[6] ,
    \ram_clk_delay_sel[5] }));
 clk_skew_adjust u_clk_skew_adjust_2 (.clk_in(wb_clk_i),
    .clk_out(data_arrays_0_0_ext_ram_clk1),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\ram_clk_delay_sel[14] ,
    \ram_clk_delay_sel[13] ,
    \ram_clk_delay_sel[12] ,
    \ram_clk_delay_sel[11] ,
    \ram_clk_delay_sel[10] }));
 clk_skew_adjust u_clk_skew_adjust_3 (.clk_in(wb_clk_i),
    .clk_out(data_arrays_0_0_ext_ram_clk2),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\ram_clk_delay_sel[19] ,
    \ram_clk_delay_sel[18] ,
    \ram_clk_delay_sel[17] ,
    \ram_clk_delay_sel[16] ,
    \ram_clk_delay_sel[15] }));
 clk_skew_adjust u_clk_skew_adjust_4 (.clk_in(wb_clk_i),
    .clk_out(data_arrays_0_0_ext_ram_clk3),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\ram_clk_delay_sel[24] ,
    \ram_clk_delay_sel[23] ,
    \ram_clk_delay_sel[22] ,
    \ram_clk_delay_sel[21] ,
    \ram_clk_delay_sel[20] }));
endmodule
