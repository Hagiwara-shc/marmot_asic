VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Marmot
  CLASS BLOCK ;
  FOREIGN Marmot ;
  ORIGIN 0.000 0.000 ;
  SIZE 1767.395 BY 1778.115 ;
  PIN data_arrays_0_0_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END data_arrays_0_0_ext_ram_addr1[0]
  PIN data_arrays_0_0_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END data_arrays_0_0_ext_ram_addr1[1]
  PIN data_arrays_0_0_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 772.520 4.000 773.120 ;
    END
  END data_arrays_0_0_ext_ram_addr1[2]
  PIN data_arrays_0_0_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.920 4.000 776.520 ;
    END
  END data_arrays_0_0_ext_ram_addr1[3]
  PIN data_arrays_0_0_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END data_arrays_0_0_ext_ram_addr1[4]
  PIN data_arrays_0_0_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END data_arrays_0_0_ext_ram_addr1[5]
  PIN data_arrays_0_0_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END data_arrays_0_0_ext_ram_addr1[6]
  PIN data_arrays_0_0_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 789.520 4.000 790.120 ;
    END
  END data_arrays_0_0_ext_ram_addr1[7]
  PIN data_arrays_0_0_ext_ram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 793.600 4.000 794.200 ;
    END
  END data_arrays_0_0_ext_ram_addr1[8]
  PIN data_arrays_0_0_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END data_arrays_0_0_ext_ram_addr[0]
  PIN data_arrays_0_0_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END data_arrays_0_0_ext_ram_addr[1]
  PIN data_arrays_0_0_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END data_arrays_0_0_ext_ram_addr[2]
  PIN data_arrays_0_0_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END data_arrays_0_0_ext_ram_addr[3]
  PIN data_arrays_0_0_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END data_arrays_0_0_ext_ram_addr[4]
  PIN data_arrays_0_0_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END data_arrays_0_0_ext_ram_addr[5]
  PIN data_arrays_0_0_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END data_arrays_0_0_ext_ram_addr[6]
  PIN data_arrays_0_0_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END data_arrays_0_0_ext_ram_addr[7]
  PIN data_arrays_0_0_ext_ram_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END data_arrays_0_0_ext_ram_addr[8]
  PIN data_arrays_0_0_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 483.520 4.000 484.120 ;
    END
  END data_arrays_0_0_ext_ram_clk
  PIN data_arrays_0_0_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END data_arrays_0_0_ext_ram_csb1[0]
  PIN data_arrays_0_0_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 740.560 4.000 741.160 ;
    END
  END data_arrays_0_0_ext_ram_csb1[1]
  PIN data_arrays_0_0_ext_ram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END data_arrays_0_0_ext_ram_csb1[2]
  PIN data_arrays_0_0_ext_ram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 747.360 4.000 747.960 ;
    END
  END data_arrays_0_0_ext_ram_csb1[3]
  PIN data_arrays_0_0_ext_ram_csb1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.760 4.000 751.360 ;
    END
  END data_arrays_0_0_ext_ram_csb1[4]
  PIN data_arrays_0_0_ext_ram_csb1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END data_arrays_0_0_ext_ram_csb1[5]
  PIN data_arrays_0_0_ext_ram_csb1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END data_arrays_0_0_ext_ram_csb1[6]
  PIN data_arrays_0_0_ext_ram_csb1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END data_arrays_0_0_ext_ram_csb1[7]
  PIN data_arrays_0_0_ext_ram_csb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END data_arrays_0_0_ext_ram_csb[0]
  PIN data_arrays_0_0_ext_ram_csb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END data_arrays_0_0_ext_ram_csb[1]
  PIN data_arrays_0_0_ext_ram_csb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END data_arrays_0_0_ext_ram_csb[2]
  PIN data_arrays_0_0_ext_ram_csb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END data_arrays_0_0_ext_ram_csb[3]
  PIN data_arrays_0_0_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[0]
  PIN data_arrays_0_0_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[10]
  PIN data_arrays_0_0_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[11]
  PIN data_arrays_0_0_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[12]
  PIN data_arrays_0_0_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[13]
  PIN data_arrays_0_0_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[14]
  PIN data_arrays_0_0_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[15]
  PIN data_arrays_0_0_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[16]
  PIN data_arrays_0_0_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[17]
  PIN data_arrays_0_0_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[18]
  PIN data_arrays_0_0_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[19]
  PIN data_arrays_0_0_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[1]
  PIN data_arrays_0_0_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[20]
  PIN data_arrays_0_0_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[21]
  PIN data_arrays_0_0_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[22]
  PIN data_arrays_0_0_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[23]
  PIN data_arrays_0_0_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[24]
  PIN data_arrays_0_0_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[25]
  PIN data_arrays_0_0_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[26]
  PIN data_arrays_0_0_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[27]
  PIN data_arrays_0_0_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[28]
  PIN data_arrays_0_0_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[29]
  PIN data_arrays_0_0_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[2]
  PIN data_arrays_0_0_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[30]
  PIN data_arrays_0_0_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[31]
  PIN data_arrays_0_0_ext_ram_rdata0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[32]
  PIN data_arrays_0_0_ext_ram_rdata0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[33]
  PIN data_arrays_0_0_ext_ram_rdata0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[34]
  PIN data_arrays_0_0_ext_ram_rdata0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[35]
  PIN data_arrays_0_0_ext_ram_rdata0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[36]
  PIN data_arrays_0_0_ext_ram_rdata0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[37]
  PIN data_arrays_0_0_ext_ram_rdata0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[38]
  PIN data_arrays_0_0_ext_ram_rdata0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[39]
  PIN data_arrays_0_0_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[3]
  PIN data_arrays_0_0_ext_ram_rdata0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[40]
  PIN data_arrays_0_0_ext_ram_rdata0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[41]
  PIN data_arrays_0_0_ext_ram_rdata0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[42]
  PIN data_arrays_0_0_ext_ram_rdata0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[43]
  PIN data_arrays_0_0_ext_ram_rdata0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[44]
  PIN data_arrays_0_0_ext_ram_rdata0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[45]
  PIN data_arrays_0_0_ext_ram_rdata0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[46]
  PIN data_arrays_0_0_ext_ram_rdata0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[47]
  PIN data_arrays_0_0_ext_ram_rdata0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[48]
  PIN data_arrays_0_0_ext_ram_rdata0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[49]
  PIN data_arrays_0_0_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[4]
  PIN data_arrays_0_0_ext_ram_rdata0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[50]
  PIN data_arrays_0_0_ext_ram_rdata0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[51]
  PIN data_arrays_0_0_ext_ram_rdata0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[52]
  PIN data_arrays_0_0_ext_ram_rdata0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[53]
  PIN data_arrays_0_0_ext_ram_rdata0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[54]
  PIN data_arrays_0_0_ext_ram_rdata0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[55]
  PIN data_arrays_0_0_ext_ram_rdata0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[56]
  PIN data_arrays_0_0_ext_ram_rdata0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[57]
  PIN data_arrays_0_0_ext_ram_rdata0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[58]
  PIN data_arrays_0_0_ext_ram_rdata0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[59]
  PIN data_arrays_0_0_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[5]
  PIN data_arrays_0_0_ext_ram_rdata0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[60]
  PIN data_arrays_0_0_ext_ram_rdata0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[61]
  PIN data_arrays_0_0_ext_ram_rdata0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[62]
  PIN data_arrays_0_0_ext_ram_rdata0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[63]
  PIN data_arrays_0_0_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[6]
  PIN data_arrays_0_0_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[7]
  PIN data_arrays_0_0_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[8]
  PIN data_arrays_0_0_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata0[9]
  PIN data_arrays_0_0_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[0]
  PIN data_arrays_0_0_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[10]
  PIN data_arrays_0_0_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[11]
  PIN data_arrays_0_0_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[12]
  PIN data_arrays_0_0_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[13]
  PIN data_arrays_0_0_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[14]
  PIN data_arrays_0_0_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[15]
  PIN data_arrays_0_0_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[16]
  PIN data_arrays_0_0_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[17]
  PIN data_arrays_0_0_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[18]
  PIN data_arrays_0_0_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[19]
  PIN data_arrays_0_0_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[1]
  PIN data_arrays_0_0_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[20]
  PIN data_arrays_0_0_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[21]
  PIN data_arrays_0_0_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[22]
  PIN data_arrays_0_0_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[23]
  PIN data_arrays_0_0_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[24]
  PIN data_arrays_0_0_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[25]
  PIN data_arrays_0_0_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[26]
  PIN data_arrays_0_0_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[27]
  PIN data_arrays_0_0_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[28]
  PIN data_arrays_0_0_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[29]
  PIN data_arrays_0_0_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[2]
  PIN data_arrays_0_0_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[30]
  PIN data_arrays_0_0_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[31]
  PIN data_arrays_0_0_ext_ram_rdata1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[32]
  PIN data_arrays_0_0_ext_ram_rdata1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[33]
  PIN data_arrays_0_0_ext_ram_rdata1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[34]
  PIN data_arrays_0_0_ext_ram_rdata1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[35]
  PIN data_arrays_0_0_ext_ram_rdata1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[36]
  PIN data_arrays_0_0_ext_ram_rdata1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[37]
  PIN data_arrays_0_0_ext_ram_rdata1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[38]
  PIN data_arrays_0_0_ext_ram_rdata1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[39]
  PIN data_arrays_0_0_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[3]
  PIN data_arrays_0_0_ext_ram_rdata1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[40]
  PIN data_arrays_0_0_ext_ram_rdata1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[41]
  PIN data_arrays_0_0_ext_ram_rdata1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[42]
  PIN data_arrays_0_0_ext_ram_rdata1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[43]
  PIN data_arrays_0_0_ext_ram_rdata1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[44]
  PIN data_arrays_0_0_ext_ram_rdata1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[45]
  PIN data_arrays_0_0_ext_ram_rdata1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[46]
  PIN data_arrays_0_0_ext_ram_rdata1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[47]
  PIN data_arrays_0_0_ext_ram_rdata1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[48]
  PIN data_arrays_0_0_ext_ram_rdata1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[49]
  PIN data_arrays_0_0_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[4]
  PIN data_arrays_0_0_ext_ram_rdata1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[50]
  PIN data_arrays_0_0_ext_ram_rdata1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[51]
  PIN data_arrays_0_0_ext_ram_rdata1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[52]
  PIN data_arrays_0_0_ext_ram_rdata1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[53]
  PIN data_arrays_0_0_ext_ram_rdata1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 4.000 417.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[54]
  PIN data_arrays_0_0_ext_ram_rdata1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[55]
  PIN data_arrays_0_0_ext_ram_rdata1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[56]
  PIN data_arrays_0_0_ext_ram_rdata1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[57]
  PIN data_arrays_0_0_ext_ram_rdata1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[58]
  PIN data_arrays_0_0_ext_ram_rdata1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[59]
  PIN data_arrays_0_0_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[5]
  PIN data_arrays_0_0_ext_ram_rdata1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[60]
  PIN data_arrays_0_0_ext_ram_rdata1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[61]
  PIN data_arrays_0_0_ext_ram_rdata1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[62]
  PIN data_arrays_0_0_ext_ram_rdata1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.160 4.000 448.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[63]
  PIN data_arrays_0_0_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[6]
  PIN data_arrays_0_0_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[7]
  PIN data_arrays_0_0_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[8]
  PIN data_arrays_0_0_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata1[9]
  PIN data_arrays_0_0_ext_ram_rdata2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[0]
  PIN data_arrays_0_0_ext_ram_rdata2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[10]
  PIN data_arrays_0_0_ext_ram_rdata2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.760 4.000 836.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[11]
  PIN data_arrays_0_0_ext_ram_rdata2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[12]
  PIN data_arrays_0_0_ext_ram_rdata2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 842.560 4.000 843.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[13]
  PIN data_arrays_0_0_ext_ram_rdata2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.960 4.000 846.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[14]
  PIN data_arrays_0_0_ext_ram_rdata2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 849.360 4.000 849.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[15]
  PIN data_arrays_0_0_ext_ram_rdata2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[16]
  PIN data_arrays_0_0_ext_ram_rdata2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[17]
  PIN data_arrays_0_0_ext_ram_rdata2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[18]
  PIN data_arrays_0_0_ext_ram_rdata2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[19]
  PIN data_arrays_0_0_ext_ram_rdata2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 800.400 4.000 801.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[1]
  PIN data_arrays_0_0_ext_ram_rdata2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[20]
  PIN data_arrays_0_0_ext_ram_rdata2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.120 4.000 871.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[21]
  PIN data_arrays_0_0_ext_ram_rdata2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 874.520 4.000 875.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[22]
  PIN data_arrays_0_0_ext_ram_rdata2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.920 4.000 878.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[23]
  PIN data_arrays_0_0_ext_ram_rdata2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[24]
  PIN data_arrays_0_0_ext_ram_rdata2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.720 4.000 885.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[25]
  PIN data_arrays_0_0_ext_ram_rdata2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[26]
  PIN data_arrays_0_0_ext_ram_rdata2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[27]
  PIN data_arrays_0_0_ext_ram_rdata2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 895.600 4.000 896.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[28]
  PIN data_arrays_0_0_ext_ram_rdata2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[29]
  PIN data_arrays_0_0_ext_ram_rdata2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.800 4.000 804.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[2]
  PIN data_arrays_0_0_ext_ram_rdata2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 902.400 4.000 903.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[30]
  PIN data_arrays_0_0_ext_ram_rdata2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[31]
  PIN data_arrays_0_0_ext_ram_rdata2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.200 4.000 909.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[32]
  PIN data_arrays_0_0_ext_ram_rdata2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.280 4.000 913.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[33]
  PIN data_arrays_0_0_ext_ram_rdata2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[34]
  PIN data_arrays_0_0_ext_ram_rdata2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[35]
  PIN data_arrays_0_0_ext_ram_rdata2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 923.480 4.000 924.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[36]
  PIN data_arrays_0_0_ext_ram_rdata2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.880 4.000 927.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[37]
  PIN data_arrays_0_0_ext_ram_rdata2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[38]
  PIN data_arrays_0_0_ext_ram_rdata2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 4.000 934.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[39]
  PIN data_arrays_0_0_ext_ram_rdata2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.200 4.000 807.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[3]
  PIN data_arrays_0_0_ext_ram_rdata2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.760 4.000 938.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[40]
  PIN data_arrays_0_0_ext_ram_rdata2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[41]
  PIN data_arrays_0_0_ext_ram_rdata2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 944.560 4.000 945.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[42]
  PIN data_arrays_0_0_ext_ram_rdata2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[43]
  PIN data_arrays_0_0_ext_ram_rdata2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[44]
  PIN data_arrays_0_0_ext_ram_rdata2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[45]
  PIN data_arrays_0_0_ext_ram_rdata2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[46]
  PIN data_arrays_0_0_ext_ram_rdata2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[47]
  PIN data_arrays_0_0_ext_ram_rdata2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[48]
  PIN data_arrays_0_0_ext_ram_rdata2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.720 4.000 970.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[49]
  PIN data_arrays_0_0_ext_ram_rdata2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[4]
  PIN data_arrays_0_0_ext_ram_rdata2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.120 4.000 973.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[50]
  PIN data_arrays_0_0_ext_ram_rdata2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 976.520 4.000 977.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[51]
  PIN data_arrays_0_0_ext_ram_rdata2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.920 4.000 980.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[52]
  PIN data_arrays_0_0_ext_ram_rdata2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[53]
  PIN data_arrays_0_0_ext_ram_rdata2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.720 4.000 987.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[54]
  PIN data_arrays_0_0_ext_ram_rdata2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.800 4.000 991.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[55]
  PIN data_arrays_0_0_ext_ram_rdata2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[56]
  PIN data_arrays_0_0_ext_ram_rdata2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 997.600 4.000 998.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[57]
  PIN data_arrays_0_0_ext_ram_rdata2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.000 4.000 1001.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[58]
  PIN data_arrays_0_0_ext_ram_rdata2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1004.400 4.000 1005.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[59]
  PIN data_arrays_0_0_ext_ram_rdata2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[5]
  PIN data_arrays_0_0_ext_ram_rdata2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[60]
  PIN data_arrays_0_0_ext_ram_rdata2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[61]
  PIN data_arrays_0_0_ext_ram_rdata2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1015.280 4.000 1015.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[62]
  PIN data_arrays_0_0_ext_ram_rdata2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.680 4.000 1019.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[63]
  PIN data_arrays_0_0_ext_ram_rdata2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[6]
  PIN data_arrays_0_0_ext_ram_rdata2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 821.480 4.000 822.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[7]
  PIN data_arrays_0_0_ext_ram_rdata2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.880 4.000 825.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[8]
  PIN data_arrays_0_0_ext_ram_rdata2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata2[9]
  PIN data_arrays_0_0_ext_ram_rdata3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1022.080 4.000 1022.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[0]
  PIN data_arrays_0_0_ext_ram_rdata3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[10]
  PIN data_arrays_0_0_ext_ram_rdata3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[11]
  PIN data_arrays_0_0_ext_ram_rdata3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[12]
  PIN data_arrays_0_0_ext_ram_rdata3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1068.320 4.000 1068.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[13]
  PIN data_arrays_0_0_ext_ram_rdata3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.720 4.000 1072.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[14]
  PIN data_arrays_0_0_ext_ram_rdata3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.120 4.000 1075.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[15]
  PIN data_arrays_0_0_ext_ram_rdata3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1078.520 4.000 1079.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[16]
  PIN data_arrays_0_0_ext_ram_rdata3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.920 4.000 1082.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[17]
  PIN data_arrays_0_0_ext_ram_rdata3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1085.320 4.000 1085.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[18]
  PIN data_arrays_0_0_ext_ram_rdata3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1089.400 4.000 1090.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[19]
  PIN data_arrays_0_0_ext_ram_rdata3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[1]
  PIN data_arrays_0_0_ext_ram_rdata3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1092.800 4.000 1093.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[20]
  PIN data_arrays_0_0_ext_ram_rdata3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.200 4.000 1096.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[21]
  PIN data_arrays_0_0_ext_ram_rdata3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[22]
  PIN data_arrays_0_0_ext_ram_rdata3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1103.000 4.000 1103.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[23]
  PIN data_arrays_0_0_ext_ram_rdata3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1106.400 4.000 1107.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[24]
  PIN data_arrays_0_0_ext_ram_rdata3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1110.480 4.000 1111.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[25]
  PIN data_arrays_0_0_ext_ram_rdata3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1113.880 4.000 1114.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[26]
  PIN data_arrays_0_0_ext_ram_rdata3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.280 4.000 1117.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[27]
  PIN data_arrays_0_0_ext_ram_rdata3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.680 4.000 1121.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[28]
  PIN data_arrays_0_0_ext_ram_rdata3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.080 4.000 1124.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[29]
  PIN data_arrays_0_0_ext_ram_rdata3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[2]
  PIN data_arrays_0_0_ext_ram_rdata3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.160 4.000 1128.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[30]
  PIN data_arrays_0_0_ext_ram_rdata3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1131.560 4.000 1132.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[31]
  PIN data_arrays_0_0_ext_ram_rdata3[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1134.960 4.000 1135.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[32]
  PIN data_arrays_0_0_ext_ram_rdata3[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1138.360 4.000 1138.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[33]
  PIN data_arrays_0_0_ext_ram_rdata3[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.760 4.000 1142.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[34]
  PIN data_arrays_0_0_ext_ram_rdata3[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.160 4.000 1145.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[35]
  PIN data_arrays_0_0_ext_ram_rdata3[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[36]
  PIN data_arrays_0_0_ext_ram_rdata3[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[37]
  PIN data_arrays_0_0_ext_ram_rdata3[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[38]
  PIN data_arrays_0_0_ext_ram_rdata3[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[39]
  PIN data_arrays_0_0_ext_ram_rdata3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.960 4.000 1033.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[3]
  PIN data_arrays_0_0_ext_ram_rdata3[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[40]
  PIN data_arrays_0_0_ext_ram_rdata3[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[41]
  PIN data_arrays_0_0_ext_ram_rdata3[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1170.320 4.000 1170.920 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[42]
  PIN data_arrays_0_0_ext_ram_rdata3[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.720 4.000 1174.320 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[43]
  PIN data_arrays_0_0_ext_ram_rdata3[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.120 4.000 1177.720 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[44]
  PIN data_arrays_0_0_ext_ram_rdata3[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1180.520 4.000 1181.120 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[45]
  PIN data_arrays_0_0_ext_ram_rdata3[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.920 4.000 1184.520 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[46]
  PIN data_arrays_0_0_ext_ram_rdata3[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1188.000 4.000 1188.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[47]
  PIN data_arrays_0_0_ext_ram_rdata3[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1191.400 4.000 1192.000 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[48]
  PIN data_arrays_0_0_ext_ram_rdata3[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.800 4.000 1195.400 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[49]
  PIN data_arrays_0_0_ext_ram_rdata3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[4]
  PIN data_arrays_0_0_ext_ram_rdata3[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1198.200 4.000 1198.800 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[50]
  PIN data_arrays_0_0_ext_ram_rdata3[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1201.600 4.000 1202.200 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[51]
  PIN data_arrays_0_0_ext_ram_rdata3[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1205.000 4.000 1205.600 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[52]
  PIN data_arrays_0_0_ext_ram_rdata3[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1209.080 4.000 1209.680 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[53]
  PIN data_arrays_0_0_ext_ram_rdata3[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1212.480 4.000 1213.080 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[54]
  PIN data_arrays_0_0_ext_ram_rdata3[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1215.880 4.000 1216.480 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[55]
  PIN data_arrays_0_0_ext_ram_rdata3[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1219.280 4.000 1219.880 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[56]
  PIN data_arrays_0_0_ext_ram_rdata3[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1222.680 4.000 1223.280 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[57]
  PIN data_arrays_0_0_ext_ram_rdata3[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1226.760 4.000 1227.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[58]
  PIN data_arrays_0_0_ext_ram_rdata3[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.160 4.000 1230.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[59]
  PIN data_arrays_0_0_ext_ram_rdata3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1039.760 4.000 1040.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[5]
  PIN data_arrays_0_0_ext_ram_rdata3[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1233.560 4.000 1234.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[60]
  PIN data_arrays_0_0_ext_ram_rdata3[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.960 4.000 1237.560 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[61]
  PIN data_arrays_0_0_ext_ram_rdata3[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1240.360 4.000 1240.960 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[62]
  PIN data_arrays_0_0_ext_ram_rdata3[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.760 4.000 1244.360 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[63]
  PIN data_arrays_0_0_ext_ram_rdata3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.160 4.000 1043.760 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[6]
  PIN data_arrays_0_0_ext_ram_rdata3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1046.560 4.000 1047.160 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[7]
  PIN data_arrays_0_0_ext_ram_rdata3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[8]
  PIN data_arrays_0_0_ext_ram_rdata3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END data_arrays_0_0_ext_ram_rdata3[9]
  PIN data_arrays_0_0_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[0]
  PIN data_arrays_0_0_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata[10]
  PIN data_arrays_0_0_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata[11]
  PIN data_arrays_0_0_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[12]
  PIN data_arrays_0_0_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 532.480 4.000 533.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[13]
  PIN data_arrays_0_0_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[14]
  PIN data_arrays_0_0_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata[15]
  PIN data_arrays_0_0_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata[16]
  PIN data_arrays_0_0_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata[17]
  PIN data_arrays_0_0_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[18]
  PIN data_arrays_0_0_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[19]
  PIN data_arrays_0_0_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 490.320 4.000 490.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[1]
  PIN data_arrays_0_0_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[20]
  PIN data_arrays_0_0_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata[21]
  PIN data_arrays_0_0_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata[22]
  PIN data_arrays_0_0_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata[23]
  PIN data_arrays_0_0_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata[24]
  PIN data_arrays_0_0_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[25]
  PIN data_arrays_0_0_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[26]
  PIN data_arrays_0_0_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata[27]
  PIN data_arrays_0_0_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[28]
  PIN data_arrays_0_0_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[29]
  PIN data_arrays_0_0_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[2]
  PIN data_arrays_0_0_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[30]
  PIN data_arrays_0_0_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[31]
  PIN data_arrays_0_0_ext_ram_wdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[32]
  PIN data_arrays_0_0_ext_ram_wdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[33]
  PIN data_arrays_0_0_ext_ram_wdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[34]
  PIN data_arrays_0_0_ext_ram_wdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.000 4.000 610.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[35]
  PIN data_arrays_0_0_ext_ram_wdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.080 4.000 614.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[36]
  PIN data_arrays_0_0_ext_ram_wdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[37]
  PIN data_arrays_0_0_ext_ram_wdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.880 4.000 621.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[38]
  PIN data_arrays_0_0_ext_ram_wdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END data_arrays_0_0_ext_ram_wdata[39]
  PIN data_arrays_0_0_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[3]
  PIN data_arrays_0_0_ext_ram_wdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END data_arrays_0_0_ext_ram_wdata[40]
  PIN data_arrays_0_0_ext_ram_wdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END data_arrays_0_0_ext_ram_wdata[41]
  PIN data_arrays_0_0_ext_ram_wdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[42]
  PIN data_arrays_0_0_ext_ram_wdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END data_arrays_0_0_ext_ram_wdata[43]
  PIN data_arrays_0_0_ext_ram_wdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END data_arrays_0_0_ext_ram_wdata[44]
  PIN data_arrays_0_0_ext_ram_wdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 645.360 4.000 645.960 ;
    END
  END data_arrays_0_0_ext_ram_wdata[45]
  PIN data_arrays_0_0_ext_ram_wdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END data_arrays_0_0_ext_ram_wdata[46]
  PIN data_arrays_0_0_ext_ram_wdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END data_arrays_0_0_ext_ram_wdata[47]
  PIN data_arrays_0_0_ext_ram_wdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END data_arrays_0_0_ext_ram_wdata[48]
  PIN data_arrays_0_0_ext_ram_wdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END data_arrays_0_0_ext_ram_wdata[49]
  PIN data_arrays_0_0_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[4]
  PIN data_arrays_0_0_ext_ram_wdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END data_arrays_0_0_ext_ram_wdata[50]
  PIN data_arrays_0_0_ext_ram_wdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END data_arrays_0_0_ext_ram_wdata[51]
  PIN data_arrays_0_0_ext_ram_wdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END data_arrays_0_0_ext_ram_wdata[52]
  PIN data_arrays_0_0_ext_ram_wdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[53]
  PIN data_arrays_0_0_ext_ram_wdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END data_arrays_0_0_ext_ram_wdata[54]
  PIN data_arrays_0_0_ext_ram_wdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END data_arrays_0_0_ext_ram_wdata[55]
  PIN data_arrays_0_0_ext_ram_wdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END data_arrays_0_0_ext_ram_wdata[56]
  PIN data_arrays_0_0_ext_ram_wdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.520 4.000 688.120 ;
    END
  END data_arrays_0_0_ext_ram_wdata[57]
  PIN data_arrays_0_0_ext_ram_wdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END data_arrays_0_0_ext_ram_wdata[58]
  PIN data_arrays_0_0_ext_ram_wdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[59]
  PIN data_arrays_0_0_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[5]
  PIN data_arrays_0_0_ext_ram_wdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 698.400 4.000 699.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[60]
  PIN data_arrays_0_0_ext_ram_wdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END data_arrays_0_0_ext_ram_wdata[61]
  PIN data_arrays_0_0_ext_ram_wdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 4.000 705.800 ;
    END
  END data_arrays_0_0_ext_ram_wdata[62]
  PIN data_arrays_0_0_ext_ram_wdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END data_arrays_0_0_ext_ram_wdata[63]
  PIN data_arrays_0_0_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END data_arrays_0_0_ext_ram_wdata[6]
  PIN data_arrays_0_0_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END data_arrays_0_0_ext_ram_wdata[7]
  PIN data_arrays_0_0_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END data_arrays_0_0_ext_ram_wdata[8]
  PIN data_arrays_0_0_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END data_arrays_0_0_ext_ram_wdata[9]
  PIN data_arrays_0_0_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.760 4.000 734.360 ;
    END
  END data_arrays_0_0_ext_ram_web
  PIN data_arrays_0_0_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END data_arrays_0_0_ext_ram_wmask[0]
  PIN data_arrays_0_0_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END data_arrays_0_0_ext_ram_wmask[1]
  PIN data_arrays_0_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1702.080 1767.395 1702.680 ;
    END
  END data_arrays_0_ext_ram_addr1[0]
  PIN data_arrays_0_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1710.920 1767.395 1711.520 ;
    END
  END data_arrays_0_ext_ram_addr1[1]
  PIN data_arrays_0_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1719.760 1767.395 1720.360 ;
    END
  END data_arrays_0_ext_ram_addr1[2]
  PIN data_arrays_0_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1728.600 1767.395 1729.200 ;
    END
  END data_arrays_0_ext_ram_addr1[3]
  PIN data_arrays_0_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1737.440 1767.395 1738.040 ;
    END
  END data_arrays_0_ext_ram_addr1[4]
  PIN data_arrays_0_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1746.280 1767.395 1746.880 ;
    END
  END data_arrays_0_ext_ram_addr1[5]
  PIN data_arrays_0_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1755.120 1767.395 1755.720 ;
    END
  END data_arrays_0_ext_ram_addr1[6]
  PIN data_arrays_0_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1763.960 1767.395 1764.560 ;
    END
  END data_arrays_0_ext_ram_addr1[7]
  PIN data_arrays_0_ext_ram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1772.800 1767.395 1773.400 ;
    END
  END data_arrays_0_ext_ram_addr1[8]
  PIN data_arrays_0_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1141.760 1767.395 1142.360 ;
    END
  END data_arrays_0_ext_ram_addr[0]
  PIN data_arrays_0_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1150.600 1767.395 1151.200 ;
    END
  END data_arrays_0_ext_ram_addr[1]
  PIN data_arrays_0_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1159.440 1767.395 1160.040 ;
    END
  END data_arrays_0_ext_ram_addr[2]
  PIN data_arrays_0_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1168.280 1767.395 1168.880 ;
    END
  END data_arrays_0_ext_ram_addr[3]
  PIN data_arrays_0_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1177.120 1767.395 1177.720 ;
    END
  END data_arrays_0_ext_ram_addr[4]
  PIN data_arrays_0_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1185.960 1767.395 1186.560 ;
    END
  END data_arrays_0_ext_ram_addr[5]
  PIN data_arrays_0_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1195.480 1767.395 1196.080 ;
    END
  END data_arrays_0_ext_ram_addr[6]
  PIN data_arrays_0_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1204.320 1767.395 1204.920 ;
    END
  END data_arrays_0_ext_ram_addr[7]
  PIN data_arrays_0_ext_ram_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1213.160 1767.395 1213.760 ;
    END
  END data_arrays_0_ext_ram_addr[8]
  PIN data_arrays_0_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1222.000 1767.395 1222.600 ;
    END
  END data_arrays_0_ext_ram_clk
  PIN data_arrays_0_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1630.680 1767.395 1631.280 ;
    END
  END data_arrays_0_ext_ram_csb1[0]
  PIN data_arrays_0_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1639.520 1767.395 1640.120 ;
    END
  END data_arrays_0_ext_ram_csb1[1]
  PIN data_arrays_0_ext_ram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1648.360 1767.395 1648.960 ;
    END
  END data_arrays_0_ext_ram_csb1[2]
  PIN data_arrays_0_ext_ram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1657.200 1767.395 1657.800 ;
    END
  END data_arrays_0_ext_ram_csb1[3]
  PIN data_arrays_0_ext_ram_csb1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1666.720 1767.395 1667.320 ;
    END
  END data_arrays_0_ext_ram_csb1[4]
  PIN data_arrays_0_ext_ram_csb1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1675.560 1767.395 1676.160 ;
    END
  END data_arrays_0_ext_ram_csb1[5]
  PIN data_arrays_0_ext_ram_csb1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1684.400 1767.395 1685.000 ;
    END
  END data_arrays_0_ext_ram_csb1[6]
  PIN data_arrays_0_ext_ram_csb1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1693.240 1767.395 1693.840 ;
    END
  END data_arrays_0_ext_ram_csb1[7]
  PIN data_arrays_0_ext_ram_csb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1551.120 1767.395 1551.720 ;
    END
  END data_arrays_0_ext_ram_csb[0]
  PIN data_arrays_0_ext_ram_csb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1559.960 1767.395 1560.560 ;
    END
  END data_arrays_0_ext_ram_csb[1]
  PIN data_arrays_0_ext_ram_csb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1568.800 1767.395 1569.400 ;
    END
  END data_arrays_0_ext_ram_csb[2]
  PIN data_arrays_0_ext_ram_csb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1577.640 1767.395 1578.240 ;
    END
  END data_arrays_0_ext_ram_csb[3]
  PIN data_arrays_0_ext_ram_csb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1586.480 1767.395 1587.080 ;
    END
  END data_arrays_0_ext_ram_csb[4]
  PIN data_arrays_0_ext_ram_csb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1595.320 1767.395 1595.920 ;
    END
  END data_arrays_0_ext_ram_csb[5]
  PIN data_arrays_0_ext_ram_csb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1604.160 1767.395 1604.760 ;
    END
  END data_arrays_0_ext_ram_csb[6]
  PIN data_arrays_0_ext_ram_csb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1613.000 1767.395 1613.600 ;
    END
  END data_arrays_0_ext_ram_csb[7]
  PIN data_arrays_0_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 4.120 1767.395 4.720 ;
    END
  END data_arrays_0_ext_ram_rdata0[0]
  PIN data_arrays_0_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 92.520 1767.395 93.120 ;
    END
  END data_arrays_0_ext_ram_rdata0[10]
  PIN data_arrays_0_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 101.360 1767.395 101.960 ;
    END
  END data_arrays_0_ext_ram_rdata0[11]
  PIN data_arrays_0_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 110.200 1767.395 110.800 ;
    END
  END data_arrays_0_ext_ram_rdata0[12]
  PIN data_arrays_0_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 119.040 1767.395 119.640 ;
    END
  END data_arrays_0_ext_ram_rdata0[13]
  PIN data_arrays_0_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 128.560 1767.395 129.160 ;
    END
  END data_arrays_0_ext_ram_rdata0[14]
  PIN data_arrays_0_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 137.400 1767.395 138.000 ;
    END
  END data_arrays_0_ext_ram_rdata0[15]
  PIN data_arrays_0_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 146.240 1767.395 146.840 ;
    END
  END data_arrays_0_ext_ram_rdata0[16]
  PIN data_arrays_0_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 155.080 1767.395 155.680 ;
    END
  END data_arrays_0_ext_ram_rdata0[17]
  PIN data_arrays_0_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 163.920 1767.395 164.520 ;
    END
  END data_arrays_0_ext_ram_rdata0[18]
  PIN data_arrays_0_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 172.760 1767.395 173.360 ;
    END
  END data_arrays_0_ext_ram_rdata0[19]
  PIN data_arrays_0_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 12.960 1767.395 13.560 ;
    END
  END data_arrays_0_ext_ram_rdata0[1]
  PIN data_arrays_0_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 181.600 1767.395 182.200 ;
    END
  END data_arrays_0_ext_ram_rdata0[20]
  PIN data_arrays_0_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 190.440 1767.395 191.040 ;
    END
  END data_arrays_0_ext_ram_rdata0[21]
  PIN data_arrays_0_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 199.280 1767.395 199.880 ;
    END
  END data_arrays_0_ext_ram_rdata0[22]
  PIN data_arrays_0_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 208.120 1767.395 208.720 ;
    END
  END data_arrays_0_ext_ram_rdata0[23]
  PIN data_arrays_0_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 216.960 1767.395 217.560 ;
    END
  END data_arrays_0_ext_ram_rdata0[24]
  PIN data_arrays_0_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 225.800 1767.395 226.400 ;
    END
  END data_arrays_0_ext_ram_rdata0[25]
  PIN data_arrays_0_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 234.640 1767.395 235.240 ;
    END
  END data_arrays_0_ext_ram_rdata0[26]
  PIN data_arrays_0_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 244.160 1767.395 244.760 ;
    END
  END data_arrays_0_ext_ram_rdata0[27]
  PIN data_arrays_0_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 253.000 1767.395 253.600 ;
    END
  END data_arrays_0_ext_ram_rdata0[28]
  PIN data_arrays_0_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 261.840 1767.395 262.440 ;
    END
  END data_arrays_0_ext_ram_rdata0[29]
  PIN data_arrays_0_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 21.800 1767.395 22.400 ;
    END
  END data_arrays_0_ext_ram_rdata0[2]
  PIN data_arrays_0_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 270.680 1767.395 271.280 ;
    END
  END data_arrays_0_ext_ram_rdata0[30]
  PIN data_arrays_0_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 279.520 1767.395 280.120 ;
    END
  END data_arrays_0_ext_ram_rdata0[31]
  PIN data_arrays_0_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 30.640 1767.395 31.240 ;
    END
  END data_arrays_0_ext_ram_rdata0[3]
  PIN data_arrays_0_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 39.480 1767.395 40.080 ;
    END
  END data_arrays_0_ext_ram_rdata0[4]
  PIN data_arrays_0_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 48.320 1767.395 48.920 ;
    END
  END data_arrays_0_ext_ram_rdata0[5]
  PIN data_arrays_0_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 57.160 1767.395 57.760 ;
    END
  END data_arrays_0_ext_ram_rdata0[6]
  PIN data_arrays_0_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 66.000 1767.395 66.600 ;
    END
  END data_arrays_0_ext_ram_rdata0[7]
  PIN data_arrays_0_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 74.840 1767.395 75.440 ;
    END
  END data_arrays_0_ext_ram_rdata0[8]
  PIN data_arrays_0_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 83.680 1767.395 84.280 ;
    END
  END data_arrays_0_ext_ram_rdata0[9]
  PIN data_arrays_0_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 288.360 1767.395 288.960 ;
    END
  END data_arrays_0_ext_ram_rdata1[0]
  PIN data_arrays_0_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 377.440 1767.395 378.040 ;
    END
  END data_arrays_0_ext_ram_rdata1[10]
  PIN data_arrays_0_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 386.280 1767.395 386.880 ;
    END
  END data_arrays_0_ext_ram_rdata1[11]
  PIN data_arrays_0_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 395.120 1767.395 395.720 ;
    END
  END data_arrays_0_ext_ram_rdata1[12]
  PIN data_arrays_0_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 403.960 1767.395 404.560 ;
    END
  END data_arrays_0_ext_ram_rdata1[13]
  PIN data_arrays_0_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 412.800 1767.395 413.400 ;
    END
  END data_arrays_0_ext_ram_rdata1[14]
  PIN data_arrays_0_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 421.640 1767.395 422.240 ;
    END
  END data_arrays_0_ext_ram_rdata1[15]
  PIN data_arrays_0_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 430.480 1767.395 431.080 ;
    END
  END data_arrays_0_ext_ram_rdata1[16]
  PIN data_arrays_0_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 439.320 1767.395 439.920 ;
    END
  END data_arrays_0_ext_ram_rdata1[17]
  PIN data_arrays_0_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 448.160 1767.395 448.760 ;
    END
  END data_arrays_0_ext_ram_rdata1[18]
  PIN data_arrays_0_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 457.000 1767.395 457.600 ;
    END
  END data_arrays_0_ext_ram_rdata1[19]
  PIN data_arrays_0_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 297.200 1767.395 297.800 ;
    END
  END data_arrays_0_ext_ram_rdata1[1]
  PIN data_arrays_0_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 465.840 1767.395 466.440 ;
    END
  END data_arrays_0_ext_ram_rdata1[20]
  PIN data_arrays_0_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 474.680 1767.395 475.280 ;
    END
  END data_arrays_0_ext_ram_rdata1[21]
  PIN data_arrays_0_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 484.200 1767.395 484.800 ;
    END
  END data_arrays_0_ext_ram_rdata1[22]
  PIN data_arrays_0_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 493.040 1767.395 493.640 ;
    END
  END data_arrays_0_ext_ram_rdata1[23]
  PIN data_arrays_0_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 501.880 1767.395 502.480 ;
    END
  END data_arrays_0_ext_ram_rdata1[24]
  PIN data_arrays_0_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 510.720 1767.395 511.320 ;
    END
  END data_arrays_0_ext_ram_rdata1[25]
  PIN data_arrays_0_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 519.560 1767.395 520.160 ;
    END
  END data_arrays_0_ext_ram_rdata1[26]
  PIN data_arrays_0_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 528.400 1767.395 529.000 ;
    END
  END data_arrays_0_ext_ram_rdata1[27]
  PIN data_arrays_0_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 537.240 1767.395 537.840 ;
    END
  END data_arrays_0_ext_ram_rdata1[28]
  PIN data_arrays_0_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 546.080 1767.395 546.680 ;
    END
  END data_arrays_0_ext_ram_rdata1[29]
  PIN data_arrays_0_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 306.040 1767.395 306.640 ;
    END
  END data_arrays_0_ext_ram_rdata1[2]
  PIN data_arrays_0_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 554.920 1767.395 555.520 ;
    END
  END data_arrays_0_ext_ram_rdata1[30]
  PIN data_arrays_0_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 563.760 1767.395 564.360 ;
    END
  END data_arrays_0_ext_ram_rdata1[31]
  PIN data_arrays_0_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 314.880 1767.395 315.480 ;
    END
  END data_arrays_0_ext_ram_rdata1[3]
  PIN data_arrays_0_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 323.720 1767.395 324.320 ;
    END
  END data_arrays_0_ext_ram_rdata1[4]
  PIN data_arrays_0_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 332.560 1767.395 333.160 ;
    END
  END data_arrays_0_ext_ram_rdata1[5]
  PIN data_arrays_0_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 341.400 1767.395 342.000 ;
    END
  END data_arrays_0_ext_ram_rdata1[6]
  PIN data_arrays_0_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 350.240 1767.395 350.840 ;
    END
  END data_arrays_0_ext_ram_rdata1[7]
  PIN data_arrays_0_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 359.760 1767.395 360.360 ;
    END
  END data_arrays_0_ext_ram_rdata1[8]
  PIN data_arrays_0_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 368.600 1767.395 369.200 ;
    END
  END data_arrays_0_ext_ram_rdata1[9]
  PIN data_arrays_0_ext_ram_rdata2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 572.600 1767.395 573.200 ;
    END
  END data_arrays_0_ext_ram_rdata2[0]
  PIN data_arrays_0_ext_ram_rdata2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 661.680 1767.395 662.280 ;
    END
  END data_arrays_0_ext_ram_rdata2[10]
  PIN data_arrays_0_ext_ram_rdata2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 670.520 1767.395 671.120 ;
    END
  END data_arrays_0_ext_ram_rdata2[11]
  PIN data_arrays_0_ext_ram_rdata2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 679.360 1767.395 679.960 ;
    END
  END data_arrays_0_ext_ram_rdata2[12]
  PIN data_arrays_0_ext_ram_rdata2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 688.200 1767.395 688.800 ;
    END
  END data_arrays_0_ext_ram_rdata2[13]
  PIN data_arrays_0_ext_ram_rdata2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 697.040 1767.395 697.640 ;
    END
  END data_arrays_0_ext_ram_rdata2[14]
  PIN data_arrays_0_ext_ram_rdata2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 705.880 1767.395 706.480 ;
    END
  END data_arrays_0_ext_ram_rdata2[15]
  PIN data_arrays_0_ext_ram_rdata2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 715.400 1767.395 716.000 ;
    END
  END data_arrays_0_ext_ram_rdata2[16]
  PIN data_arrays_0_ext_ram_rdata2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 724.240 1767.395 724.840 ;
    END
  END data_arrays_0_ext_ram_rdata2[17]
  PIN data_arrays_0_ext_ram_rdata2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 733.080 1767.395 733.680 ;
    END
  END data_arrays_0_ext_ram_rdata2[18]
  PIN data_arrays_0_ext_ram_rdata2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 741.920 1767.395 742.520 ;
    END
  END data_arrays_0_ext_ram_rdata2[19]
  PIN data_arrays_0_ext_ram_rdata2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 581.440 1767.395 582.040 ;
    END
  END data_arrays_0_ext_ram_rdata2[1]
  PIN data_arrays_0_ext_ram_rdata2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 750.760 1767.395 751.360 ;
    END
  END data_arrays_0_ext_ram_rdata2[20]
  PIN data_arrays_0_ext_ram_rdata2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 759.600 1767.395 760.200 ;
    END
  END data_arrays_0_ext_ram_rdata2[21]
  PIN data_arrays_0_ext_ram_rdata2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 768.440 1767.395 769.040 ;
    END
  END data_arrays_0_ext_ram_rdata2[22]
  PIN data_arrays_0_ext_ram_rdata2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 777.280 1767.395 777.880 ;
    END
  END data_arrays_0_ext_ram_rdata2[23]
  PIN data_arrays_0_ext_ram_rdata2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 786.120 1767.395 786.720 ;
    END
  END data_arrays_0_ext_ram_rdata2[24]
  PIN data_arrays_0_ext_ram_rdata2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 794.960 1767.395 795.560 ;
    END
  END data_arrays_0_ext_ram_rdata2[25]
  PIN data_arrays_0_ext_ram_rdata2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 803.800 1767.395 804.400 ;
    END
  END data_arrays_0_ext_ram_rdata2[26]
  PIN data_arrays_0_ext_ram_rdata2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 812.640 1767.395 813.240 ;
    END
  END data_arrays_0_ext_ram_rdata2[27]
  PIN data_arrays_0_ext_ram_rdata2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 821.480 1767.395 822.080 ;
    END
  END data_arrays_0_ext_ram_rdata2[28]
  PIN data_arrays_0_ext_ram_rdata2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 830.320 1767.395 830.920 ;
    END
  END data_arrays_0_ext_ram_rdata2[29]
  PIN data_arrays_0_ext_ram_rdata2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 590.280 1767.395 590.880 ;
    END
  END data_arrays_0_ext_ram_rdata2[2]
  PIN data_arrays_0_ext_ram_rdata2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 839.840 1767.395 840.440 ;
    END
  END data_arrays_0_ext_ram_rdata2[30]
  PIN data_arrays_0_ext_ram_rdata2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 848.680 1767.395 849.280 ;
    END
  END data_arrays_0_ext_ram_rdata2[31]
  PIN data_arrays_0_ext_ram_rdata2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 599.800 1767.395 600.400 ;
    END
  END data_arrays_0_ext_ram_rdata2[3]
  PIN data_arrays_0_ext_ram_rdata2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 608.640 1767.395 609.240 ;
    END
  END data_arrays_0_ext_ram_rdata2[4]
  PIN data_arrays_0_ext_ram_rdata2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 617.480 1767.395 618.080 ;
    END
  END data_arrays_0_ext_ram_rdata2[5]
  PIN data_arrays_0_ext_ram_rdata2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 626.320 1767.395 626.920 ;
    END
  END data_arrays_0_ext_ram_rdata2[6]
  PIN data_arrays_0_ext_ram_rdata2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 635.160 1767.395 635.760 ;
    END
  END data_arrays_0_ext_ram_rdata2[7]
  PIN data_arrays_0_ext_ram_rdata2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 644.000 1767.395 644.600 ;
    END
  END data_arrays_0_ext_ram_rdata2[8]
  PIN data_arrays_0_ext_ram_rdata2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 652.840 1767.395 653.440 ;
    END
  END data_arrays_0_ext_ram_rdata2[9]
  PIN data_arrays_0_ext_ram_rdata3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 857.520 1767.395 858.120 ;
    END
  END data_arrays_0_ext_ram_rdata3[0]
  PIN data_arrays_0_ext_ram_rdata3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 945.920 1767.395 946.520 ;
    END
  END data_arrays_0_ext_ram_rdata3[10]
  PIN data_arrays_0_ext_ram_rdata3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 955.440 1767.395 956.040 ;
    END
  END data_arrays_0_ext_ram_rdata3[11]
  PIN data_arrays_0_ext_ram_rdata3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 964.280 1767.395 964.880 ;
    END
  END data_arrays_0_ext_ram_rdata3[12]
  PIN data_arrays_0_ext_ram_rdata3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 973.120 1767.395 973.720 ;
    END
  END data_arrays_0_ext_ram_rdata3[13]
  PIN data_arrays_0_ext_ram_rdata3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 981.960 1767.395 982.560 ;
    END
  END data_arrays_0_ext_ram_rdata3[14]
  PIN data_arrays_0_ext_ram_rdata3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 990.800 1767.395 991.400 ;
    END
  END data_arrays_0_ext_ram_rdata3[15]
  PIN data_arrays_0_ext_ram_rdata3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 999.640 1767.395 1000.240 ;
    END
  END data_arrays_0_ext_ram_rdata3[16]
  PIN data_arrays_0_ext_ram_rdata3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1008.480 1767.395 1009.080 ;
    END
  END data_arrays_0_ext_ram_rdata3[17]
  PIN data_arrays_0_ext_ram_rdata3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1017.320 1767.395 1017.920 ;
    END
  END data_arrays_0_ext_ram_rdata3[18]
  PIN data_arrays_0_ext_ram_rdata3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1026.160 1767.395 1026.760 ;
    END
  END data_arrays_0_ext_ram_rdata3[19]
  PIN data_arrays_0_ext_ram_rdata3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 866.360 1767.395 866.960 ;
    END
  END data_arrays_0_ext_ram_rdata3[1]
  PIN data_arrays_0_ext_ram_rdata3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1035.000 1767.395 1035.600 ;
    END
  END data_arrays_0_ext_ram_rdata3[20]
  PIN data_arrays_0_ext_ram_rdata3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1043.840 1767.395 1044.440 ;
    END
  END data_arrays_0_ext_ram_rdata3[21]
  PIN data_arrays_0_ext_ram_rdata3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1052.680 1767.395 1053.280 ;
    END
  END data_arrays_0_ext_ram_rdata3[22]
  PIN data_arrays_0_ext_ram_rdata3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1061.520 1767.395 1062.120 ;
    END
  END data_arrays_0_ext_ram_rdata3[23]
  PIN data_arrays_0_ext_ram_rdata3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1071.040 1767.395 1071.640 ;
    END
  END data_arrays_0_ext_ram_rdata3[24]
  PIN data_arrays_0_ext_ram_rdata3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1079.880 1767.395 1080.480 ;
    END
  END data_arrays_0_ext_ram_rdata3[25]
  PIN data_arrays_0_ext_ram_rdata3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1088.720 1767.395 1089.320 ;
    END
  END data_arrays_0_ext_ram_rdata3[26]
  PIN data_arrays_0_ext_ram_rdata3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1097.560 1767.395 1098.160 ;
    END
  END data_arrays_0_ext_ram_rdata3[27]
  PIN data_arrays_0_ext_ram_rdata3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1106.400 1767.395 1107.000 ;
    END
  END data_arrays_0_ext_ram_rdata3[28]
  PIN data_arrays_0_ext_ram_rdata3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1115.240 1767.395 1115.840 ;
    END
  END data_arrays_0_ext_ram_rdata3[29]
  PIN data_arrays_0_ext_ram_rdata3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 875.200 1767.395 875.800 ;
    END
  END data_arrays_0_ext_ram_rdata3[2]
  PIN data_arrays_0_ext_ram_rdata3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1124.080 1767.395 1124.680 ;
    END
  END data_arrays_0_ext_ram_rdata3[30]
  PIN data_arrays_0_ext_ram_rdata3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1132.920 1767.395 1133.520 ;
    END
  END data_arrays_0_ext_ram_rdata3[31]
  PIN data_arrays_0_ext_ram_rdata3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 884.040 1767.395 884.640 ;
    END
  END data_arrays_0_ext_ram_rdata3[3]
  PIN data_arrays_0_ext_ram_rdata3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 892.880 1767.395 893.480 ;
    END
  END data_arrays_0_ext_ram_rdata3[4]
  PIN data_arrays_0_ext_ram_rdata3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 901.720 1767.395 902.320 ;
    END
  END data_arrays_0_ext_ram_rdata3[5]
  PIN data_arrays_0_ext_ram_rdata3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 910.560 1767.395 911.160 ;
    END
  END data_arrays_0_ext_ram_rdata3[6]
  PIN data_arrays_0_ext_ram_rdata3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 919.400 1767.395 920.000 ;
    END
  END data_arrays_0_ext_ram_rdata3[7]
  PIN data_arrays_0_ext_ram_rdata3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 928.240 1767.395 928.840 ;
    END
  END data_arrays_0_ext_ram_rdata3[8]
  PIN data_arrays_0_ext_ram_rdata3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 937.080 1767.395 937.680 ;
    END
  END data_arrays_0_ext_ram_rdata3[9]
  PIN data_arrays_0_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1230.840 1767.395 1231.440 ;
    END
  END data_arrays_0_ext_ram_wdata[0]
  PIN data_arrays_0_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1319.920 1767.395 1320.520 ;
    END
  END data_arrays_0_ext_ram_wdata[10]
  PIN data_arrays_0_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1328.760 1767.395 1329.360 ;
    END
  END data_arrays_0_ext_ram_wdata[11]
  PIN data_arrays_0_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1337.600 1767.395 1338.200 ;
    END
  END data_arrays_0_ext_ram_wdata[12]
  PIN data_arrays_0_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1346.440 1767.395 1347.040 ;
    END
  END data_arrays_0_ext_ram_wdata[13]
  PIN data_arrays_0_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1355.280 1767.395 1355.880 ;
    END
  END data_arrays_0_ext_ram_wdata[14]
  PIN data_arrays_0_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1364.120 1767.395 1364.720 ;
    END
  END data_arrays_0_ext_ram_wdata[15]
  PIN data_arrays_0_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1372.960 1767.395 1373.560 ;
    END
  END data_arrays_0_ext_ram_wdata[16]
  PIN data_arrays_0_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1381.800 1767.395 1382.400 ;
    END
  END data_arrays_0_ext_ram_wdata[17]
  PIN data_arrays_0_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1390.640 1767.395 1391.240 ;
    END
  END data_arrays_0_ext_ram_wdata[18]
  PIN data_arrays_0_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1399.480 1767.395 1400.080 ;
    END
  END data_arrays_0_ext_ram_wdata[19]
  PIN data_arrays_0_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1239.680 1767.395 1240.280 ;
    END
  END data_arrays_0_ext_ram_wdata[1]
  PIN data_arrays_0_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1408.320 1767.395 1408.920 ;
    END
  END data_arrays_0_ext_ram_wdata[20]
  PIN data_arrays_0_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1417.160 1767.395 1417.760 ;
    END
  END data_arrays_0_ext_ram_wdata[21]
  PIN data_arrays_0_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1426.680 1767.395 1427.280 ;
    END
  END data_arrays_0_ext_ram_wdata[22]
  PIN data_arrays_0_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1435.520 1767.395 1436.120 ;
    END
  END data_arrays_0_ext_ram_wdata[23]
  PIN data_arrays_0_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1444.360 1767.395 1444.960 ;
    END
  END data_arrays_0_ext_ram_wdata[24]
  PIN data_arrays_0_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1453.200 1767.395 1453.800 ;
    END
  END data_arrays_0_ext_ram_wdata[25]
  PIN data_arrays_0_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1462.040 1767.395 1462.640 ;
    END
  END data_arrays_0_ext_ram_wdata[26]
  PIN data_arrays_0_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1470.880 1767.395 1471.480 ;
    END
  END data_arrays_0_ext_ram_wdata[27]
  PIN data_arrays_0_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1479.720 1767.395 1480.320 ;
    END
  END data_arrays_0_ext_ram_wdata[28]
  PIN data_arrays_0_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1488.560 1767.395 1489.160 ;
    END
  END data_arrays_0_ext_ram_wdata[29]
  PIN data_arrays_0_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1248.520 1767.395 1249.120 ;
    END
  END data_arrays_0_ext_ram_wdata[2]
  PIN data_arrays_0_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1497.400 1767.395 1498.000 ;
    END
  END data_arrays_0_ext_ram_wdata[30]
  PIN data_arrays_0_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1506.240 1767.395 1506.840 ;
    END
  END data_arrays_0_ext_ram_wdata[31]
  PIN data_arrays_0_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1257.360 1767.395 1257.960 ;
    END
  END data_arrays_0_ext_ram_wdata[3]
  PIN data_arrays_0_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1266.200 1767.395 1266.800 ;
    END
  END data_arrays_0_ext_ram_wdata[4]
  PIN data_arrays_0_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1275.040 1767.395 1275.640 ;
    END
  END data_arrays_0_ext_ram_wdata[5]
  PIN data_arrays_0_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1283.880 1767.395 1284.480 ;
    END
  END data_arrays_0_ext_ram_wdata[6]
  PIN data_arrays_0_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1292.720 1767.395 1293.320 ;
    END
  END data_arrays_0_ext_ram_wdata[7]
  PIN data_arrays_0_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1301.560 1767.395 1302.160 ;
    END
  END data_arrays_0_ext_ram_wdata[8]
  PIN data_arrays_0_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1311.080 1767.395 1311.680 ;
    END
  END data_arrays_0_ext_ram_wdata[9]
  PIN data_arrays_0_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1621.840 1767.395 1622.440 ;
    END
  END data_arrays_0_ext_ram_web
  PIN data_arrays_0_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1515.080 1767.395 1515.680 ;
    END
  END data_arrays_0_ext_ram_wmask[0]
  PIN data_arrays_0_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1523.920 1767.395 1524.520 ;
    END
  END data_arrays_0_ext_ram_wmask[1]
  PIN data_arrays_0_ext_ram_wmask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1532.760 1767.395 1533.360 ;
    END
  END data_arrays_0_ext_ram_wmask[2]
  PIN data_arrays_0_ext_ram_wmask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1763.395 1541.600 1767.395 1542.200 ;
    END
  END data_arrays_0_ext_ram_wmask[3]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 1774.115 7.730 1778.115 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 1774.115 472.790 1778.115 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 1774.115 519.250 1778.115 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 1774.115 565.710 1778.115 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1774.115 612.170 1778.115 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 1774.115 658.630 1778.115 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 1774.115 705.090 1778.115 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 1774.115 751.550 1778.115 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 1774.115 798.010 1778.115 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 1774.115 844.470 1778.115 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 1774.115 891.390 1778.115 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 1774.115 54.190 1778.115 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 1774.115 937.850 1778.115 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 1774.115 984.310 1778.115 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 1774.115 1030.770 1778.115 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 1774.115 1077.230 1778.115 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.410 1774.115 1123.690 1778.115 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 1774.115 1170.150 1778.115 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.330 1774.115 1216.610 1778.115 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.790 1774.115 1263.070 1778.115 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.250 1774.115 1309.530 1778.115 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.170 1774.115 1356.450 1778.115 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 1774.115 100.650 1778.115 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.630 1774.115 1402.910 1778.115 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 1774.115 1449.370 1778.115 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.550 1774.115 1495.830 1778.115 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.010 1774.115 1542.290 1778.115 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.470 1774.115 1588.750 1778.115 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.930 1774.115 1635.210 1778.115 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.390 1774.115 1681.670 1778.115 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.850 1774.115 1728.130 1778.115 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 1774.115 147.110 1778.115 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1774.115 193.570 1778.115 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 1774.115 240.030 1778.115 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 1774.115 286.490 1778.115 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 1774.115 332.950 1778.115 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 1774.115 379.410 1778.115 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 1774.115 425.870 1778.115 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1774.115 22.910 1778.115 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 1774.115 487.970 1778.115 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 1774.115 534.430 1778.115 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 1774.115 580.890 1778.115 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 1774.115 627.810 1778.115 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 1774.115 674.270 1778.115 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 1774.115 720.730 1778.115 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 1774.115 767.190 1778.115 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 1774.115 813.650 1778.115 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 1774.115 860.110 1778.115 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.290 1774.115 906.570 1778.115 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 1774.115 69.370 1778.115 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 1774.115 953.030 1778.115 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 1774.115 999.490 1778.115 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 1774.115 1046.410 1778.115 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 1774.115 1092.870 1778.115 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.050 1774.115 1139.330 1778.115 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.510 1774.115 1185.790 1778.115 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.970 1774.115 1232.250 1778.115 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 1774.115 1278.710 1778.115 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.890 1774.115 1325.170 1778.115 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.350 1774.115 1371.630 1778.115 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 1774.115 115.830 1778.115 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.810 1774.115 1418.090 1778.115 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 1774.115 1464.550 1778.115 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.190 1774.115 1511.470 1778.115 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.650 1774.115 1557.930 1778.115 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.110 1774.115 1604.390 1778.115 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.570 1774.115 1650.850 1778.115 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.030 1774.115 1697.310 1778.115 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.490 1774.115 1743.770 1778.115 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 1774.115 162.750 1778.115 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 1774.115 209.210 1778.115 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 1774.115 255.670 1778.115 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 1774.115 302.130 1778.115 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 1774.115 348.590 1778.115 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 1774.115 395.050 1778.115 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 1774.115 441.510 1778.115 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 1774.115 38.550 1778.115 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 1774.115 503.610 1778.115 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 1774.115 550.070 1778.115 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 1774.115 596.530 1778.115 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 1774.115 642.990 1778.115 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1774.115 689.450 1778.115 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 1774.115 735.910 1778.115 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 1774.115 782.830 1778.115 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 1774.115 829.290 1778.115 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.470 1774.115 875.750 1778.115 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 1774.115 922.210 1778.115 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 1774.115 85.010 1778.115 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 1774.115 968.670 1778.115 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.850 1774.115 1015.130 1778.115 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 1774.115 1061.590 1778.115 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 1774.115 1108.050 1778.115 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.230 1774.115 1154.510 1778.115 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 1774.115 1201.430 1778.115 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 1774.115 1247.890 1778.115 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.070 1774.115 1294.350 1778.115 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.530 1774.115 1340.810 1778.115 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.990 1774.115 1387.270 1778.115 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 1774.115 131.470 1778.115 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.450 1774.115 1433.730 1778.115 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.910 1774.115 1480.190 1778.115 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 1774.115 1526.650 1778.115 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.830 1774.115 1573.110 1778.115 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.290 1774.115 1619.570 1778.115 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.210 1774.115 1666.490 1778.115 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.670 1774.115 1712.950 1778.115 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1759.130 1774.115 1759.410 1778.115 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 1774.115 177.930 1778.115 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 1774.115 224.390 1778.115 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 1774.115 270.850 1778.115 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 1774.115 317.770 1778.115 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1774.115 364.230 1778.115 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 1774.115 410.690 1778.115 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 1774.115 457.150 1778.115 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.750 0.000 1758.030 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 0.000 1761.710 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.110 0.000 1765.390 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.910 0.000 1457.190 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.490 0.000 1467.770 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 0.000 1478.350 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 0.000 1489.390 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 0.000 1499.970 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.310 0.000 1521.590 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.890 0.000 1532.170 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 0.000 1543.210 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.510 0.000 1553.790 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.090 0.000 1564.370 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.130 0.000 1575.410 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.710 0.000 1585.990 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.290 0.000 1596.570 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.330 0.000 1607.610 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.910 0.000 1618.190 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.950 0.000 1629.230 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.530 0.000 1639.810 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 0.000 1650.390 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.150 0.000 1661.430 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.730 0.000 1672.010 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.310 0.000 1682.590 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.350 0.000 1693.630 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.930 0.000 1704.210 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.970 0.000 1715.250 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.550 0.000 1725.830 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.130 0.000 1736.410 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 0.000 1747.450 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 0.000 510.510 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 0.000 725.790 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 0.000 746.950 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 0.000 757.990 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 0.000 800.770 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 0.000 854.590 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 0.000 865.630 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.170 0.000 919.450 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 0.000 930.030 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 0.000 951.650 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 0.000 962.230 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 0.000 983.850 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 0.000 994.430 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 0.000 1016.050 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 0.000 1026.630 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 0.000 1048.250 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 0.000 1058.830 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.170 0.000 1080.450 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 0.000 1102.070 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.370 0.000 1112.650 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.410 0.000 1123.690 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.990 0.000 1134.270 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.610 0.000 1155.890 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.190 0.000 1166.470 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 0.000 1177.510 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 0.000 1188.090 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 0.000 1198.670 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.430 0.000 1209.710 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.010 0.000 1220.290 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 0.000 1231.330 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.630 0.000 1241.910 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.210 0.000 1252.490 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.250 0.000 1263.530 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 0.000 1274.110 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.410 0.000 1284.690 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.450 0.000 1295.730 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.030 0.000 1306.310 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.650 0.000 1327.930 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.230 0.000 1338.510 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.850 0.000 1360.130 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 0.000 1370.710 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 0.000 1381.750 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.050 0.000 1392.330 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 0.000 1403.370 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.250 0.000 1424.530 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 0.000 1435.570 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 0.000 1446.150 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.130 0.000 1460.410 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.170 0.000 1471.450 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.750 0.000 1482.030 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.330 0.000 1492.610 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.370 0.000 1503.650 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.950 0.000 1514.230 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.990 0.000 1525.270 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.570 0.000 1535.850 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.150 0.000 1546.430 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 0.000 1557.470 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.770 0.000 1568.050 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.350 0.000 1578.630 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.390 0.000 1589.670 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.970 0.000 1600.250 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.010 0.000 1611.290 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.590 0.000 1621.870 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.170 0.000 1632.450 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.210 0.000 1643.490 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.790 0.000 1654.070 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.830 0.000 1665.110 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.410 0.000 1675.690 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.990 0.000 1686.270 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.030 0.000 1697.310 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1707.610 0.000 1707.890 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 0.000 1718.470 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 0.000 1729.510 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.810 0.000 1740.090 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.850 0.000 1751.130 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 0.000 675.650 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 0.000 696.810 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 0.000 826.070 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 0.000 836.650 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 0.000 847.690 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 0.000 858.270 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 0.000 868.850 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 0.000 912.090 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 0.000 922.670 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 0.000 933.710 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.590 0.000 954.870 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.630 0.000 965.910 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 0.000 998.110 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 0.000 1008.690 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.450 0.000 1019.730 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.030 0.000 1030.310 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.070 0.000 1041.350 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 0.000 1051.930 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.230 0.000 1062.510 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 0.000 1073.550 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.850 0.000 1084.130 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.430 0.000 1094.710 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.470 0.000 1105.750 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.050 0.000 1116.330 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.670 0.000 1137.950 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.250 0.000 1148.530 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 0.000 1170.150 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.450 0.000 1180.730 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 0.000 1191.770 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 0.000 1202.350 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.110 0.000 1213.390 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.270 0.000 1234.550 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.310 0.000 1245.590 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.470 0.000 1266.750 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 0.000 1277.790 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 0.000 1309.990 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 0.000 1320.570 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.330 0.000 1331.610 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.910 0.000 1342.190 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.530 0.000 1363.810 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.110 0.000 1374.390 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.730 0.000 1396.010 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.310 0.000 1406.590 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 0.000 1417.630 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.930 0.000 1428.210 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.970 0.000 1439.250 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.550 0.000 1449.830 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.810 0.000 1464.090 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.390 0.000 1474.670 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.430 0.000 1485.710 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.010 0.000 1496.290 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 0.000 1507.330 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.630 0.000 1517.910 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.210 0.000 1528.490 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 0.000 1539.530 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.830 0.000 1550.110 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.870 0.000 1561.150 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.030 0.000 1582.310 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.070 0.000 1593.350 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 0.000 1603.930 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.230 0.000 1614.510 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.270 0.000 1625.550 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 0.000 1636.130 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.890 0.000 1647.170 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.470 0.000 1657.750 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 0.000 1668.330 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.090 0.000 1679.370 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.670 0.000 1689.950 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 0.000 1700.530 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.290 0.000 1711.570 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.870 0.000 1722.150 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.910 0.000 1733.190 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.490 0.000 1743.770 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.070 0.000 1754.350 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 0.000 625.510 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 0.000 722.110 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 0.000 743.730 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 0.000 840.330 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 0.000 850.910 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 0.000 883.570 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 0.000 894.150 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.450 0.000 904.730 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 0.000 915.770 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 0.000 926.350 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.690 0.000 947.970 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.270 0.000 958.550 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 0.000 980.170 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 0.000 990.750 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.090 0.000 1012.370 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 0.000 1023.410 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 0.000 1044.570 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.330 0.000 1055.610 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 0.000 1076.770 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 0.000 1087.810 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 0.000 1109.430 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.730 0.000 1120.010 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 0.000 1141.630 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.550 0.000 1173.830 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.130 0.000 1184.410 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.750 0.000 1206.030 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.330 0.000 1216.610 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 0.000 1227.650 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.950 0.000 1238.230 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990 0.000 1249.270 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.570 0.000 1259.850 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1270.150 0.000 1270.430 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.190 0.000 1281.470 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.770 0.000 1292.050 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.350 0.000 1302.630 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.390 0.000 1313.670 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.970 0.000 1324.250 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.010 0.000 1335.290 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.590 0.000 1345.870 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.170 0.000 1356.450 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.210 0.000 1367.490 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.790 0.000 1378.070 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.370 0.000 1388.650 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.410 0.000 1399.690 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.990 0.000 1410.270 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 0.000 1421.310 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.610 0.000 1431.890 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.190 0.000 1442.470 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.230 0.000 1453.510 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END la_oenb[9]
  PIN tag_array_ext_ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.160 4.000 1638.760 ;
    END
  END tag_array_ext_ram_addr1[0]
  PIN tag_array_ext_ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1642.240 4.000 1642.840 ;
    END
  END tag_array_ext_ram_addr1[1]
  PIN tag_array_ext_ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1645.640 4.000 1646.240 ;
    END
  END tag_array_ext_ram_addr1[2]
  PIN tag_array_ext_ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1649.040 4.000 1649.640 ;
    END
  END tag_array_ext_ram_addr1[3]
  PIN tag_array_ext_ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1652.440 4.000 1653.040 ;
    END
  END tag_array_ext_ram_addr1[4]
  PIN tag_array_ext_ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1655.840 4.000 1656.440 ;
    END
  END tag_array_ext_ram_addr1[5]
  PIN tag_array_ext_ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END tag_array_ext_ram_addr1[6]
  PIN tag_array_ext_ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1663.320 4.000 1663.920 ;
    END
  END tag_array_ext_ram_addr1[7]
  PIN tag_array_ext_ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END tag_array_ext_ram_addr[0]
  PIN tag_array_ext_ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1363.440 4.000 1364.040 ;
    END
  END tag_array_ext_ram_addr[1]
  PIN tag_array_ext_ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1367.520 4.000 1368.120 ;
    END
  END tag_array_ext_ram_addr[2]
  PIN tag_array_ext_ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.920 4.000 1371.520 ;
    END
  END tag_array_ext_ram_addr[3]
  PIN tag_array_ext_ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1374.320 4.000 1374.920 ;
    END
  END tag_array_ext_ram_addr[4]
  PIN tag_array_ext_ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.720 4.000 1378.320 ;
    END
  END tag_array_ext_ram_addr[5]
  PIN tag_array_ext_ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1381.120 4.000 1381.720 ;
    END
  END tag_array_ext_ram_addr[6]
  PIN tag_array_ext_ram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1385.200 4.000 1385.800 ;
    END
  END tag_array_ext_ram_addr[7]
  PIN tag_array_ext_ram_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1388.600 4.000 1389.200 ;
    END
  END tag_array_ext_ram_clk
  PIN tag_array_ext_ram_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1624.560 4.000 1625.160 ;
    END
  END tag_array_ext_ram_csb
  PIN tag_array_ext_ram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1631.360 4.000 1631.960 ;
    END
  END tag_array_ext_ram_csb1[0]
  PIN tag_array_ext_ram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1634.760 4.000 1635.360 ;
    END
  END tag_array_ext_ram_csb1[1]
  PIN tag_array_ext_ram_rdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END tag_array_ext_ram_rdata0[0]
  PIN tag_array_ext_ram_rdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1282.520 4.000 1283.120 ;
    END
  END tag_array_ext_ram_rdata0[10]
  PIN tag_array_ext_ram_rdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1286.600 4.000 1287.200 ;
    END
  END tag_array_ext_ram_rdata0[11]
  PIN tag_array_ext_ram_rdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1290.000 4.000 1290.600 ;
    END
  END tag_array_ext_ram_rdata0[12]
  PIN tag_array_ext_ram_rdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END tag_array_ext_ram_rdata0[13]
  PIN tag_array_ext_ram_rdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1296.800 4.000 1297.400 ;
    END
  END tag_array_ext_ram_rdata0[14]
  PIN tag_array_ext_ram_rdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.200 4.000 1300.800 ;
    END
  END tag_array_ext_ram_rdata0[15]
  PIN tag_array_ext_ram_rdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1303.600 4.000 1304.200 ;
    END
  END tag_array_ext_ram_rdata0[16]
  PIN tag_array_ext_ram_rdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1307.680 4.000 1308.280 ;
    END
  END tag_array_ext_ram_rdata0[17]
  PIN tag_array_ext_ram_rdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1311.080 4.000 1311.680 ;
    END
  END tag_array_ext_ram_rdata0[18]
  PIN tag_array_ext_ram_rdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1314.480 4.000 1315.080 ;
    END
  END tag_array_ext_ram_rdata0[19]
  PIN tag_array_ext_ram_rdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.240 4.000 1251.840 ;
    END
  END tag_array_ext_ram_rdata0[1]
  PIN tag_array_ext_ram_rdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1317.880 4.000 1318.480 ;
    END
  END tag_array_ext_ram_rdata0[20]
  PIN tag_array_ext_ram_rdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1321.280 4.000 1321.880 ;
    END
  END tag_array_ext_ram_rdata0[21]
  PIN tag_array_ext_ram_rdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1325.360 4.000 1325.960 ;
    END
  END tag_array_ext_ram_rdata0[22]
  PIN tag_array_ext_ram_rdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1328.760 4.000 1329.360 ;
    END
  END tag_array_ext_ram_rdata0[23]
  PIN tag_array_ext_ram_rdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.160 4.000 1332.760 ;
    END
  END tag_array_ext_ram_rdata0[24]
  PIN tag_array_ext_ram_rdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1335.560 4.000 1336.160 ;
    END
  END tag_array_ext_ram_rdata0[25]
  PIN tag_array_ext_ram_rdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1338.960 4.000 1339.560 ;
    END
  END tag_array_ext_ram_rdata0[26]
  PIN tag_array_ext_ram_rdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1342.360 4.000 1342.960 ;
    END
  END tag_array_ext_ram_rdata0[27]
  PIN tag_array_ext_ram_rdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1346.440 4.000 1347.040 ;
    END
  END tag_array_ext_ram_rdata0[28]
  PIN tag_array_ext_ram_rdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.840 4.000 1350.440 ;
    END
  END tag_array_ext_ram_rdata0[29]
  PIN tag_array_ext_ram_rdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END tag_array_ext_ram_rdata0[2]
  PIN tag_array_ext_ram_rdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END tag_array_ext_ram_rdata0[30]
  PIN tag_array_ext_ram_rdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1356.640 4.000 1357.240 ;
    END
  END tag_array_ext_ram_rdata0[31]
  PIN tag_array_ext_ram_rdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END tag_array_ext_ram_rdata0[3]
  PIN tag_array_ext_ram_rdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END tag_array_ext_ram_rdata0[4]
  PIN tag_array_ext_ram_rdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END tag_array_ext_ram_rdata0[5]
  PIN tag_array_ext_ram_rdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.920 4.000 1269.520 ;
    END
  END tag_array_ext_ram_rdata0[6]
  PIN tag_array_ext_ram_rdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1272.320 4.000 1272.920 ;
    END
  END tag_array_ext_ram_rdata0[7]
  PIN tag_array_ext_ram_rdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.720 4.000 1276.320 ;
    END
  END tag_array_ext_ram_rdata0[8]
  PIN tag_array_ext_ram_rdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.120 4.000 1279.720 ;
    END
  END tag_array_ext_ram_rdata0[9]
  PIN tag_array_ext_ram_rdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.720 4.000 1667.320 ;
    END
  END tag_array_ext_ram_rdata1[0]
  PIN tag_array_ext_ram_rdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1702.080 4.000 1702.680 ;
    END
  END tag_array_ext_ram_rdata1[10]
  PIN tag_array_ext_ram_rdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1705.480 4.000 1706.080 ;
    END
  END tag_array_ext_ram_rdata1[11]
  PIN tag_array_ext_ram_rdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1708.880 4.000 1709.480 ;
    END
  END tag_array_ext_ram_rdata1[12]
  PIN tag_array_ext_ram_rdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1712.280 4.000 1712.880 ;
    END
  END tag_array_ext_ram_rdata1[13]
  PIN tag_array_ext_ram_rdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.680 4.000 1716.280 ;
    END
  END tag_array_ext_ram_rdata1[14]
  PIN tag_array_ext_ram_rdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1719.080 4.000 1719.680 ;
    END
  END tag_array_ext_ram_rdata1[15]
  PIN tag_array_ext_ram_rdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.160 4.000 1723.760 ;
    END
  END tag_array_ext_ram_rdata1[16]
  PIN tag_array_ext_ram_rdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1726.560 4.000 1727.160 ;
    END
  END tag_array_ext_ram_rdata1[17]
  PIN tag_array_ext_ram_rdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1729.960 4.000 1730.560 ;
    END
  END tag_array_ext_ram_rdata1[18]
  PIN tag_array_ext_ram_rdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1733.360 4.000 1733.960 ;
    END
  END tag_array_ext_ram_rdata1[19]
  PIN tag_array_ext_ram_rdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1670.120 4.000 1670.720 ;
    END
  END tag_array_ext_ram_rdata1[1]
  PIN tag_array_ext_ram_rdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1736.760 4.000 1737.360 ;
    END
  END tag_array_ext_ram_rdata1[20]
  PIN tag_array_ext_ram_rdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1740.840 4.000 1741.440 ;
    END
  END tag_array_ext_ram_rdata1[21]
  PIN tag_array_ext_ram_rdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1744.240 4.000 1744.840 ;
    END
  END tag_array_ext_ram_rdata1[22]
  PIN tag_array_ext_ram_rdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END tag_array_ext_ram_rdata1[23]
  PIN tag_array_ext_ram_rdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.040 4.000 1751.640 ;
    END
  END tag_array_ext_ram_rdata1[24]
  PIN tag_array_ext_ram_rdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1754.440 4.000 1755.040 ;
    END
  END tag_array_ext_ram_rdata1[25]
  PIN tag_array_ext_ram_rdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.840 4.000 1758.440 ;
    END
  END tag_array_ext_ram_rdata1[26]
  PIN tag_array_ext_ram_rdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1761.920 4.000 1762.520 ;
    END
  END tag_array_ext_ram_rdata1[27]
  PIN tag_array_ext_ram_rdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1765.320 4.000 1765.920 ;
    END
  END tag_array_ext_ram_rdata1[28]
  PIN tag_array_ext_ram_rdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.720 4.000 1769.320 ;
    END
  END tag_array_ext_ram_rdata1[29]
  PIN tag_array_ext_ram_rdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1673.520 4.000 1674.120 ;
    END
  END tag_array_ext_ram_rdata1[2]
  PIN tag_array_ext_ram_rdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1772.120 4.000 1772.720 ;
    END
  END tag_array_ext_ram_rdata1[30]
  PIN tag_array_ext_ram_rdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1775.520 4.000 1776.120 ;
    END
  END tag_array_ext_ram_rdata1[31]
  PIN tag_array_ext_ram_rdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1676.920 4.000 1677.520 ;
    END
  END tag_array_ext_ram_rdata1[3]
  PIN tag_array_ext_ram_rdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1681.000 4.000 1681.600 ;
    END
  END tag_array_ext_ram_rdata1[4]
  PIN tag_array_ext_ram_rdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1684.400 4.000 1685.000 ;
    END
  END tag_array_ext_ram_rdata1[5]
  PIN tag_array_ext_ram_rdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1687.800 4.000 1688.400 ;
    END
  END tag_array_ext_ram_rdata1[6]
  PIN tag_array_ext_ram_rdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1691.200 4.000 1691.800 ;
    END
  END tag_array_ext_ram_rdata1[7]
  PIN tag_array_ext_ram_rdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1694.600 4.000 1695.200 ;
    END
  END tag_array_ext_ram_rdata1[8]
  PIN tag_array_ext_ram_rdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1698.000 4.000 1698.600 ;
    END
  END tag_array_ext_ram_rdata1[9]
  PIN tag_array_ext_ram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.000 4.000 1392.600 ;
    END
  END tag_array_ext_ram_wdata[0]
  PIN tag_array_ext_ram_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1427.360 4.000 1427.960 ;
    END
  END tag_array_ext_ram_wdata[10]
  PIN tag_array_ext_ram_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1430.760 4.000 1431.360 ;
    END
  END tag_array_ext_ram_wdata[11]
  PIN tag_array_ext_ram_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.160 4.000 1434.760 ;
    END
  END tag_array_ext_ram_wdata[12]
  PIN tag_array_ext_ram_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1437.560 4.000 1438.160 ;
    END
  END tag_array_ext_ram_wdata[13]
  PIN tag_array_ext_ram_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1440.960 4.000 1441.560 ;
    END
  END tag_array_ext_ram_wdata[14]
  PIN tag_array_ext_ram_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.040 4.000 1445.640 ;
    END
  END tag_array_ext_ram_wdata[15]
  PIN tag_array_ext_ram_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 4.000 1449.040 ;
    END
  END tag_array_ext_ram_wdata[16]
  PIN tag_array_ext_ram_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.840 4.000 1452.440 ;
    END
  END tag_array_ext_ram_wdata[17]
  PIN tag_array_ext_ram_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END tag_array_ext_ram_wdata[18]
  PIN tag_array_ext_ram_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END tag_array_ext_ram_wdata[19]
  PIN tag_array_ext_ram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1395.400 4.000 1396.000 ;
    END
  END tag_array_ext_ram_wdata[1]
  PIN tag_array_ext_ram_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END tag_array_ext_ram_wdata[20]
  PIN tag_array_ext_ram_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1466.120 4.000 1466.720 ;
    END
  END tag_array_ext_ram_wdata[21]
  PIN tag_array_ext_ram_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1469.520 4.000 1470.120 ;
    END
  END tag_array_ext_ram_wdata[22]
  PIN tag_array_ext_ram_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.920 4.000 1473.520 ;
    END
  END tag_array_ext_ram_wdata[23]
  PIN tag_array_ext_ram_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1476.320 4.000 1476.920 ;
    END
  END tag_array_ext_ram_wdata[24]
  PIN tag_array_ext_ram_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.720 4.000 1480.320 ;
    END
  END tag_array_ext_ram_wdata[25]
  PIN tag_array_ext_ram_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1483.800 4.000 1484.400 ;
    END
  END tag_array_ext_ram_wdata[26]
  PIN tag_array_ext_ram_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1487.200 4.000 1487.800 ;
    END
  END tag_array_ext_ram_wdata[27]
  PIN tag_array_ext_ram_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1490.600 4.000 1491.200 ;
    END
  END tag_array_ext_ram_wdata[28]
  PIN tag_array_ext_ram_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1494.000 4.000 1494.600 ;
    END
  END tag_array_ext_ram_wdata[29]
  PIN tag_array_ext_ram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1398.800 4.000 1399.400 ;
    END
  END tag_array_ext_ram_wdata[2]
  PIN tag_array_ext_ram_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1497.400 4.000 1498.000 ;
    END
  END tag_array_ext_ram_wdata[30]
  PIN tag_array_ext_ram_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1500.800 4.000 1501.400 ;
    END
  END tag_array_ext_ram_wdata[31]
  PIN tag_array_ext_ram_wdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1504.880 4.000 1505.480 ;
    END
  END tag_array_ext_ram_wdata[32]
  PIN tag_array_ext_ram_wdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1508.280 4.000 1508.880 ;
    END
  END tag_array_ext_ram_wdata[33]
  PIN tag_array_ext_ram_wdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1511.680 4.000 1512.280 ;
    END
  END tag_array_ext_ram_wdata[34]
  PIN tag_array_ext_ram_wdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1515.080 4.000 1515.680 ;
    END
  END tag_array_ext_ram_wdata[35]
  PIN tag_array_ext_ram_wdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1518.480 4.000 1519.080 ;
    END
  END tag_array_ext_ram_wdata[36]
  PIN tag_array_ext_ram_wdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1521.880 4.000 1522.480 ;
    END
  END tag_array_ext_ram_wdata[37]
  PIN tag_array_ext_ram_wdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1525.960 4.000 1526.560 ;
    END
  END tag_array_ext_ram_wdata[38]
  PIN tag_array_ext_ram_wdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1529.360 4.000 1529.960 ;
    END
  END tag_array_ext_ram_wdata[39]
  PIN tag_array_ext_ram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1402.200 4.000 1402.800 ;
    END
  END tag_array_ext_ram_wdata[3]
  PIN tag_array_ext_ram_wdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1532.760 4.000 1533.360 ;
    END
  END tag_array_ext_ram_wdata[40]
  PIN tag_array_ext_ram_wdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.160 4.000 1536.760 ;
    END
  END tag_array_ext_ram_wdata[41]
  PIN tag_array_ext_ram_wdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1539.560 4.000 1540.160 ;
    END
  END tag_array_ext_ram_wdata[42]
  PIN tag_array_ext_ram_wdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END tag_array_ext_ram_wdata[43]
  PIN tag_array_ext_ram_wdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.040 4.000 1547.640 ;
    END
  END tag_array_ext_ram_wdata[44]
  PIN tag_array_ext_ram_wdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END tag_array_ext_ram_wdata[45]
  PIN tag_array_ext_ram_wdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.840 4.000 1554.440 ;
    END
  END tag_array_ext_ram_wdata[46]
  PIN tag_array_ext_ram_wdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1557.240 4.000 1557.840 ;
    END
  END tag_array_ext_ram_wdata[47]
  PIN tag_array_ext_ram_wdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1560.640 4.000 1561.240 ;
    END
  END tag_array_ext_ram_wdata[48]
  PIN tag_array_ext_ram_wdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.720 4.000 1565.320 ;
    END
  END tag_array_ext_ram_wdata[49]
  PIN tag_array_ext_ram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1406.280 4.000 1406.880 ;
    END
  END tag_array_ext_ram_wdata[4]
  PIN tag_array_ext_ram_wdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1568.120 4.000 1568.720 ;
    END
  END tag_array_ext_ram_wdata[50]
  PIN tag_array_ext_ram_wdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1571.520 4.000 1572.120 ;
    END
  END tag_array_ext_ram_wdata[51]
  PIN tag_array_ext_ram_wdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.920 4.000 1575.520 ;
    END
  END tag_array_ext_ram_wdata[52]
  PIN tag_array_ext_ram_wdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1578.320 4.000 1578.920 ;
    END
  END tag_array_ext_ram_wdata[53]
  PIN tag_array_ext_ram_wdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1582.400 4.000 1583.000 ;
    END
  END tag_array_ext_ram_wdata[54]
  PIN tag_array_ext_ram_wdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1585.800 4.000 1586.400 ;
    END
  END tag_array_ext_ram_wdata[55]
  PIN tag_array_ext_ram_wdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1589.200 4.000 1589.800 ;
    END
  END tag_array_ext_ram_wdata[56]
  PIN tag_array_ext_ram_wdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1592.600 4.000 1593.200 ;
    END
  END tag_array_ext_ram_wdata[57]
  PIN tag_array_ext_ram_wdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1596.000 4.000 1596.600 ;
    END
  END tag_array_ext_ram_wdata[58]
  PIN tag_array_ext_ram_wdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1599.400 4.000 1600.000 ;
    END
  END tag_array_ext_ram_wdata[59]
  PIN tag_array_ext_ram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.680 4.000 1410.280 ;
    END
  END tag_array_ext_ram_wdata[5]
  PIN tag_array_ext_ram_wdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1603.480 4.000 1604.080 ;
    END
  END tag_array_ext_ram_wdata[60]
  PIN tag_array_ext_ram_wdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1606.880 4.000 1607.480 ;
    END
  END tag_array_ext_ram_wdata[61]
  PIN tag_array_ext_ram_wdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1610.280 4.000 1610.880 ;
    END
  END tag_array_ext_ram_wdata[62]
  PIN tag_array_ext_ram_wdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1613.680 4.000 1614.280 ;
    END
  END tag_array_ext_ram_wdata[63]
  PIN tag_array_ext_ram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1413.080 4.000 1413.680 ;
    END
  END tag_array_ext_ram_wdata[6]
  PIN tag_array_ext_ram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1416.480 4.000 1417.080 ;
    END
  END tag_array_ext_ram_wdata[7]
  PIN tag_array_ext_ram_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1419.880 4.000 1420.480 ;
    END
  END tag_array_ext_ram_wdata[8]
  PIN tag_array_ext_ram_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1423.960 4.000 1424.560 ;
    END
  END tag_array_ext_ram_wdata[9]
  PIN tag_array_ext_ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1627.960 4.000 1628.560 ;
    END
  END tag_array_ext_ram_web
  PIN tag_array_ext_ram_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1617.080 4.000 1617.680 ;
    END
  END tag_array_ext_ram_wmask[0]
  PIN tag_array_ext_ram_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1620.480 4.000 1621.080 ;
    END
  END tag_array_ext_ram_wmask[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1765.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1765.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1765.520 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1761.800 1765.365 ;
      LAYER met1 ;
        RECT 0.990 0.040 1767.250 1773.740 ;
      LAYER met2 ;
        RECT 1.020 1773.835 7.170 1774.530 ;
        RECT 8.010 1773.835 22.350 1774.530 ;
        RECT 23.190 1773.835 37.990 1774.530 ;
        RECT 38.830 1773.835 53.630 1774.530 ;
        RECT 54.470 1773.835 68.810 1774.530 ;
        RECT 69.650 1773.835 84.450 1774.530 ;
        RECT 85.290 1773.835 100.090 1774.530 ;
        RECT 100.930 1773.835 115.270 1774.530 ;
        RECT 116.110 1773.835 130.910 1774.530 ;
        RECT 131.750 1773.835 146.550 1774.530 ;
        RECT 147.390 1773.835 162.190 1774.530 ;
        RECT 163.030 1773.835 177.370 1774.530 ;
        RECT 178.210 1773.835 193.010 1774.530 ;
        RECT 193.850 1773.835 208.650 1774.530 ;
        RECT 209.490 1773.835 223.830 1774.530 ;
        RECT 224.670 1773.835 239.470 1774.530 ;
        RECT 240.310 1773.835 255.110 1774.530 ;
        RECT 255.950 1773.835 270.290 1774.530 ;
        RECT 271.130 1773.835 285.930 1774.530 ;
        RECT 286.770 1773.835 301.570 1774.530 ;
        RECT 302.410 1773.835 317.210 1774.530 ;
        RECT 318.050 1773.835 332.390 1774.530 ;
        RECT 333.230 1773.835 348.030 1774.530 ;
        RECT 348.870 1773.835 363.670 1774.530 ;
        RECT 364.510 1773.835 378.850 1774.530 ;
        RECT 379.690 1773.835 394.490 1774.530 ;
        RECT 395.330 1773.835 410.130 1774.530 ;
        RECT 410.970 1773.835 425.310 1774.530 ;
        RECT 426.150 1773.835 440.950 1774.530 ;
        RECT 441.790 1773.835 456.590 1774.530 ;
        RECT 457.430 1773.835 472.230 1774.530 ;
        RECT 473.070 1773.835 487.410 1774.530 ;
        RECT 488.250 1773.835 503.050 1774.530 ;
        RECT 503.890 1773.835 518.690 1774.530 ;
        RECT 519.530 1773.835 533.870 1774.530 ;
        RECT 534.710 1773.835 549.510 1774.530 ;
        RECT 550.350 1773.835 565.150 1774.530 ;
        RECT 565.990 1773.835 580.330 1774.530 ;
        RECT 581.170 1773.835 595.970 1774.530 ;
        RECT 596.810 1773.835 611.610 1774.530 ;
        RECT 612.450 1773.835 627.250 1774.530 ;
        RECT 628.090 1773.835 642.430 1774.530 ;
        RECT 643.270 1773.835 658.070 1774.530 ;
        RECT 658.910 1773.835 673.710 1774.530 ;
        RECT 674.550 1773.835 688.890 1774.530 ;
        RECT 689.730 1773.835 704.530 1774.530 ;
        RECT 705.370 1773.835 720.170 1774.530 ;
        RECT 721.010 1773.835 735.350 1774.530 ;
        RECT 736.190 1773.835 750.990 1774.530 ;
        RECT 751.830 1773.835 766.630 1774.530 ;
        RECT 767.470 1773.835 782.270 1774.530 ;
        RECT 783.110 1773.835 797.450 1774.530 ;
        RECT 798.290 1773.835 813.090 1774.530 ;
        RECT 813.930 1773.835 828.730 1774.530 ;
        RECT 829.570 1773.835 843.910 1774.530 ;
        RECT 844.750 1773.835 859.550 1774.530 ;
        RECT 860.390 1773.835 875.190 1774.530 ;
        RECT 876.030 1773.835 890.830 1774.530 ;
        RECT 891.670 1773.835 906.010 1774.530 ;
        RECT 906.850 1773.835 921.650 1774.530 ;
        RECT 922.490 1773.835 937.290 1774.530 ;
        RECT 938.130 1773.835 952.470 1774.530 ;
        RECT 953.310 1773.835 968.110 1774.530 ;
        RECT 968.950 1773.835 983.750 1774.530 ;
        RECT 984.590 1773.835 998.930 1774.530 ;
        RECT 999.770 1773.835 1014.570 1774.530 ;
        RECT 1015.410 1773.835 1030.210 1774.530 ;
        RECT 1031.050 1773.835 1045.850 1774.530 ;
        RECT 1046.690 1773.835 1061.030 1774.530 ;
        RECT 1061.870 1773.835 1076.670 1774.530 ;
        RECT 1077.510 1773.835 1092.310 1774.530 ;
        RECT 1093.150 1773.835 1107.490 1774.530 ;
        RECT 1108.330 1773.835 1123.130 1774.530 ;
        RECT 1123.970 1773.835 1138.770 1774.530 ;
        RECT 1139.610 1773.835 1153.950 1774.530 ;
        RECT 1154.790 1773.835 1169.590 1774.530 ;
        RECT 1170.430 1773.835 1185.230 1774.530 ;
        RECT 1186.070 1773.835 1200.870 1774.530 ;
        RECT 1201.710 1773.835 1216.050 1774.530 ;
        RECT 1216.890 1773.835 1231.690 1774.530 ;
        RECT 1232.530 1773.835 1247.330 1774.530 ;
        RECT 1248.170 1773.835 1262.510 1774.530 ;
        RECT 1263.350 1773.835 1278.150 1774.530 ;
        RECT 1278.990 1773.835 1293.790 1774.530 ;
        RECT 1294.630 1773.835 1308.970 1774.530 ;
        RECT 1309.810 1773.835 1324.610 1774.530 ;
        RECT 1325.450 1773.835 1340.250 1774.530 ;
        RECT 1341.090 1773.835 1355.890 1774.530 ;
        RECT 1356.730 1773.835 1371.070 1774.530 ;
        RECT 1371.910 1773.835 1386.710 1774.530 ;
        RECT 1387.550 1773.835 1402.350 1774.530 ;
        RECT 1403.190 1773.835 1417.530 1774.530 ;
        RECT 1418.370 1773.835 1433.170 1774.530 ;
        RECT 1434.010 1773.835 1448.810 1774.530 ;
        RECT 1449.650 1773.835 1463.990 1774.530 ;
        RECT 1464.830 1773.835 1479.630 1774.530 ;
        RECT 1480.470 1773.835 1495.270 1774.530 ;
        RECT 1496.110 1773.835 1510.910 1774.530 ;
        RECT 1511.750 1773.835 1526.090 1774.530 ;
        RECT 1526.930 1773.835 1541.730 1774.530 ;
        RECT 1542.570 1773.835 1557.370 1774.530 ;
        RECT 1558.210 1773.835 1572.550 1774.530 ;
        RECT 1573.390 1773.835 1588.190 1774.530 ;
        RECT 1589.030 1773.835 1603.830 1774.530 ;
        RECT 1604.670 1773.835 1619.010 1774.530 ;
        RECT 1619.850 1773.835 1634.650 1774.530 ;
        RECT 1635.490 1773.835 1650.290 1774.530 ;
        RECT 1651.130 1773.835 1665.930 1774.530 ;
        RECT 1666.770 1773.835 1681.110 1774.530 ;
        RECT 1681.950 1773.835 1696.750 1774.530 ;
        RECT 1697.590 1773.835 1712.390 1774.530 ;
        RECT 1713.230 1773.835 1727.570 1774.530 ;
        RECT 1728.410 1773.835 1743.210 1774.530 ;
        RECT 1744.050 1773.835 1758.850 1774.530 ;
        RECT 1759.690 1773.835 1767.230 1774.530 ;
        RECT 1.020 4.280 1767.230 1773.835 ;
        RECT 1.020 0.010 1.190 4.280 ;
        RECT 2.030 0.010 4.410 4.280 ;
        RECT 5.250 0.010 8.090 4.280 ;
        RECT 8.930 0.010 11.770 4.280 ;
        RECT 12.610 0.010 15.450 4.280 ;
        RECT 16.290 0.010 18.670 4.280 ;
        RECT 19.510 0.010 22.350 4.280 ;
        RECT 23.190 0.010 26.030 4.280 ;
        RECT 26.870 0.010 29.710 4.280 ;
        RECT 30.550 0.010 33.390 4.280 ;
        RECT 34.230 0.010 36.610 4.280 ;
        RECT 37.450 0.010 40.290 4.280 ;
        RECT 41.130 0.010 43.970 4.280 ;
        RECT 44.810 0.010 47.650 4.280 ;
        RECT 48.490 0.010 51.330 4.280 ;
        RECT 52.170 0.010 54.550 4.280 ;
        RECT 55.390 0.010 58.230 4.280 ;
        RECT 59.070 0.010 61.910 4.280 ;
        RECT 62.750 0.010 65.590 4.280 ;
        RECT 66.430 0.010 69.270 4.280 ;
        RECT 70.110 0.010 72.490 4.280 ;
        RECT 73.330 0.010 76.170 4.280 ;
        RECT 77.010 0.010 79.850 4.280 ;
        RECT 80.690 0.010 83.530 4.280 ;
        RECT 84.370 0.010 87.210 4.280 ;
        RECT 88.050 0.010 90.430 4.280 ;
        RECT 91.270 0.010 94.110 4.280 ;
        RECT 94.950 0.010 97.790 4.280 ;
        RECT 98.630 0.010 101.470 4.280 ;
        RECT 102.310 0.010 105.150 4.280 ;
        RECT 105.990 0.010 108.370 4.280 ;
        RECT 109.210 0.010 112.050 4.280 ;
        RECT 112.890 0.010 115.730 4.280 ;
        RECT 116.570 0.010 119.410 4.280 ;
        RECT 120.250 0.010 122.630 4.280 ;
        RECT 123.470 0.010 126.310 4.280 ;
        RECT 127.150 0.010 129.990 4.280 ;
        RECT 130.830 0.010 133.670 4.280 ;
        RECT 134.510 0.010 137.350 4.280 ;
        RECT 138.190 0.010 140.570 4.280 ;
        RECT 141.410 0.010 144.250 4.280 ;
        RECT 145.090 0.010 147.930 4.280 ;
        RECT 148.770 0.010 151.610 4.280 ;
        RECT 152.450 0.010 155.290 4.280 ;
        RECT 156.130 0.010 158.510 4.280 ;
        RECT 159.350 0.010 162.190 4.280 ;
        RECT 163.030 0.010 165.870 4.280 ;
        RECT 166.710 0.010 169.550 4.280 ;
        RECT 170.390 0.010 173.230 4.280 ;
        RECT 174.070 0.010 176.450 4.280 ;
        RECT 177.290 0.010 180.130 4.280 ;
        RECT 180.970 0.010 183.810 4.280 ;
        RECT 184.650 0.010 187.490 4.280 ;
        RECT 188.330 0.010 191.170 4.280 ;
        RECT 192.010 0.010 194.390 4.280 ;
        RECT 195.230 0.010 198.070 4.280 ;
        RECT 198.910 0.010 201.750 4.280 ;
        RECT 202.590 0.010 205.430 4.280 ;
        RECT 206.270 0.010 209.110 4.280 ;
        RECT 209.950 0.010 212.330 4.280 ;
        RECT 213.170 0.010 216.010 4.280 ;
        RECT 216.850 0.010 219.690 4.280 ;
        RECT 220.530 0.010 223.370 4.280 ;
        RECT 224.210 0.010 226.590 4.280 ;
        RECT 227.430 0.010 230.270 4.280 ;
        RECT 231.110 0.010 233.950 4.280 ;
        RECT 234.790 0.010 237.630 4.280 ;
        RECT 238.470 0.010 241.310 4.280 ;
        RECT 242.150 0.010 244.530 4.280 ;
        RECT 245.370 0.010 248.210 4.280 ;
        RECT 249.050 0.010 251.890 4.280 ;
        RECT 252.730 0.010 255.570 4.280 ;
        RECT 256.410 0.010 259.250 4.280 ;
        RECT 260.090 0.010 262.470 4.280 ;
        RECT 263.310 0.010 266.150 4.280 ;
        RECT 266.990 0.010 269.830 4.280 ;
        RECT 270.670 0.010 273.510 4.280 ;
        RECT 274.350 0.010 277.190 4.280 ;
        RECT 278.030 0.010 280.410 4.280 ;
        RECT 281.250 0.010 284.090 4.280 ;
        RECT 284.930 0.010 287.770 4.280 ;
        RECT 288.610 0.010 291.450 4.280 ;
        RECT 292.290 0.010 295.130 4.280 ;
        RECT 295.970 0.010 298.350 4.280 ;
        RECT 299.190 0.010 302.030 4.280 ;
        RECT 302.870 0.010 305.710 4.280 ;
        RECT 306.550 0.010 309.390 4.280 ;
        RECT 310.230 0.010 313.070 4.280 ;
        RECT 313.910 0.010 316.290 4.280 ;
        RECT 317.130 0.010 319.970 4.280 ;
        RECT 320.810 0.010 323.650 4.280 ;
        RECT 324.490 0.010 327.330 4.280 ;
        RECT 328.170 0.010 330.550 4.280 ;
        RECT 331.390 0.010 334.230 4.280 ;
        RECT 335.070 0.010 337.910 4.280 ;
        RECT 338.750 0.010 341.590 4.280 ;
        RECT 342.430 0.010 345.270 4.280 ;
        RECT 346.110 0.010 348.490 4.280 ;
        RECT 349.330 0.010 352.170 4.280 ;
        RECT 353.010 0.010 355.850 4.280 ;
        RECT 356.690 0.010 359.530 4.280 ;
        RECT 360.370 0.010 363.210 4.280 ;
        RECT 364.050 0.010 366.430 4.280 ;
        RECT 367.270 0.010 370.110 4.280 ;
        RECT 370.950 0.010 373.790 4.280 ;
        RECT 374.630 0.010 377.470 4.280 ;
        RECT 378.310 0.010 381.150 4.280 ;
        RECT 381.990 0.010 384.370 4.280 ;
        RECT 385.210 0.010 388.050 4.280 ;
        RECT 388.890 0.010 391.730 4.280 ;
        RECT 392.570 0.010 395.410 4.280 ;
        RECT 396.250 0.010 399.090 4.280 ;
        RECT 399.930 0.010 402.310 4.280 ;
        RECT 403.150 0.010 405.990 4.280 ;
        RECT 406.830 0.010 409.670 4.280 ;
        RECT 410.510 0.010 413.350 4.280 ;
        RECT 414.190 0.010 417.030 4.280 ;
        RECT 417.870 0.010 420.250 4.280 ;
        RECT 421.090 0.010 423.930 4.280 ;
        RECT 424.770 0.010 427.610 4.280 ;
        RECT 428.450 0.010 431.290 4.280 ;
        RECT 432.130 0.010 434.510 4.280 ;
        RECT 435.350 0.010 438.190 4.280 ;
        RECT 439.030 0.010 441.870 4.280 ;
        RECT 442.710 0.010 445.550 4.280 ;
        RECT 446.390 0.010 449.230 4.280 ;
        RECT 450.070 0.010 452.450 4.280 ;
        RECT 453.290 0.010 456.130 4.280 ;
        RECT 456.970 0.010 459.810 4.280 ;
        RECT 460.650 0.010 463.490 4.280 ;
        RECT 464.330 0.010 467.170 4.280 ;
        RECT 468.010 0.010 470.390 4.280 ;
        RECT 471.230 0.010 474.070 4.280 ;
        RECT 474.910 0.010 477.750 4.280 ;
        RECT 478.590 0.010 481.430 4.280 ;
        RECT 482.270 0.010 485.110 4.280 ;
        RECT 485.950 0.010 488.330 4.280 ;
        RECT 489.170 0.010 492.010 4.280 ;
        RECT 492.850 0.010 495.690 4.280 ;
        RECT 496.530 0.010 499.370 4.280 ;
        RECT 500.210 0.010 503.050 4.280 ;
        RECT 503.890 0.010 506.270 4.280 ;
        RECT 507.110 0.010 509.950 4.280 ;
        RECT 510.790 0.010 513.630 4.280 ;
        RECT 514.470 0.010 517.310 4.280 ;
        RECT 518.150 0.010 520.990 4.280 ;
        RECT 521.830 0.010 524.210 4.280 ;
        RECT 525.050 0.010 527.890 4.280 ;
        RECT 528.730 0.010 531.570 4.280 ;
        RECT 532.410 0.010 535.250 4.280 ;
        RECT 536.090 0.010 538.470 4.280 ;
        RECT 539.310 0.010 542.150 4.280 ;
        RECT 542.990 0.010 545.830 4.280 ;
        RECT 546.670 0.010 549.510 4.280 ;
        RECT 550.350 0.010 553.190 4.280 ;
        RECT 554.030 0.010 556.410 4.280 ;
        RECT 557.250 0.010 560.090 4.280 ;
        RECT 560.930 0.010 563.770 4.280 ;
        RECT 564.610 0.010 567.450 4.280 ;
        RECT 568.290 0.010 571.130 4.280 ;
        RECT 571.970 0.010 574.350 4.280 ;
        RECT 575.190 0.010 578.030 4.280 ;
        RECT 578.870 0.010 581.710 4.280 ;
        RECT 582.550 0.010 585.390 4.280 ;
        RECT 586.230 0.010 589.070 4.280 ;
        RECT 589.910 0.010 592.290 4.280 ;
        RECT 593.130 0.010 595.970 4.280 ;
        RECT 596.810 0.010 599.650 4.280 ;
        RECT 600.490 0.010 603.330 4.280 ;
        RECT 604.170 0.010 607.010 4.280 ;
        RECT 607.850 0.010 610.230 4.280 ;
        RECT 611.070 0.010 613.910 4.280 ;
        RECT 614.750 0.010 617.590 4.280 ;
        RECT 618.430 0.010 621.270 4.280 ;
        RECT 622.110 0.010 624.950 4.280 ;
        RECT 625.790 0.010 628.170 4.280 ;
        RECT 629.010 0.010 631.850 4.280 ;
        RECT 632.690 0.010 635.530 4.280 ;
        RECT 636.370 0.010 639.210 4.280 ;
        RECT 640.050 0.010 642.430 4.280 ;
        RECT 643.270 0.010 646.110 4.280 ;
        RECT 646.950 0.010 649.790 4.280 ;
        RECT 650.630 0.010 653.470 4.280 ;
        RECT 654.310 0.010 657.150 4.280 ;
        RECT 657.990 0.010 660.370 4.280 ;
        RECT 661.210 0.010 664.050 4.280 ;
        RECT 664.890 0.010 667.730 4.280 ;
        RECT 668.570 0.010 671.410 4.280 ;
        RECT 672.250 0.010 675.090 4.280 ;
        RECT 675.930 0.010 678.310 4.280 ;
        RECT 679.150 0.010 681.990 4.280 ;
        RECT 682.830 0.010 685.670 4.280 ;
        RECT 686.510 0.010 689.350 4.280 ;
        RECT 690.190 0.010 693.030 4.280 ;
        RECT 693.870 0.010 696.250 4.280 ;
        RECT 697.090 0.010 699.930 4.280 ;
        RECT 700.770 0.010 703.610 4.280 ;
        RECT 704.450 0.010 707.290 4.280 ;
        RECT 708.130 0.010 710.970 4.280 ;
        RECT 711.810 0.010 714.190 4.280 ;
        RECT 715.030 0.010 717.870 4.280 ;
        RECT 718.710 0.010 721.550 4.280 ;
        RECT 722.390 0.010 725.230 4.280 ;
        RECT 726.070 0.010 728.910 4.280 ;
        RECT 729.750 0.010 732.130 4.280 ;
        RECT 732.970 0.010 735.810 4.280 ;
        RECT 736.650 0.010 739.490 4.280 ;
        RECT 740.330 0.010 743.170 4.280 ;
        RECT 744.010 0.010 746.390 4.280 ;
        RECT 747.230 0.010 750.070 4.280 ;
        RECT 750.910 0.010 753.750 4.280 ;
        RECT 754.590 0.010 757.430 4.280 ;
        RECT 758.270 0.010 761.110 4.280 ;
        RECT 761.950 0.010 764.330 4.280 ;
        RECT 765.170 0.010 768.010 4.280 ;
        RECT 768.850 0.010 771.690 4.280 ;
        RECT 772.530 0.010 775.370 4.280 ;
        RECT 776.210 0.010 779.050 4.280 ;
        RECT 779.890 0.010 782.270 4.280 ;
        RECT 783.110 0.010 785.950 4.280 ;
        RECT 786.790 0.010 789.630 4.280 ;
        RECT 790.470 0.010 793.310 4.280 ;
        RECT 794.150 0.010 796.990 4.280 ;
        RECT 797.830 0.010 800.210 4.280 ;
        RECT 801.050 0.010 803.890 4.280 ;
        RECT 804.730 0.010 807.570 4.280 ;
        RECT 808.410 0.010 811.250 4.280 ;
        RECT 812.090 0.010 814.930 4.280 ;
        RECT 815.770 0.010 818.150 4.280 ;
        RECT 818.990 0.010 821.830 4.280 ;
        RECT 822.670 0.010 825.510 4.280 ;
        RECT 826.350 0.010 829.190 4.280 ;
        RECT 830.030 0.010 832.870 4.280 ;
        RECT 833.710 0.010 836.090 4.280 ;
        RECT 836.930 0.010 839.770 4.280 ;
        RECT 840.610 0.010 843.450 4.280 ;
        RECT 844.290 0.010 847.130 4.280 ;
        RECT 847.970 0.010 850.350 4.280 ;
        RECT 851.190 0.010 854.030 4.280 ;
        RECT 854.870 0.010 857.710 4.280 ;
        RECT 858.550 0.010 861.390 4.280 ;
        RECT 862.230 0.010 865.070 4.280 ;
        RECT 865.910 0.010 868.290 4.280 ;
        RECT 869.130 0.010 871.970 4.280 ;
        RECT 872.810 0.010 875.650 4.280 ;
        RECT 876.490 0.010 879.330 4.280 ;
        RECT 880.170 0.010 883.010 4.280 ;
        RECT 883.850 0.010 886.230 4.280 ;
        RECT 887.070 0.010 889.910 4.280 ;
        RECT 890.750 0.010 893.590 4.280 ;
        RECT 894.430 0.010 897.270 4.280 ;
        RECT 898.110 0.010 900.950 4.280 ;
        RECT 901.790 0.010 904.170 4.280 ;
        RECT 905.010 0.010 907.850 4.280 ;
        RECT 908.690 0.010 911.530 4.280 ;
        RECT 912.370 0.010 915.210 4.280 ;
        RECT 916.050 0.010 918.890 4.280 ;
        RECT 919.730 0.010 922.110 4.280 ;
        RECT 922.950 0.010 925.790 4.280 ;
        RECT 926.630 0.010 929.470 4.280 ;
        RECT 930.310 0.010 933.150 4.280 ;
        RECT 933.990 0.010 936.830 4.280 ;
        RECT 937.670 0.010 940.050 4.280 ;
        RECT 940.890 0.010 943.730 4.280 ;
        RECT 944.570 0.010 947.410 4.280 ;
        RECT 948.250 0.010 951.090 4.280 ;
        RECT 951.930 0.010 954.310 4.280 ;
        RECT 955.150 0.010 957.990 4.280 ;
        RECT 958.830 0.010 961.670 4.280 ;
        RECT 962.510 0.010 965.350 4.280 ;
        RECT 966.190 0.010 969.030 4.280 ;
        RECT 969.870 0.010 972.250 4.280 ;
        RECT 973.090 0.010 975.930 4.280 ;
        RECT 976.770 0.010 979.610 4.280 ;
        RECT 980.450 0.010 983.290 4.280 ;
        RECT 984.130 0.010 986.970 4.280 ;
        RECT 987.810 0.010 990.190 4.280 ;
        RECT 991.030 0.010 993.870 4.280 ;
        RECT 994.710 0.010 997.550 4.280 ;
        RECT 998.390 0.010 1001.230 4.280 ;
        RECT 1002.070 0.010 1004.910 4.280 ;
        RECT 1005.750 0.010 1008.130 4.280 ;
        RECT 1008.970 0.010 1011.810 4.280 ;
        RECT 1012.650 0.010 1015.490 4.280 ;
        RECT 1016.330 0.010 1019.170 4.280 ;
        RECT 1020.010 0.010 1022.850 4.280 ;
        RECT 1023.690 0.010 1026.070 4.280 ;
        RECT 1026.910 0.010 1029.750 4.280 ;
        RECT 1030.590 0.010 1033.430 4.280 ;
        RECT 1034.270 0.010 1037.110 4.280 ;
        RECT 1037.950 0.010 1040.790 4.280 ;
        RECT 1041.630 0.010 1044.010 4.280 ;
        RECT 1044.850 0.010 1047.690 4.280 ;
        RECT 1048.530 0.010 1051.370 4.280 ;
        RECT 1052.210 0.010 1055.050 4.280 ;
        RECT 1055.890 0.010 1058.270 4.280 ;
        RECT 1059.110 0.010 1061.950 4.280 ;
        RECT 1062.790 0.010 1065.630 4.280 ;
        RECT 1066.470 0.010 1069.310 4.280 ;
        RECT 1070.150 0.010 1072.990 4.280 ;
        RECT 1073.830 0.010 1076.210 4.280 ;
        RECT 1077.050 0.010 1079.890 4.280 ;
        RECT 1080.730 0.010 1083.570 4.280 ;
        RECT 1084.410 0.010 1087.250 4.280 ;
        RECT 1088.090 0.010 1090.930 4.280 ;
        RECT 1091.770 0.010 1094.150 4.280 ;
        RECT 1094.990 0.010 1097.830 4.280 ;
        RECT 1098.670 0.010 1101.510 4.280 ;
        RECT 1102.350 0.010 1105.190 4.280 ;
        RECT 1106.030 0.010 1108.870 4.280 ;
        RECT 1109.710 0.010 1112.090 4.280 ;
        RECT 1112.930 0.010 1115.770 4.280 ;
        RECT 1116.610 0.010 1119.450 4.280 ;
        RECT 1120.290 0.010 1123.130 4.280 ;
        RECT 1123.970 0.010 1126.810 4.280 ;
        RECT 1127.650 0.010 1130.030 4.280 ;
        RECT 1130.870 0.010 1133.710 4.280 ;
        RECT 1134.550 0.010 1137.390 4.280 ;
        RECT 1138.230 0.010 1141.070 4.280 ;
        RECT 1141.910 0.010 1144.750 4.280 ;
        RECT 1145.590 0.010 1147.970 4.280 ;
        RECT 1148.810 0.010 1151.650 4.280 ;
        RECT 1152.490 0.010 1155.330 4.280 ;
        RECT 1156.170 0.010 1159.010 4.280 ;
        RECT 1159.850 0.010 1162.230 4.280 ;
        RECT 1163.070 0.010 1165.910 4.280 ;
        RECT 1166.750 0.010 1169.590 4.280 ;
        RECT 1170.430 0.010 1173.270 4.280 ;
        RECT 1174.110 0.010 1176.950 4.280 ;
        RECT 1177.790 0.010 1180.170 4.280 ;
        RECT 1181.010 0.010 1183.850 4.280 ;
        RECT 1184.690 0.010 1187.530 4.280 ;
        RECT 1188.370 0.010 1191.210 4.280 ;
        RECT 1192.050 0.010 1194.890 4.280 ;
        RECT 1195.730 0.010 1198.110 4.280 ;
        RECT 1198.950 0.010 1201.790 4.280 ;
        RECT 1202.630 0.010 1205.470 4.280 ;
        RECT 1206.310 0.010 1209.150 4.280 ;
        RECT 1209.990 0.010 1212.830 4.280 ;
        RECT 1213.670 0.010 1216.050 4.280 ;
        RECT 1216.890 0.010 1219.730 4.280 ;
        RECT 1220.570 0.010 1223.410 4.280 ;
        RECT 1224.250 0.010 1227.090 4.280 ;
        RECT 1227.930 0.010 1230.770 4.280 ;
        RECT 1231.610 0.010 1233.990 4.280 ;
        RECT 1234.830 0.010 1237.670 4.280 ;
        RECT 1238.510 0.010 1241.350 4.280 ;
        RECT 1242.190 0.010 1245.030 4.280 ;
        RECT 1245.870 0.010 1248.710 4.280 ;
        RECT 1249.550 0.010 1251.930 4.280 ;
        RECT 1252.770 0.010 1255.610 4.280 ;
        RECT 1256.450 0.010 1259.290 4.280 ;
        RECT 1260.130 0.010 1262.970 4.280 ;
        RECT 1263.810 0.010 1266.190 4.280 ;
        RECT 1267.030 0.010 1269.870 4.280 ;
        RECT 1270.710 0.010 1273.550 4.280 ;
        RECT 1274.390 0.010 1277.230 4.280 ;
        RECT 1278.070 0.010 1280.910 4.280 ;
        RECT 1281.750 0.010 1284.130 4.280 ;
        RECT 1284.970 0.010 1287.810 4.280 ;
        RECT 1288.650 0.010 1291.490 4.280 ;
        RECT 1292.330 0.010 1295.170 4.280 ;
        RECT 1296.010 0.010 1298.850 4.280 ;
        RECT 1299.690 0.010 1302.070 4.280 ;
        RECT 1302.910 0.010 1305.750 4.280 ;
        RECT 1306.590 0.010 1309.430 4.280 ;
        RECT 1310.270 0.010 1313.110 4.280 ;
        RECT 1313.950 0.010 1316.790 4.280 ;
        RECT 1317.630 0.010 1320.010 4.280 ;
        RECT 1320.850 0.010 1323.690 4.280 ;
        RECT 1324.530 0.010 1327.370 4.280 ;
        RECT 1328.210 0.010 1331.050 4.280 ;
        RECT 1331.890 0.010 1334.730 4.280 ;
        RECT 1335.570 0.010 1337.950 4.280 ;
        RECT 1338.790 0.010 1341.630 4.280 ;
        RECT 1342.470 0.010 1345.310 4.280 ;
        RECT 1346.150 0.010 1348.990 4.280 ;
        RECT 1349.830 0.010 1352.670 4.280 ;
        RECT 1353.510 0.010 1355.890 4.280 ;
        RECT 1356.730 0.010 1359.570 4.280 ;
        RECT 1360.410 0.010 1363.250 4.280 ;
        RECT 1364.090 0.010 1366.930 4.280 ;
        RECT 1367.770 0.010 1370.150 4.280 ;
        RECT 1370.990 0.010 1373.830 4.280 ;
        RECT 1374.670 0.010 1377.510 4.280 ;
        RECT 1378.350 0.010 1381.190 4.280 ;
        RECT 1382.030 0.010 1384.870 4.280 ;
        RECT 1385.710 0.010 1388.090 4.280 ;
        RECT 1388.930 0.010 1391.770 4.280 ;
        RECT 1392.610 0.010 1395.450 4.280 ;
        RECT 1396.290 0.010 1399.130 4.280 ;
        RECT 1399.970 0.010 1402.810 4.280 ;
        RECT 1403.650 0.010 1406.030 4.280 ;
        RECT 1406.870 0.010 1409.710 4.280 ;
        RECT 1410.550 0.010 1413.390 4.280 ;
        RECT 1414.230 0.010 1417.070 4.280 ;
        RECT 1417.910 0.010 1420.750 4.280 ;
        RECT 1421.590 0.010 1423.970 4.280 ;
        RECT 1424.810 0.010 1427.650 4.280 ;
        RECT 1428.490 0.010 1431.330 4.280 ;
        RECT 1432.170 0.010 1435.010 4.280 ;
        RECT 1435.850 0.010 1438.690 4.280 ;
        RECT 1439.530 0.010 1441.910 4.280 ;
        RECT 1442.750 0.010 1445.590 4.280 ;
        RECT 1446.430 0.010 1449.270 4.280 ;
        RECT 1450.110 0.010 1452.950 4.280 ;
        RECT 1453.790 0.010 1456.630 4.280 ;
        RECT 1457.470 0.010 1459.850 4.280 ;
        RECT 1460.690 0.010 1463.530 4.280 ;
        RECT 1464.370 0.010 1467.210 4.280 ;
        RECT 1468.050 0.010 1470.890 4.280 ;
        RECT 1471.730 0.010 1474.110 4.280 ;
        RECT 1474.950 0.010 1477.790 4.280 ;
        RECT 1478.630 0.010 1481.470 4.280 ;
        RECT 1482.310 0.010 1485.150 4.280 ;
        RECT 1485.990 0.010 1488.830 4.280 ;
        RECT 1489.670 0.010 1492.050 4.280 ;
        RECT 1492.890 0.010 1495.730 4.280 ;
        RECT 1496.570 0.010 1499.410 4.280 ;
        RECT 1500.250 0.010 1503.090 4.280 ;
        RECT 1503.930 0.010 1506.770 4.280 ;
        RECT 1507.610 0.010 1509.990 4.280 ;
        RECT 1510.830 0.010 1513.670 4.280 ;
        RECT 1514.510 0.010 1517.350 4.280 ;
        RECT 1518.190 0.010 1521.030 4.280 ;
        RECT 1521.870 0.010 1524.710 4.280 ;
        RECT 1525.550 0.010 1527.930 4.280 ;
        RECT 1528.770 0.010 1531.610 4.280 ;
        RECT 1532.450 0.010 1535.290 4.280 ;
        RECT 1536.130 0.010 1538.970 4.280 ;
        RECT 1539.810 0.010 1542.650 4.280 ;
        RECT 1543.490 0.010 1545.870 4.280 ;
        RECT 1546.710 0.010 1549.550 4.280 ;
        RECT 1550.390 0.010 1553.230 4.280 ;
        RECT 1554.070 0.010 1556.910 4.280 ;
        RECT 1557.750 0.010 1560.590 4.280 ;
        RECT 1561.430 0.010 1563.810 4.280 ;
        RECT 1564.650 0.010 1567.490 4.280 ;
        RECT 1568.330 0.010 1571.170 4.280 ;
        RECT 1572.010 0.010 1574.850 4.280 ;
        RECT 1575.690 0.010 1578.070 4.280 ;
        RECT 1578.910 0.010 1581.750 4.280 ;
        RECT 1582.590 0.010 1585.430 4.280 ;
        RECT 1586.270 0.010 1589.110 4.280 ;
        RECT 1589.950 0.010 1592.790 4.280 ;
        RECT 1593.630 0.010 1596.010 4.280 ;
        RECT 1596.850 0.010 1599.690 4.280 ;
        RECT 1600.530 0.010 1603.370 4.280 ;
        RECT 1604.210 0.010 1607.050 4.280 ;
        RECT 1607.890 0.010 1610.730 4.280 ;
        RECT 1611.570 0.010 1613.950 4.280 ;
        RECT 1614.790 0.010 1617.630 4.280 ;
        RECT 1618.470 0.010 1621.310 4.280 ;
        RECT 1622.150 0.010 1624.990 4.280 ;
        RECT 1625.830 0.010 1628.670 4.280 ;
        RECT 1629.510 0.010 1631.890 4.280 ;
        RECT 1632.730 0.010 1635.570 4.280 ;
        RECT 1636.410 0.010 1639.250 4.280 ;
        RECT 1640.090 0.010 1642.930 4.280 ;
        RECT 1643.770 0.010 1646.610 4.280 ;
        RECT 1647.450 0.010 1649.830 4.280 ;
        RECT 1650.670 0.010 1653.510 4.280 ;
        RECT 1654.350 0.010 1657.190 4.280 ;
        RECT 1658.030 0.010 1660.870 4.280 ;
        RECT 1661.710 0.010 1664.550 4.280 ;
        RECT 1665.390 0.010 1667.770 4.280 ;
        RECT 1668.610 0.010 1671.450 4.280 ;
        RECT 1672.290 0.010 1675.130 4.280 ;
        RECT 1675.970 0.010 1678.810 4.280 ;
        RECT 1679.650 0.010 1682.030 4.280 ;
        RECT 1682.870 0.010 1685.710 4.280 ;
        RECT 1686.550 0.010 1689.390 4.280 ;
        RECT 1690.230 0.010 1693.070 4.280 ;
        RECT 1693.910 0.010 1696.750 4.280 ;
        RECT 1697.590 0.010 1699.970 4.280 ;
        RECT 1700.810 0.010 1703.650 4.280 ;
        RECT 1704.490 0.010 1707.330 4.280 ;
        RECT 1708.170 0.010 1711.010 4.280 ;
        RECT 1711.850 0.010 1714.690 4.280 ;
        RECT 1715.530 0.010 1717.910 4.280 ;
        RECT 1718.750 0.010 1721.590 4.280 ;
        RECT 1722.430 0.010 1725.270 4.280 ;
        RECT 1726.110 0.010 1728.950 4.280 ;
        RECT 1729.790 0.010 1732.630 4.280 ;
        RECT 1733.470 0.010 1735.850 4.280 ;
        RECT 1736.690 0.010 1739.530 4.280 ;
        RECT 1740.370 0.010 1743.210 4.280 ;
        RECT 1744.050 0.010 1746.890 4.280 ;
        RECT 1747.730 0.010 1750.570 4.280 ;
        RECT 1751.410 0.010 1753.790 4.280 ;
        RECT 1754.630 0.010 1757.470 4.280 ;
        RECT 1758.310 0.010 1761.150 4.280 ;
        RECT 1761.990 0.010 1764.830 4.280 ;
        RECT 1765.670 0.010 1767.230 4.280 ;
      LAYER met3 ;
        RECT 1.445 1773.120 1762.995 1773.265 ;
        RECT 4.400 1772.400 1762.995 1773.120 ;
        RECT 4.400 1771.720 1767.255 1772.400 ;
        RECT 1.445 1769.720 1767.255 1771.720 ;
        RECT 4.400 1768.320 1767.255 1769.720 ;
        RECT 1.445 1766.320 1767.255 1768.320 ;
        RECT 4.400 1764.960 1767.255 1766.320 ;
        RECT 4.400 1764.920 1762.995 1764.960 ;
        RECT 1.445 1763.560 1762.995 1764.920 ;
        RECT 1.445 1762.920 1767.255 1763.560 ;
        RECT 4.400 1761.520 1767.255 1762.920 ;
        RECT 1.445 1758.840 1767.255 1761.520 ;
        RECT 4.400 1757.440 1767.255 1758.840 ;
        RECT 1.445 1756.120 1767.255 1757.440 ;
        RECT 1.445 1755.440 1762.995 1756.120 ;
        RECT 4.400 1754.720 1762.995 1755.440 ;
        RECT 4.400 1754.040 1767.255 1754.720 ;
        RECT 1.445 1752.040 1767.255 1754.040 ;
        RECT 4.400 1750.640 1767.255 1752.040 ;
        RECT 1.445 1748.640 1767.255 1750.640 ;
        RECT 4.400 1747.280 1767.255 1748.640 ;
        RECT 4.400 1747.240 1762.995 1747.280 ;
        RECT 1.445 1745.880 1762.995 1747.240 ;
        RECT 1.445 1745.240 1767.255 1745.880 ;
        RECT 4.400 1743.840 1767.255 1745.240 ;
        RECT 1.445 1741.840 1767.255 1743.840 ;
        RECT 4.400 1740.440 1767.255 1741.840 ;
        RECT 1.445 1738.440 1767.255 1740.440 ;
        RECT 1.445 1737.760 1762.995 1738.440 ;
        RECT 4.400 1737.040 1762.995 1737.760 ;
        RECT 4.400 1736.360 1767.255 1737.040 ;
        RECT 1.445 1734.360 1767.255 1736.360 ;
        RECT 4.400 1732.960 1767.255 1734.360 ;
        RECT 1.445 1730.960 1767.255 1732.960 ;
        RECT 4.400 1729.600 1767.255 1730.960 ;
        RECT 4.400 1729.560 1762.995 1729.600 ;
        RECT 1.445 1728.200 1762.995 1729.560 ;
        RECT 1.445 1727.560 1767.255 1728.200 ;
        RECT 4.400 1726.160 1767.255 1727.560 ;
        RECT 1.445 1724.160 1767.255 1726.160 ;
        RECT 4.400 1722.760 1767.255 1724.160 ;
        RECT 1.445 1720.760 1767.255 1722.760 ;
        RECT 1.445 1720.080 1762.995 1720.760 ;
        RECT 4.400 1719.360 1762.995 1720.080 ;
        RECT 4.400 1718.680 1767.255 1719.360 ;
        RECT 1.445 1716.680 1767.255 1718.680 ;
        RECT 4.400 1715.280 1767.255 1716.680 ;
        RECT 1.445 1713.280 1767.255 1715.280 ;
        RECT 4.400 1711.920 1767.255 1713.280 ;
        RECT 4.400 1711.880 1762.995 1711.920 ;
        RECT 1.445 1710.520 1762.995 1711.880 ;
        RECT 1.445 1709.880 1767.255 1710.520 ;
        RECT 4.400 1708.480 1767.255 1709.880 ;
        RECT 1.445 1706.480 1767.255 1708.480 ;
        RECT 4.400 1705.080 1767.255 1706.480 ;
        RECT 1.445 1703.080 1767.255 1705.080 ;
        RECT 4.400 1701.680 1762.995 1703.080 ;
        RECT 1.445 1699.000 1767.255 1701.680 ;
        RECT 4.400 1697.600 1767.255 1699.000 ;
        RECT 1.445 1695.600 1767.255 1697.600 ;
        RECT 4.400 1694.240 1767.255 1695.600 ;
        RECT 4.400 1694.200 1762.995 1694.240 ;
        RECT 1.445 1692.840 1762.995 1694.200 ;
        RECT 1.445 1692.200 1767.255 1692.840 ;
        RECT 4.400 1690.800 1767.255 1692.200 ;
        RECT 1.445 1688.800 1767.255 1690.800 ;
        RECT 4.400 1687.400 1767.255 1688.800 ;
        RECT 1.445 1685.400 1767.255 1687.400 ;
        RECT 4.400 1684.000 1762.995 1685.400 ;
        RECT 1.445 1682.000 1767.255 1684.000 ;
        RECT 4.400 1680.600 1767.255 1682.000 ;
        RECT 1.445 1677.920 1767.255 1680.600 ;
        RECT 4.400 1676.560 1767.255 1677.920 ;
        RECT 4.400 1676.520 1762.995 1676.560 ;
        RECT 1.445 1675.160 1762.995 1676.520 ;
        RECT 1.445 1674.520 1767.255 1675.160 ;
        RECT 4.400 1673.120 1767.255 1674.520 ;
        RECT 1.445 1671.120 1767.255 1673.120 ;
        RECT 4.400 1669.720 1767.255 1671.120 ;
        RECT 1.445 1667.720 1767.255 1669.720 ;
        RECT 4.400 1666.320 1762.995 1667.720 ;
        RECT 1.445 1664.320 1767.255 1666.320 ;
        RECT 4.400 1662.920 1767.255 1664.320 ;
        RECT 1.445 1660.240 1767.255 1662.920 ;
        RECT 4.400 1658.840 1767.255 1660.240 ;
        RECT 1.445 1658.200 1767.255 1658.840 ;
        RECT 1.445 1656.840 1762.995 1658.200 ;
        RECT 4.400 1656.800 1762.995 1656.840 ;
        RECT 4.400 1655.440 1767.255 1656.800 ;
        RECT 1.445 1653.440 1767.255 1655.440 ;
        RECT 4.400 1652.040 1767.255 1653.440 ;
        RECT 1.445 1650.040 1767.255 1652.040 ;
        RECT 4.400 1649.360 1767.255 1650.040 ;
        RECT 4.400 1648.640 1762.995 1649.360 ;
        RECT 1.445 1647.960 1762.995 1648.640 ;
        RECT 1.445 1646.640 1767.255 1647.960 ;
        RECT 4.400 1645.240 1767.255 1646.640 ;
        RECT 1.445 1643.240 1767.255 1645.240 ;
        RECT 4.400 1641.840 1767.255 1643.240 ;
        RECT 1.445 1640.520 1767.255 1641.840 ;
        RECT 1.445 1639.160 1762.995 1640.520 ;
        RECT 4.400 1639.120 1762.995 1639.160 ;
        RECT 4.400 1637.760 1767.255 1639.120 ;
        RECT 1.445 1635.760 1767.255 1637.760 ;
        RECT 4.400 1634.360 1767.255 1635.760 ;
        RECT 1.445 1632.360 1767.255 1634.360 ;
        RECT 4.400 1631.680 1767.255 1632.360 ;
        RECT 4.400 1630.960 1762.995 1631.680 ;
        RECT 1.445 1630.280 1762.995 1630.960 ;
        RECT 1.445 1628.960 1767.255 1630.280 ;
        RECT 4.400 1627.560 1767.255 1628.960 ;
        RECT 1.445 1625.560 1767.255 1627.560 ;
        RECT 4.400 1624.160 1767.255 1625.560 ;
        RECT 1.445 1622.840 1767.255 1624.160 ;
        RECT 1.445 1621.480 1762.995 1622.840 ;
        RECT 4.400 1621.440 1762.995 1621.480 ;
        RECT 4.400 1620.080 1767.255 1621.440 ;
        RECT 1.445 1618.080 1767.255 1620.080 ;
        RECT 4.400 1616.680 1767.255 1618.080 ;
        RECT 1.445 1614.680 1767.255 1616.680 ;
        RECT 4.400 1614.000 1767.255 1614.680 ;
        RECT 4.400 1613.280 1762.995 1614.000 ;
        RECT 1.445 1612.600 1762.995 1613.280 ;
        RECT 1.445 1611.280 1767.255 1612.600 ;
        RECT 4.400 1609.880 1767.255 1611.280 ;
        RECT 1.445 1607.880 1767.255 1609.880 ;
        RECT 4.400 1606.480 1767.255 1607.880 ;
        RECT 1.445 1605.160 1767.255 1606.480 ;
        RECT 1.445 1604.480 1762.995 1605.160 ;
        RECT 4.400 1603.760 1762.995 1604.480 ;
        RECT 4.400 1603.080 1767.255 1603.760 ;
        RECT 1.445 1600.400 1767.255 1603.080 ;
        RECT 4.400 1599.000 1767.255 1600.400 ;
        RECT 1.445 1597.000 1767.255 1599.000 ;
        RECT 4.400 1596.320 1767.255 1597.000 ;
        RECT 4.400 1595.600 1762.995 1596.320 ;
        RECT 1.445 1594.920 1762.995 1595.600 ;
        RECT 1.445 1593.600 1767.255 1594.920 ;
        RECT 4.400 1592.200 1767.255 1593.600 ;
        RECT 1.445 1590.200 1767.255 1592.200 ;
        RECT 4.400 1588.800 1767.255 1590.200 ;
        RECT 1.445 1587.480 1767.255 1588.800 ;
        RECT 1.445 1586.800 1762.995 1587.480 ;
        RECT 4.400 1586.080 1762.995 1586.800 ;
        RECT 4.400 1585.400 1767.255 1586.080 ;
        RECT 1.445 1583.400 1767.255 1585.400 ;
        RECT 4.400 1582.000 1767.255 1583.400 ;
        RECT 1.445 1579.320 1767.255 1582.000 ;
        RECT 4.400 1578.640 1767.255 1579.320 ;
        RECT 4.400 1577.920 1762.995 1578.640 ;
        RECT 1.445 1577.240 1762.995 1577.920 ;
        RECT 1.445 1575.920 1767.255 1577.240 ;
        RECT 4.400 1574.520 1767.255 1575.920 ;
        RECT 1.445 1572.520 1767.255 1574.520 ;
        RECT 4.400 1571.120 1767.255 1572.520 ;
        RECT 1.445 1569.800 1767.255 1571.120 ;
        RECT 1.445 1569.120 1762.995 1569.800 ;
        RECT 4.400 1568.400 1762.995 1569.120 ;
        RECT 4.400 1567.720 1767.255 1568.400 ;
        RECT 1.445 1565.720 1767.255 1567.720 ;
        RECT 4.400 1564.320 1767.255 1565.720 ;
        RECT 1.445 1561.640 1767.255 1564.320 ;
        RECT 4.400 1560.960 1767.255 1561.640 ;
        RECT 4.400 1560.240 1762.995 1560.960 ;
        RECT 1.445 1559.560 1762.995 1560.240 ;
        RECT 1.445 1558.240 1767.255 1559.560 ;
        RECT 4.400 1556.840 1767.255 1558.240 ;
        RECT 1.445 1554.840 1767.255 1556.840 ;
        RECT 4.400 1553.440 1767.255 1554.840 ;
        RECT 1.445 1552.120 1767.255 1553.440 ;
        RECT 1.445 1551.440 1762.995 1552.120 ;
        RECT 4.400 1550.720 1762.995 1551.440 ;
        RECT 4.400 1550.040 1767.255 1550.720 ;
        RECT 1.445 1548.040 1767.255 1550.040 ;
        RECT 4.400 1546.640 1767.255 1548.040 ;
        RECT 1.445 1544.640 1767.255 1546.640 ;
        RECT 4.400 1543.240 1767.255 1544.640 ;
        RECT 1.445 1542.600 1767.255 1543.240 ;
        RECT 1.445 1541.200 1762.995 1542.600 ;
        RECT 1.445 1540.560 1767.255 1541.200 ;
        RECT 4.400 1539.160 1767.255 1540.560 ;
        RECT 1.445 1537.160 1767.255 1539.160 ;
        RECT 4.400 1535.760 1767.255 1537.160 ;
        RECT 1.445 1533.760 1767.255 1535.760 ;
        RECT 4.400 1532.360 1762.995 1533.760 ;
        RECT 1.445 1530.360 1767.255 1532.360 ;
        RECT 4.400 1528.960 1767.255 1530.360 ;
        RECT 1.445 1526.960 1767.255 1528.960 ;
        RECT 4.400 1525.560 1767.255 1526.960 ;
        RECT 1.445 1524.920 1767.255 1525.560 ;
        RECT 1.445 1523.520 1762.995 1524.920 ;
        RECT 1.445 1522.880 1767.255 1523.520 ;
        RECT 4.400 1521.480 1767.255 1522.880 ;
        RECT 1.445 1519.480 1767.255 1521.480 ;
        RECT 4.400 1518.080 1767.255 1519.480 ;
        RECT 1.445 1516.080 1767.255 1518.080 ;
        RECT 4.400 1514.680 1762.995 1516.080 ;
        RECT 1.445 1512.680 1767.255 1514.680 ;
        RECT 4.400 1511.280 1767.255 1512.680 ;
        RECT 1.445 1509.280 1767.255 1511.280 ;
        RECT 4.400 1507.880 1767.255 1509.280 ;
        RECT 1.445 1507.240 1767.255 1507.880 ;
        RECT 1.445 1505.880 1762.995 1507.240 ;
        RECT 4.400 1505.840 1762.995 1505.880 ;
        RECT 4.400 1504.480 1767.255 1505.840 ;
        RECT 1.445 1501.800 1767.255 1504.480 ;
        RECT 4.400 1500.400 1767.255 1501.800 ;
        RECT 1.445 1498.400 1767.255 1500.400 ;
        RECT 4.400 1497.000 1762.995 1498.400 ;
        RECT 1.445 1495.000 1767.255 1497.000 ;
        RECT 4.400 1493.600 1767.255 1495.000 ;
        RECT 1.445 1491.600 1767.255 1493.600 ;
        RECT 4.400 1490.200 1767.255 1491.600 ;
        RECT 1.445 1489.560 1767.255 1490.200 ;
        RECT 1.445 1488.200 1762.995 1489.560 ;
        RECT 4.400 1488.160 1762.995 1488.200 ;
        RECT 4.400 1486.800 1767.255 1488.160 ;
        RECT 1.445 1484.800 1767.255 1486.800 ;
        RECT 4.400 1483.400 1767.255 1484.800 ;
        RECT 1.445 1480.720 1767.255 1483.400 ;
        RECT 4.400 1479.320 1762.995 1480.720 ;
        RECT 1.445 1477.320 1767.255 1479.320 ;
        RECT 4.400 1475.920 1767.255 1477.320 ;
        RECT 1.445 1473.920 1767.255 1475.920 ;
        RECT 4.400 1472.520 1767.255 1473.920 ;
        RECT 1.445 1471.880 1767.255 1472.520 ;
        RECT 1.445 1470.520 1762.995 1471.880 ;
        RECT 4.400 1470.480 1762.995 1470.520 ;
        RECT 4.400 1469.120 1767.255 1470.480 ;
        RECT 1.445 1467.120 1767.255 1469.120 ;
        RECT 4.400 1465.720 1767.255 1467.120 ;
        RECT 1.445 1463.040 1767.255 1465.720 ;
        RECT 4.400 1461.640 1762.995 1463.040 ;
        RECT 1.445 1459.640 1767.255 1461.640 ;
        RECT 4.400 1458.240 1767.255 1459.640 ;
        RECT 1.445 1456.240 1767.255 1458.240 ;
        RECT 4.400 1454.840 1767.255 1456.240 ;
        RECT 1.445 1454.200 1767.255 1454.840 ;
        RECT 1.445 1452.840 1762.995 1454.200 ;
        RECT 4.400 1452.800 1762.995 1452.840 ;
        RECT 4.400 1451.440 1767.255 1452.800 ;
        RECT 1.445 1449.440 1767.255 1451.440 ;
        RECT 4.400 1448.040 1767.255 1449.440 ;
        RECT 1.445 1446.040 1767.255 1448.040 ;
        RECT 4.400 1445.360 1767.255 1446.040 ;
        RECT 4.400 1444.640 1762.995 1445.360 ;
        RECT 1.445 1443.960 1762.995 1444.640 ;
        RECT 1.445 1441.960 1767.255 1443.960 ;
        RECT 4.400 1440.560 1767.255 1441.960 ;
        RECT 1.445 1438.560 1767.255 1440.560 ;
        RECT 4.400 1437.160 1767.255 1438.560 ;
        RECT 1.445 1436.520 1767.255 1437.160 ;
        RECT 1.445 1435.160 1762.995 1436.520 ;
        RECT 4.400 1435.120 1762.995 1435.160 ;
        RECT 4.400 1433.760 1767.255 1435.120 ;
        RECT 1.445 1431.760 1767.255 1433.760 ;
        RECT 4.400 1430.360 1767.255 1431.760 ;
        RECT 1.445 1428.360 1767.255 1430.360 ;
        RECT 4.400 1427.680 1767.255 1428.360 ;
        RECT 4.400 1426.960 1762.995 1427.680 ;
        RECT 1.445 1426.280 1762.995 1426.960 ;
        RECT 1.445 1424.960 1767.255 1426.280 ;
        RECT 4.400 1423.560 1767.255 1424.960 ;
        RECT 1.445 1420.880 1767.255 1423.560 ;
        RECT 4.400 1419.480 1767.255 1420.880 ;
        RECT 1.445 1418.160 1767.255 1419.480 ;
        RECT 1.445 1417.480 1762.995 1418.160 ;
        RECT 4.400 1416.760 1762.995 1417.480 ;
        RECT 4.400 1416.080 1767.255 1416.760 ;
        RECT 1.445 1414.080 1767.255 1416.080 ;
        RECT 4.400 1412.680 1767.255 1414.080 ;
        RECT 1.445 1410.680 1767.255 1412.680 ;
        RECT 4.400 1409.320 1767.255 1410.680 ;
        RECT 4.400 1409.280 1762.995 1409.320 ;
        RECT 1.445 1407.920 1762.995 1409.280 ;
        RECT 1.445 1407.280 1767.255 1407.920 ;
        RECT 4.400 1405.880 1767.255 1407.280 ;
        RECT 1.445 1403.200 1767.255 1405.880 ;
        RECT 4.400 1401.800 1767.255 1403.200 ;
        RECT 1.445 1400.480 1767.255 1401.800 ;
        RECT 1.445 1399.800 1762.995 1400.480 ;
        RECT 4.400 1399.080 1762.995 1399.800 ;
        RECT 4.400 1398.400 1767.255 1399.080 ;
        RECT 1.445 1396.400 1767.255 1398.400 ;
        RECT 4.400 1395.000 1767.255 1396.400 ;
        RECT 1.445 1393.000 1767.255 1395.000 ;
        RECT 4.400 1391.640 1767.255 1393.000 ;
        RECT 4.400 1391.600 1762.995 1391.640 ;
        RECT 1.445 1390.240 1762.995 1391.600 ;
        RECT 1.445 1389.600 1767.255 1390.240 ;
        RECT 4.400 1388.200 1767.255 1389.600 ;
        RECT 1.445 1386.200 1767.255 1388.200 ;
        RECT 4.400 1384.800 1767.255 1386.200 ;
        RECT 1.445 1382.800 1767.255 1384.800 ;
        RECT 1.445 1382.120 1762.995 1382.800 ;
        RECT 4.400 1381.400 1762.995 1382.120 ;
        RECT 4.400 1380.720 1767.255 1381.400 ;
        RECT 1.445 1378.720 1767.255 1380.720 ;
        RECT 4.400 1377.320 1767.255 1378.720 ;
        RECT 1.445 1375.320 1767.255 1377.320 ;
        RECT 4.400 1373.960 1767.255 1375.320 ;
        RECT 4.400 1373.920 1762.995 1373.960 ;
        RECT 1.445 1372.560 1762.995 1373.920 ;
        RECT 1.445 1371.920 1767.255 1372.560 ;
        RECT 4.400 1370.520 1767.255 1371.920 ;
        RECT 1.445 1368.520 1767.255 1370.520 ;
        RECT 4.400 1367.120 1767.255 1368.520 ;
        RECT 1.445 1365.120 1767.255 1367.120 ;
        RECT 1.445 1364.440 1762.995 1365.120 ;
        RECT 4.400 1363.720 1762.995 1364.440 ;
        RECT 4.400 1363.040 1767.255 1363.720 ;
        RECT 1.445 1361.040 1767.255 1363.040 ;
        RECT 4.400 1359.640 1767.255 1361.040 ;
        RECT 1.445 1357.640 1767.255 1359.640 ;
        RECT 4.400 1356.280 1767.255 1357.640 ;
        RECT 4.400 1356.240 1762.995 1356.280 ;
        RECT 1.445 1354.880 1762.995 1356.240 ;
        RECT 1.445 1354.240 1767.255 1354.880 ;
        RECT 4.400 1352.840 1767.255 1354.240 ;
        RECT 1.445 1350.840 1767.255 1352.840 ;
        RECT 4.400 1349.440 1767.255 1350.840 ;
        RECT 1.445 1347.440 1767.255 1349.440 ;
        RECT 4.400 1346.040 1762.995 1347.440 ;
        RECT 1.445 1343.360 1767.255 1346.040 ;
        RECT 4.400 1341.960 1767.255 1343.360 ;
        RECT 1.445 1339.960 1767.255 1341.960 ;
        RECT 4.400 1338.600 1767.255 1339.960 ;
        RECT 4.400 1338.560 1762.995 1338.600 ;
        RECT 1.445 1337.200 1762.995 1338.560 ;
        RECT 1.445 1336.560 1767.255 1337.200 ;
        RECT 4.400 1335.160 1767.255 1336.560 ;
        RECT 1.445 1333.160 1767.255 1335.160 ;
        RECT 4.400 1331.760 1767.255 1333.160 ;
        RECT 1.445 1329.760 1767.255 1331.760 ;
        RECT 4.400 1328.360 1762.995 1329.760 ;
        RECT 1.445 1326.360 1767.255 1328.360 ;
        RECT 4.400 1324.960 1767.255 1326.360 ;
        RECT 1.445 1322.280 1767.255 1324.960 ;
        RECT 4.400 1320.920 1767.255 1322.280 ;
        RECT 4.400 1320.880 1762.995 1320.920 ;
        RECT 1.445 1319.520 1762.995 1320.880 ;
        RECT 1.445 1318.880 1767.255 1319.520 ;
        RECT 4.400 1317.480 1767.255 1318.880 ;
        RECT 1.445 1315.480 1767.255 1317.480 ;
        RECT 4.400 1314.080 1767.255 1315.480 ;
        RECT 1.445 1312.080 1767.255 1314.080 ;
        RECT 4.400 1310.680 1762.995 1312.080 ;
        RECT 1.445 1308.680 1767.255 1310.680 ;
        RECT 4.400 1307.280 1767.255 1308.680 ;
        RECT 1.445 1304.600 1767.255 1307.280 ;
        RECT 4.400 1303.200 1767.255 1304.600 ;
        RECT 1.445 1302.560 1767.255 1303.200 ;
        RECT 1.445 1301.200 1762.995 1302.560 ;
        RECT 4.400 1301.160 1762.995 1301.200 ;
        RECT 4.400 1299.800 1767.255 1301.160 ;
        RECT 1.445 1297.800 1767.255 1299.800 ;
        RECT 4.400 1296.400 1767.255 1297.800 ;
        RECT 1.445 1294.400 1767.255 1296.400 ;
        RECT 4.400 1293.720 1767.255 1294.400 ;
        RECT 4.400 1293.000 1762.995 1293.720 ;
        RECT 1.445 1292.320 1762.995 1293.000 ;
        RECT 1.445 1291.000 1767.255 1292.320 ;
        RECT 4.400 1289.600 1767.255 1291.000 ;
        RECT 1.445 1287.600 1767.255 1289.600 ;
        RECT 4.400 1286.200 1767.255 1287.600 ;
        RECT 1.445 1284.880 1767.255 1286.200 ;
        RECT 1.445 1283.520 1762.995 1284.880 ;
        RECT 4.400 1283.480 1762.995 1283.520 ;
        RECT 4.400 1282.120 1767.255 1283.480 ;
        RECT 1.445 1280.120 1767.255 1282.120 ;
        RECT 4.400 1278.720 1767.255 1280.120 ;
        RECT 1.445 1276.720 1767.255 1278.720 ;
        RECT 4.400 1276.040 1767.255 1276.720 ;
        RECT 4.400 1275.320 1762.995 1276.040 ;
        RECT 1.445 1274.640 1762.995 1275.320 ;
        RECT 1.445 1273.320 1767.255 1274.640 ;
        RECT 4.400 1271.920 1767.255 1273.320 ;
        RECT 1.445 1269.920 1767.255 1271.920 ;
        RECT 4.400 1268.520 1767.255 1269.920 ;
        RECT 1.445 1267.200 1767.255 1268.520 ;
        RECT 1.445 1265.840 1762.995 1267.200 ;
        RECT 4.400 1265.800 1762.995 1265.840 ;
        RECT 4.400 1264.440 1767.255 1265.800 ;
        RECT 1.445 1262.440 1767.255 1264.440 ;
        RECT 4.400 1261.040 1767.255 1262.440 ;
        RECT 1.445 1259.040 1767.255 1261.040 ;
        RECT 4.400 1258.360 1767.255 1259.040 ;
        RECT 4.400 1257.640 1762.995 1258.360 ;
        RECT 1.445 1256.960 1762.995 1257.640 ;
        RECT 1.445 1255.640 1767.255 1256.960 ;
        RECT 4.400 1254.240 1767.255 1255.640 ;
        RECT 1.445 1252.240 1767.255 1254.240 ;
        RECT 4.400 1250.840 1767.255 1252.240 ;
        RECT 1.445 1249.520 1767.255 1250.840 ;
        RECT 1.445 1248.840 1762.995 1249.520 ;
        RECT 4.400 1248.120 1762.995 1248.840 ;
        RECT 4.400 1247.440 1767.255 1248.120 ;
        RECT 1.445 1244.760 1767.255 1247.440 ;
        RECT 4.400 1243.360 1767.255 1244.760 ;
        RECT 1.445 1241.360 1767.255 1243.360 ;
        RECT 4.400 1240.680 1767.255 1241.360 ;
        RECT 4.400 1239.960 1762.995 1240.680 ;
        RECT 1.445 1239.280 1762.995 1239.960 ;
        RECT 1.445 1237.960 1767.255 1239.280 ;
        RECT 4.400 1236.560 1767.255 1237.960 ;
        RECT 1.445 1234.560 1767.255 1236.560 ;
        RECT 4.400 1233.160 1767.255 1234.560 ;
        RECT 1.445 1231.840 1767.255 1233.160 ;
        RECT 1.445 1231.160 1762.995 1231.840 ;
        RECT 4.400 1230.440 1762.995 1231.160 ;
        RECT 4.400 1229.760 1767.255 1230.440 ;
        RECT 1.445 1227.760 1767.255 1229.760 ;
        RECT 4.400 1226.360 1767.255 1227.760 ;
        RECT 1.445 1223.680 1767.255 1226.360 ;
        RECT 4.400 1223.000 1767.255 1223.680 ;
        RECT 4.400 1222.280 1762.995 1223.000 ;
        RECT 1.445 1221.600 1762.995 1222.280 ;
        RECT 1.445 1220.280 1767.255 1221.600 ;
        RECT 4.400 1218.880 1767.255 1220.280 ;
        RECT 1.445 1216.880 1767.255 1218.880 ;
        RECT 4.400 1215.480 1767.255 1216.880 ;
        RECT 1.445 1214.160 1767.255 1215.480 ;
        RECT 1.445 1213.480 1762.995 1214.160 ;
        RECT 4.400 1212.760 1762.995 1213.480 ;
        RECT 4.400 1212.080 1767.255 1212.760 ;
        RECT 1.445 1210.080 1767.255 1212.080 ;
        RECT 4.400 1208.680 1767.255 1210.080 ;
        RECT 1.445 1206.000 1767.255 1208.680 ;
        RECT 4.400 1205.320 1767.255 1206.000 ;
        RECT 4.400 1204.600 1762.995 1205.320 ;
        RECT 1.445 1203.920 1762.995 1204.600 ;
        RECT 1.445 1202.600 1767.255 1203.920 ;
        RECT 4.400 1201.200 1767.255 1202.600 ;
        RECT 1.445 1199.200 1767.255 1201.200 ;
        RECT 4.400 1197.800 1767.255 1199.200 ;
        RECT 1.445 1196.480 1767.255 1197.800 ;
        RECT 1.445 1195.800 1762.995 1196.480 ;
        RECT 4.400 1195.080 1762.995 1195.800 ;
        RECT 4.400 1194.400 1767.255 1195.080 ;
        RECT 1.445 1192.400 1767.255 1194.400 ;
        RECT 4.400 1191.000 1767.255 1192.400 ;
        RECT 1.445 1189.000 1767.255 1191.000 ;
        RECT 4.400 1187.600 1767.255 1189.000 ;
        RECT 1.445 1186.960 1767.255 1187.600 ;
        RECT 1.445 1185.560 1762.995 1186.960 ;
        RECT 1.445 1184.920 1767.255 1185.560 ;
        RECT 4.400 1183.520 1767.255 1184.920 ;
        RECT 1.445 1181.520 1767.255 1183.520 ;
        RECT 4.400 1180.120 1767.255 1181.520 ;
        RECT 1.445 1178.120 1767.255 1180.120 ;
        RECT 4.400 1176.720 1762.995 1178.120 ;
        RECT 1.445 1174.720 1767.255 1176.720 ;
        RECT 4.400 1173.320 1767.255 1174.720 ;
        RECT 1.445 1171.320 1767.255 1173.320 ;
        RECT 4.400 1169.920 1767.255 1171.320 ;
        RECT 1.445 1169.280 1767.255 1169.920 ;
        RECT 1.445 1167.880 1762.995 1169.280 ;
        RECT 1.445 1167.240 1767.255 1167.880 ;
        RECT 4.400 1165.840 1767.255 1167.240 ;
        RECT 1.445 1163.840 1767.255 1165.840 ;
        RECT 4.400 1162.440 1767.255 1163.840 ;
        RECT 1.445 1160.440 1767.255 1162.440 ;
        RECT 4.400 1159.040 1762.995 1160.440 ;
        RECT 1.445 1157.040 1767.255 1159.040 ;
        RECT 4.400 1155.640 1767.255 1157.040 ;
        RECT 1.445 1153.640 1767.255 1155.640 ;
        RECT 4.400 1152.240 1767.255 1153.640 ;
        RECT 1.445 1151.600 1767.255 1152.240 ;
        RECT 1.445 1150.240 1762.995 1151.600 ;
        RECT 4.400 1150.200 1762.995 1150.240 ;
        RECT 4.400 1148.840 1767.255 1150.200 ;
        RECT 1.445 1146.160 1767.255 1148.840 ;
        RECT 4.400 1144.760 1767.255 1146.160 ;
        RECT 1.445 1142.760 1767.255 1144.760 ;
        RECT 4.400 1141.360 1762.995 1142.760 ;
        RECT 1.445 1139.360 1767.255 1141.360 ;
        RECT 4.400 1137.960 1767.255 1139.360 ;
        RECT 1.445 1135.960 1767.255 1137.960 ;
        RECT 4.400 1134.560 1767.255 1135.960 ;
        RECT 1.445 1133.920 1767.255 1134.560 ;
        RECT 1.445 1132.560 1762.995 1133.920 ;
        RECT 4.400 1132.520 1762.995 1132.560 ;
        RECT 4.400 1131.160 1767.255 1132.520 ;
        RECT 1.445 1129.160 1767.255 1131.160 ;
        RECT 4.400 1127.760 1767.255 1129.160 ;
        RECT 1.445 1125.080 1767.255 1127.760 ;
        RECT 4.400 1123.680 1762.995 1125.080 ;
        RECT 1.445 1121.680 1767.255 1123.680 ;
        RECT 4.400 1120.280 1767.255 1121.680 ;
        RECT 1.445 1118.280 1767.255 1120.280 ;
        RECT 4.400 1116.880 1767.255 1118.280 ;
        RECT 1.445 1116.240 1767.255 1116.880 ;
        RECT 1.445 1114.880 1762.995 1116.240 ;
        RECT 4.400 1114.840 1762.995 1114.880 ;
        RECT 4.400 1113.480 1767.255 1114.840 ;
        RECT 1.445 1111.480 1767.255 1113.480 ;
        RECT 4.400 1110.080 1767.255 1111.480 ;
        RECT 1.445 1107.400 1767.255 1110.080 ;
        RECT 4.400 1106.000 1762.995 1107.400 ;
        RECT 1.445 1104.000 1767.255 1106.000 ;
        RECT 4.400 1102.600 1767.255 1104.000 ;
        RECT 1.445 1100.600 1767.255 1102.600 ;
        RECT 4.400 1099.200 1767.255 1100.600 ;
        RECT 1.445 1098.560 1767.255 1099.200 ;
        RECT 1.445 1097.200 1762.995 1098.560 ;
        RECT 4.400 1097.160 1762.995 1097.200 ;
        RECT 4.400 1095.800 1767.255 1097.160 ;
        RECT 1.445 1093.800 1767.255 1095.800 ;
        RECT 4.400 1092.400 1767.255 1093.800 ;
        RECT 1.445 1090.400 1767.255 1092.400 ;
        RECT 4.400 1089.720 1767.255 1090.400 ;
        RECT 4.400 1089.000 1762.995 1089.720 ;
        RECT 1.445 1088.320 1762.995 1089.000 ;
        RECT 1.445 1086.320 1767.255 1088.320 ;
        RECT 4.400 1084.920 1767.255 1086.320 ;
        RECT 1.445 1082.920 1767.255 1084.920 ;
        RECT 4.400 1081.520 1767.255 1082.920 ;
        RECT 1.445 1080.880 1767.255 1081.520 ;
        RECT 1.445 1079.520 1762.995 1080.880 ;
        RECT 4.400 1079.480 1762.995 1079.520 ;
        RECT 4.400 1078.120 1767.255 1079.480 ;
        RECT 1.445 1076.120 1767.255 1078.120 ;
        RECT 4.400 1074.720 1767.255 1076.120 ;
        RECT 1.445 1072.720 1767.255 1074.720 ;
        RECT 4.400 1072.040 1767.255 1072.720 ;
        RECT 4.400 1071.320 1762.995 1072.040 ;
        RECT 1.445 1070.640 1762.995 1071.320 ;
        RECT 1.445 1069.320 1767.255 1070.640 ;
        RECT 4.400 1067.920 1767.255 1069.320 ;
        RECT 1.445 1065.240 1767.255 1067.920 ;
        RECT 4.400 1063.840 1767.255 1065.240 ;
        RECT 1.445 1062.520 1767.255 1063.840 ;
        RECT 1.445 1061.840 1762.995 1062.520 ;
        RECT 4.400 1061.120 1762.995 1061.840 ;
        RECT 4.400 1060.440 1767.255 1061.120 ;
        RECT 1.445 1058.440 1767.255 1060.440 ;
        RECT 4.400 1057.040 1767.255 1058.440 ;
        RECT 1.445 1055.040 1767.255 1057.040 ;
        RECT 4.400 1053.680 1767.255 1055.040 ;
        RECT 4.400 1053.640 1762.995 1053.680 ;
        RECT 1.445 1052.280 1762.995 1053.640 ;
        RECT 1.445 1051.640 1767.255 1052.280 ;
        RECT 4.400 1050.240 1767.255 1051.640 ;
        RECT 1.445 1047.560 1767.255 1050.240 ;
        RECT 4.400 1046.160 1767.255 1047.560 ;
        RECT 1.445 1044.840 1767.255 1046.160 ;
        RECT 1.445 1044.160 1762.995 1044.840 ;
        RECT 4.400 1043.440 1762.995 1044.160 ;
        RECT 4.400 1042.760 1767.255 1043.440 ;
        RECT 1.445 1040.760 1767.255 1042.760 ;
        RECT 4.400 1039.360 1767.255 1040.760 ;
        RECT 1.445 1037.360 1767.255 1039.360 ;
        RECT 4.400 1036.000 1767.255 1037.360 ;
        RECT 4.400 1035.960 1762.995 1036.000 ;
        RECT 1.445 1034.600 1762.995 1035.960 ;
        RECT 1.445 1033.960 1767.255 1034.600 ;
        RECT 4.400 1032.560 1767.255 1033.960 ;
        RECT 1.445 1030.560 1767.255 1032.560 ;
        RECT 4.400 1029.160 1767.255 1030.560 ;
        RECT 1.445 1027.160 1767.255 1029.160 ;
        RECT 1.445 1026.480 1762.995 1027.160 ;
        RECT 4.400 1025.760 1762.995 1026.480 ;
        RECT 4.400 1025.080 1767.255 1025.760 ;
        RECT 1.445 1023.080 1767.255 1025.080 ;
        RECT 4.400 1021.680 1767.255 1023.080 ;
        RECT 1.445 1019.680 1767.255 1021.680 ;
        RECT 4.400 1018.320 1767.255 1019.680 ;
        RECT 4.400 1018.280 1762.995 1018.320 ;
        RECT 1.445 1016.920 1762.995 1018.280 ;
        RECT 1.445 1016.280 1767.255 1016.920 ;
        RECT 4.400 1014.880 1767.255 1016.280 ;
        RECT 1.445 1012.880 1767.255 1014.880 ;
        RECT 4.400 1011.480 1767.255 1012.880 ;
        RECT 1.445 1009.480 1767.255 1011.480 ;
        RECT 1.445 1008.800 1762.995 1009.480 ;
        RECT 4.400 1008.080 1762.995 1008.800 ;
        RECT 4.400 1007.400 1767.255 1008.080 ;
        RECT 1.445 1005.400 1767.255 1007.400 ;
        RECT 4.400 1004.000 1767.255 1005.400 ;
        RECT 1.445 1002.000 1767.255 1004.000 ;
        RECT 4.400 1000.640 1767.255 1002.000 ;
        RECT 4.400 1000.600 1762.995 1000.640 ;
        RECT 1.445 999.240 1762.995 1000.600 ;
        RECT 1.445 998.600 1767.255 999.240 ;
        RECT 4.400 997.200 1767.255 998.600 ;
        RECT 1.445 995.200 1767.255 997.200 ;
        RECT 4.400 993.800 1767.255 995.200 ;
        RECT 1.445 991.800 1767.255 993.800 ;
        RECT 4.400 990.400 1762.995 991.800 ;
        RECT 1.445 987.720 1767.255 990.400 ;
        RECT 4.400 986.320 1767.255 987.720 ;
        RECT 1.445 984.320 1767.255 986.320 ;
        RECT 4.400 982.960 1767.255 984.320 ;
        RECT 4.400 982.920 1762.995 982.960 ;
        RECT 1.445 981.560 1762.995 982.920 ;
        RECT 1.445 980.920 1767.255 981.560 ;
        RECT 4.400 979.520 1767.255 980.920 ;
        RECT 1.445 977.520 1767.255 979.520 ;
        RECT 4.400 976.120 1767.255 977.520 ;
        RECT 1.445 974.120 1767.255 976.120 ;
        RECT 4.400 972.720 1762.995 974.120 ;
        RECT 1.445 970.720 1767.255 972.720 ;
        RECT 4.400 969.320 1767.255 970.720 ;
        RECT 1.445 966.640 1767.255 969.320 ;
        RECT 4.400 965.280 1767.255 966.640 ;
        RECT 4.400 965.240 1762.995 965.280 ;
        RECT 1.445 963.880 1762.995 965.240 ;
        RECT 1.445 963.240 1767.255 963.880 ;
        RECT 4.400 961.840 1767.255 963.240 ;
        RECT 1.445 959.840 1767.255 961.840 ;
        RECT 4.400 958.440 1767.255 959.840 ;
        RECT 1.445 956.440 1767.255 958.440 ;
        RECT 4.400 955.040 1762.995 956.440 ;
        RECT 1.445 953.040 1767.255 955.040 ;
        RECT 4.400 951.640 1767.255 953.040 ;
        RECT 1.445 948.960 1767.255 951.640 ;
        RECT 4.400 947.560 1767.255 948.960 ;
        RECT 1.445 946.920 1767.255 947.560 ;
        RECT 1.445 945.560 1762.995 946.920 ;
        RECT 4.400 945.520 1762.995 945.560 ;
        RECT 4.400 944.160 1767.255 945.520 ;
        RECT 1.445 942.160 1767.255 944.160 ;
        RECT 4.400 940.760 1767.255 942.160 ;
        RECT 1.445 938.760 1767.255 940.760 ;
        RECT 4.400 938.080 1767.255 938.760 ;
        RECT 4.400 937.360 1762.995 938.080 ;
        RECT 1.445 936.680 1762.995 937.360 ;
        RECT 1.445 935.360 1767.255 936.680 ;
        RECT 4.400 933.960 1767.255 935.360 ;
        RECT 1.445 931.960 1767.255 933.960 ;
        RECT 4.400 930.560 1767.255 931.960 ;
        RECT 1.445 929.240 1767.255 930.560 ;
        RECT 1.445 927.880 1762.995 929.240 ;
        RECT 4.400 927.840 1762.995 927.880 ;
        RECT 4.400 926.480 1767.255 927.840 ;
        RECT 1.445 924.480 1767.255 926.480 ;
        RECT 4.400 923.080 1767.255 924.480 ;
        RECT 1.445 921.080 1767.255 923.080 ;
        RECT 4.400 920.400 1767.255 921.080 ;
        RECT 4.400 919.680 1762.995 920.400 ;
        RECT 1.445 919.000 1762.995 919.680 ;
        RECT 1.445 917.680 1767.255 919.000 ;
        RECT 4.400 916.280 1767.255 917.680 ;
        RECT 1.445 914.280 1767.255 916.280 ;
        RECT 4.400 912.880 1767.255 914.280 ;
        RECT 1.445 911.560 1767.255 912.880 ;
        RECT 1.445 910.200 1762.995 911.560 ;
        RECT 4.400 910.160 1762.995 910.200 ;
        RECT 4.400 908.800 1767.255 910.160 ;
        RECT 1.445 906.800 1767.255 908.800 ;
        RECT 4.400 905.400 1767.255 906.800 ;
        RECT 1.445 903.400 1767.255 905.400 ;
        RECT 4.400 902.720 1767.255 903.400 ;
        RECT 4.400 902.000 1762.995 902.720 ;
        RECT 1.445 901.320 1762.995 902.000 ;
        RECT 1.445 900.000 1767.255 901.320 ;
        RECT 4.400 898.600 1767.255 900.000 ;
        RECT 1.445 896.600 1767.255 898.600 ;
        RECT 4.400 895.200 1767.255 896.600 ;
        RECT 1.445 893.880 1767.255 895.200 ;
        RECT 1.445 893.200 1762.995 893.880 ;
        RECT 4.400 892.480 1762.995 893.200 ;
        RECT 4.400 891.800 1767.255 892.480 ;
        RECT 1.445 889.120 1767.255 891.800 ;
        RECT 4.400 887.720 1767.255 889.120 ;
        RECT 1.445 885.720 1767.255 887.720 ;
        RECT 4.400 885.040 1767.255 885.720 ;
        RECT 4.400 884.320 1762.995 885.040 ;
        RECT 1.445 883.640 1762.995 884.320 ;
        RECT 1.445 882.320 1767.255 883.640 ;
        RECT 4.400 880.920 1767.255 882.320 ;
        RECT 1.445 878.920 1767.255 880.920 ;
        RECT 4.400 877.520 1767.255 878.920 ;
        RECT 1.445 876.200 1767.255 877.520 ;
        RECT 1.445 875.520 1762.995 876.200 ;
        RECT 4.400 874.800 1762.995 875.520 ;
        RECT 4.400 874.120 1767.255 874.800 ;
        RECT 1.445 872.120 1767.255 874.120 ;
        RECT 4.400 870.720 1767.255 872.120 ;
        RECT 1.445 868.040 1767.255 870.720 ;
        RECT 4.400 867.360 1767.255 868.040 ;
        RECT 4.400 866.640 1762.995 867.360 ;
        RECT 1.445 865.960 1762.995 866.640 ;
        RECT 1.445 864.640 1767.255 865.960 ;
        RECT 4.400 863.240 1767.255 864.640 ;
        RECT 1.445 861.240 1767.255 863.240 ;
        RECT 4.400 859.840 1767.255 861.240 ;
        RECT 1.445 858.520 1767.255 859.840 ;
        RECT 1.445 857.840 1762.995 858.520 ;
        RECT 4.400 857.120 1762.995 857.840 ;
        RECT 4.400 856.440 1767.255 857.120 ;
        RECT 1.445 854.440 1767.255 856.440 ;
        RECT 4.400 853.040 1767.255 854.440 ;
        RECT 1.445 850.360 1767.255 853.040 ;
        RECT 4.400 849.680 1767.255 850.360 ;
        RECT 4.400 848.960 1762.995 849.680 ;
        RECT 1.445 848.280 1762.995 848.960 ;
        RECT 1.445 846.960 1767.255 848.280 ;
        RECT 4.400 845.560 1767.255 846.960 ;
        RECT 1.445 843.560 1767.255 845.560 ;
        RECT 4.400 842.160 1767.255 843.560 ;
        RECT 1.445 840.840 1767.255 842.160 ;
        RECT 1.445 840.160 1762.995 840.840 ;
        RECT 4.400 839.440 1762.995 840.160 ;
        RECT 4.400 838.760 1767.255 839.440 ;
        RECT 1.445 836.760 1767.255 838.760 ;
        RECT 4.400 835.360 1767.255 836.760 ;
        RECT 1.445 833.360 1767.255 835.360 ;
        RECT 4.400 831.960 1767.255 833.360 ;
        RECT 1.445 831.320 1767.255 831.960 ;
        RECT 1.445 829.920 1762.995 831.320 ;
        RECT 1.445 829.280 1767.255 829.920 ;
        RECT 4.400 827.880 1767.255 829.280 ;
        RECT 1.445 825.880 1767.255 827.880 ;
        RECT 4.400 824.480 1767.255 825.880 ;
        RECT 1.445 822.480 1767.255 824.480 ;
        RECT 4.400 821.080 1762.995 822.480 ;
        RECT 1.445 819.080 1767.255 821.080 ;
        RECT 4.400 817.680 1767.255 819.080 ;
        RECT 1.445 815.680 1767.255 817.680 ;
        RECT 4.400 814.280 1767.255 815.680 ;
        RECT 1.445 813.640 1767.255 814.280 ;
        RECT 1.445 812.240 1762.995 813.640 ;
        RECT 1.445 811.600 1767.255 812.240 ;
        RECT 4.400 810.200 1767.255 811.600 ;
        RECT 1.445 808.200 1767.255 810.200 ;
        RECT 4.400 806.800 1767.255 808.200 ;
        RECT 1.445 804.800 1767.255 806.800 ;
        RECT 4.400 803.400 1762.995 804.800 ;
        RECT 1.445 801.400 1767.255 803.400 ;
        RECT 4.400 800.000 1767.255 801.400 ;
        RECT 1.445 798.000 1767.255 800.000 ;
        RECT 4.400 796.600 1767.255 798.000 ;
        RECT 1.445 795.960 1767.255 796.600 ;
        RECT 1.445 794.600 1762.995 795.960 ;
        RECT 4.400 794.560 1762.995 794.600 ;
        RECT 4.400 793.200 1767.255 794.560 ;
        RECT 1.445 790.520 1767.255 793.200 ;
        RECT 4.400 789.120 1767.255 790.520 ;
        RECT 1.445 787.120 1767.255 789.120 ;
        RECT 4.400 785.720 1762.995 787.120 ;
        RECT 1.445 783.720 1767.255 785.720 ;
        RECT 4.400 782.320 1767.255 783.720 ;
        RECT 1.445 780.320 1767.255 782.320 ;
        RECT 4.400 778.920 1767.255 780.320 ;
        RECT 1.445 778.280 1767.255 778.920 ;
        RECT 1.445 776.920 1762.995 778.280 ;
        RECT 4.400 776.880 1762.995 776.920 ;
        RECT 4.400 775.520 1767.255 776.880 ;
        RECT 1.445 773.520 1767.255 775.520 ;
        RECT 4.400 772.120 1767.255 773.520 ;
        RECT 1.445 769.440 1767.255 772.120 ;
        RECT 4.400 768.040 1762.995 769.440 ;
        RECT 1.445 766.040 1767.255 768.040 ;
        RECT 4.400 764.640 1767.255 766.040 ;
        RECT 1.445 762.640 1767.255 764.640 ;
        RECT 4.400 761.240 1767.255 762.640 ;
        RECT 1.445 760.600 1767.255 761.240 ;
        RECT 1.445 759.240 1762.995 760.600 ;
        RECT 4.400 759.200 1762.995 759.240 ;
        RECT 4.400 757.840 1767.255 759.200 ;
        RECT 1.445 755.840 1767.255 757.840 ;
        RECT 4.400 754.440 1767.255 755.840 ;
        RECT 1.445 751.760 1767.255 754.440 ;
        RECT 4.400 750.360 1762.995 751.760 ;
        RECT 1.445 748.360 1767.255 750.360 ;
        RECT 4.400 746.960 1767.255 748.360 ;
        RECT 1.445 744.960 1767.255 746.960 ;
        RECT 4.400 743.560 1767.255 744.960 ;
        RECT 1.445 742.920 1767.255 743.560 ;
        RECT 1.445 741.560 1762.995 742.920 ;
        RECT 4.400 741.520 1762.995 741.560 ;
        RECT 4.400 740.160 1767.255 741.520 ;
        RECT 1.445 738.160 1767.255 740.160 ;
        RECT 4.400 736.760 1767.255 738.160 ;
        RECT 1.445 734.760 1767.255 736.760 ;
        RECT 4.400 734.080 1767.255 734.760 ;
        RECT 4.400 733.360 1762.995 734.080 ;
        RECT 1.445 732.680 1762.995 733.360 ;
        RECT 1.445 730.680 1767.255 732.680 ;
        RECT 4.400 729.280 1767.255 730.680 ;
        RECT 1.445 727.280 1767.255 729.280 ;
        RECT 4.400 725.880 1767.255 727.280 ;
        RECT 1.445 725.240 1767.255 725.880 ;
        RECT 1.445 723.880 1762.995 725.240 ;
        RECT 4.400 723.840 1762.995 723.880 ;
        RECT 4.400 722.480 1767.255 723.840 ;
        RECT 1.445 720.480 1767.255 722.480 ;
        RECT 4.400 719.080 1767.255 720.480 ;
        RECT 1.445 717.080 1767.255 719.080 ;
        RECT 4.400 716.400 1767.255 717.080 ;
        RECT 4.400 715.680 1762.995 716.400 ;
        RECT 1.445 715.000 1762.995 715.680 ;
        RECT 1.445 713.680 1767.255 715.000 ;
        RECT 4.400 712.280 1767.255 713.680 ;
        RECT 1.445 709.600 1767.255 712.280 ;
        RECT 4.400 708.200 1767.255 709.600 ;
        RECT 1.445 706.880 1767.255 708.200 ;
        RECT 1.445 706.200 1762.995 706.880 ;
        RECT 4.400 705.480 1762.995 706.200 ;
        RECT 4.400 704.800 1767.255 705.480 ;
        RECT 1.445 702.800 1767.255 704.800 ;
        RECT 4.400 701.400 1767.255 702.800 ;
        RECT 1.445 699.400 1767.255 701.400 ;
        RECT 4.400 698.040 1767.255 699.400 ;
        RECT 4.400 698.000 1762.995 698.040 ;
        RECT 1.445 696.640 1762.995 698.000 ;
        RECT 1.445 696.000 1767.255 696.640 ;
        RECT 4.400 694.600 1767.255 696.000 ;
        RECT 1.445 691.920 1767.255 694.600 ;
        RECT 4.400 690.520 1767.255 691.920 ;
        RECT 1.445 689.200 1767.255 690.520 ;
        RECT 1.445 688.520 1762.995 689.200 ;
        RECT 4.400 687.800 1762.995 688.520 ;
        RECT 4.400 687.120 1767.255 687.800 ;
        RECT 1.445 685.120 1767.255 687.120 ;
        RECT 4.400 683.720 1767.255 685.120 ;
        RECT 1.445 681.720 1767.255 683.720 ;
        RECT 4.400 680.360 1767.255 681.720 ;
        RECT 4.400 680.320 1762.995 680.360 ;
        RECT 1.445 678.960 1762.995 680.320 ;
        RECT 1.445 678.320 1767.255 678.960 ;
        RECT 4.400 676.920 1767.255 678.320 ;
        RECT 1.445 674.920 1767.255 676.920 ;
        RECT 4.400 673.520 1767.255 674.920 ;
        RECT 1.445 671.520 1767.255 673.520 ;
        RECT 1.445 670.840 1762.995 671.520 ;
        RECT 4.400 670.120 1762.995 670.840 ;
        RECT 4.400 669.440 1767.255 670.120 ;
        RECT 1.445 667.440 1767.255 669.440 ;
        RECT 4.400 666.040 1767.255 667.440 ;
        RECT 1.445 664.040 1767.255 666.040 ;
        RECT 4.400 662.680 1767.255 664.040 ;
        RECT 4.400 662.640 1762.995 662.680 ;
        RECT 1.445 661.280 1762.995 662.640 ;
        RECT 1.445 660.640 1767.255 661.280 ;
        RECT 4.400 659.240 1767.255 660.640 ;
        RECT 1.445 657.240 1767.255 659.240 ;
        RECT 4.400 655.840 1767.255 657.240 ;
        RECT 1.445 653.840 1767.255 655.840 ;
        RECT 1.445 653.160 1762.995 653.840 ;
        RECT 4.400 652.440 1762.995 653.160 ;
        RECT 4.400 651.760 1767.255 652.440 ;
        RECT 1.445 649.760 1767.255 651.760 ;
        RECT 4.400 648.360 1767.255 649.760 ;
        RECT 1.445 646.360 1767.255 648.360 ;
        RECT 4.400 645.000 1767.255 646.360 ;
        RECT 4.400 644.960 1762.995 645.000 ;
        RECT 1.445 643.600 1762.995 644.960 ;
        RECT 1.445 642.960 1767.255 643.600 ;
        RECT 4.400 641.560 1767.255 642.960 ;
        RECT 1.445 639.560 1767.255 641.560 ;
        RECT 4.400 638.160 1767.255 639.560 ;
        RECT 1.445 636.160 1767.255 638.160 ;
        RECT 4.400 634.760 1762.995 636.160 ;
        RECT 1.445 632.080 1767.255 634.760 ;
        RECT 4.400 630.680 1767.255 632.080 ;
        RECT 1.445 628.680 1767.255 630.680 ;
        RECT 4.400 627.320 1767.255 628.680 ;
        RECT 4.400 627.280 1762.995 627.320 ;
        RECT 1.445 625.920 1762.995 627.280 ;
        RECT 1.445 625.280 1767.255 625.920 ;
        RECT 4.400 623.880 1767.255 625.280 ;
        RECT 1.445 621.880 1767.255 623.880 ;
        RECT 4.400 620.480 1767.255 621.880 ;
        RECT 1.445 618.480 1767.255 620.480 ;
        RECT 4.400 617.080 1762.995 618.480 ;
        RECT 1.445 615.080 1767.255 617.080 ;
        RECT 4.400 613.680 1767.255 615.080 ;
        RECT 1.445 611.000 1767.255 613.680 ;
        RECT 4.400 609.640 1767.255 611.000 ;
        RECT 4.400 609.600 1762.995 609.640 ;
        RECT 1.445 608.240 1762.995 609.600 ;
        RECT 1.445 607.600 1767.255 608.240 ;
        RECT 4.400 606.200 1767.255 607.600 ;
        RECT 1.445 604.200 1767.255 606.200 ;
        RECT 4.400 602.800 1767.255 604.200 ;
        RECT 1.445 600.800 1767.255 602.800 ;
        RECT 4.400 599.400 1762.995 600.800 ;
        RECT 1.445 597.400 1767.255 599.400 ;
        RECT 4.400 596.000 1767.255 597.400 ;
        RECT 1.445 593.320 1767.255 596.000 ;
        RECT 4.400 591.920 1767.255 593.320 ;
        RECT 1.445 591.280 1767.255 591.920 ;
        RECT 1.445 589.920 1762.995 591.280 ;
        RECT 4.400 589.880 1762.995 589.920 ;
        RECT 4.400 588.520 1767.255 589.880 ;
        RECT 1.445 586.520 1767.255 588.520 ;
        RECT 4.400 585.120 1767.255 586.520 ;
        RECT 1.445 583.120 1767.255 585.120 ;
        RECT 4.400 582.440 1767.255 583.120 ;
        RECT 4.400 581.720 1762.995 582.440 ;
        RECT 1.445 581.040 1762.995 581.720 ;
        RECT 1.445 579.720 1767.255 581.040 ;
        RECT 4.400 578.320 1767.255 579.720 ;
        RECT 1.445 576.320 1767.255 578.320 ;
        RECT 4.400 574.920 1767.255 576.320 ;
        RECT 1.445 573.600 1767.255 574.920 ;
        RECT 1.445 572.240 1762.995 573.600 ;
        RECT 4.400 572.200 1762.995 572.240 ;
        RECT 4.400 570.840 1767.255 572.200 ;
        RECT 1.445 568.840 1767.255 570.840 ;
        RECT 4.400 567.440 1767.255 568.840 ;
        RECT 1.445 565.440 1767.255 567.440 ;
        RECT 4.400 564.760 1767.255 565.440 ;
        RECT 4.400 564.040 1762.995 564.760 ;
        RECT 1.445 563.360 1762.995 564.040 ;
        RECT 1.445 562.040 1767.255 563.360 ;
        RECT 4.400 560.640 1767.255 562.040 ;
        RECT 1.445 558.640 1767.255 560.640 ;
        RECT 4.400 557.240 1767.255 558.640 ;
        RECT 1.445 555.920 1767.255 557.240 ;
        RECT 1.445 554.560 1762.995 555.920 ;
        RECT 4.400 554.520 1762.995 554.560 ;
        RECT 4.400 553.160 1767.255 554.520 ;
        RECT 1.445 551.160 1767.255 553.160 ;
        RECT 4.400 549.760 1767.255 551.160 ;
        RECT 1.445 547.760 1767.255 549.760 ;
        RECT 4.400 547.080 1767.255 547.760 ;
        RECT 4.400 546.360 1762.995 547.080 ;
        RECT 1.445 545.680 1762.995 546.360 ;
        RECT 1.445 544.360 1767.255 545.680 ;
        RECT 4.400 542.960 1767.255 544.360 ;
        RECT 1.445 540.960 1767.255 542.960 ;
        RECT 4.400 539.560 1767.255 540.960 ;
        RECT 1.445 538.240 1767.255 539.560 ;
        RECT 1.445 537.560 1762.995 538.240 ;
        RECT 4.400 536.840 1762.995 537.560 ;
        RECT 4.400 536.160 1767.255 536.840 ;
        RECT 1.445 533.480 1767.255 536.160 ;
        RECT 4.400 532.080 1767.255 533.480 ;
        RECT 1.445 530.080 1767.255 532.080 ;
        RECT 4.400 529.400 1767.255 530.080 ;
        RECT 4.400 528.680 1762.995 529.400 ;
        RECT 1.445 528.000 1762.995 528.680 ;
        RECT 1.445 526.680 1767.255 528.000 ;
        RECT 4.400 525.280 1767.255 526.680 ;
        RECT 1.445 523.280 1767.255 525.280 ;
        RECT 4.400 521.880 1767.255 523.280 ;
        RECT 1.445 520.560 1767.255 521.880 ;
        RECT 1.445 519.880 1762.995 520.560 ;
        RECT 4.400 519.160 1762.995 519.880 ;
        RECT 4.400 518.480 1767.255 519.160 ;
        RECT 1.445 516.480 1767.255 518.480 ;
        RECT 4.400 515.080 1767.255 516.480 ;
        RECT 1.445 512.400 1767.255 515.080 ;
        RECT 4.400 511.720 1767.255 512.400 ;
        RECT 4.400 511.000 1762.995 511.720 ;
        RECT 1.445 510.320 1762.995 511.000 ;
        RECT 1.445 509.000 1767.255 510.320 ;
        RECT 4.400 507.600 1767.255 509.000 ;
        RECT 1.445 505.600 1767.255 507.600 ;
        RECT 4.400 504.200 1767.255 505.600 ;
        RECT 1.445 502.880 1767.255 504.200 ;
        RECT 1.445 502.200 1762.995 502.880 ;
        RECT 4.400 501.480 1762.995 502.200 ;
        RECT 4.400 500.800 1767.255 501.480 ;
        RECT 1.445 498.800 1767.255 500.800 ;
        RECT 4.400 497.400 1767.255 498.800 ;
        RECT 1.445 494.720 1767.255 497.400 ;
        RECT 4.400 494.040 1767.255 494.720 ;
        RECT 4.400 493.320 1762.995 494.040 ;
        RECT 1.445 492.640 1762.995 493.320 ;
        RECT 1.445 491.320 1767.255 492.640 ;
        RECT 4.400 489.920 1767.255 491.320 ;
        RECT 1.445 487.920 1767.255 489.920 ;
        RECT 4.400 486.520 1767.255 487.920 ;
        RECT 1.445 485.200 1767.255 486.520 ;
        RECT 1.445 484.520 1762.995 485.200 ;
        RECT 4.400 483.800 1762.995 484.520 ;
        RECT 4.400 483.120 1767.255 483.800 ;
        RECT 1.445 481.120 1767.255 483.120 ;
        RECT 4.400 479.720 1767.255 481.120 ;
        RECT 1.445 477.720 1767.255 479.720 ;
        RECT 4.400 476.320 1767.255 477.720 ;
        RECT 1.445 475.680 1767.255 476.320 ;
        RECT 1.445 474.280 1762.995 475.680 ;
        RECT 1.445 473.640 1767.255 474.280 ;
        RECT 4.400 472.240 1767.255 473.640 ;
        RECT 1.445 470.240 1767.255 472.240 ;
        RECT 4.400 468.840 1767.255 470.240 ;
        RECT 1.445 466.840 1767.255 468.840 ;
        RECT 4.400 465.440 1762.995 466.840 ;
        RECT 1.445 463.440 1767.255 465.440 ;
        RECT 4.400 462.040 1767.255 463.440 ;
        RECT 1.445 460.040 1767.255 462.040 ;
        RECT 4.400 458.640 1767.255 460.040 ;
        RECT 1.445 458.000 1767.255 458.640 ;
        RECT 1.445 456.600 1762.995 458.000 ;
        RECT 1.445 455.960 1767.255 456.600 ;
        RECT 4.400 454.560 1767.255 455.960 ;
        RECT 1.445 452.560 1767.255 454.560 ;
        RECT 4.400 451.160 1767.255 452.560 ;
        RECT 1.445 449.160 1767.255 451.160 ;
        RECT 4.400 447.760 1762.995 449.160 ;
        RECT 1.445 445.760 1767.255 447.760 ;
        RECT 4.400 444.360 1767.255 445.760 ;
        RECT 1.445 442.360 1767.255 444.360 ;
        RECT 4.400 440.960 1767.255 442.360 ;
        RECT 1.445 440.320 1767.255 440.960 ;
        RECT 1.445 438.960 1762.995 440.320 ;
        RECT 4.400 438.920 1762.995 438.960 ;
        RECT 4.400 437.560 1767.255 438.920 ;
        RECT 1.445 434.880 1767.255 437.560 ;
        RECT 4.400 433.480 1767.255 434.880 ;
        RECT 1.445 431.480 1767.255 433.480 ;
        RECT 4.400 430.080 1762.995 431.480 ;
        RECT 1.445 428.080 1767.255 430.080 ;
        RECT 4.400 426.680 1767.255 428.080 ;
        RECT 1.445 424.680 1767.255 426.680 ;
        RECT 4.400 423.280 1767.255 424.680 ;
        RECT 1.445 422.640 1767.255 423.280 ;
        RECT 1.445 421.280 1762.995 422.640 ;
        RECT 4.400 421.240 1762.995 421.280 ;
        RECT 4.400 419.880 1767.255 421.240 ;
        RECT 1.445 417.880 1767.255 419.880 ;
        RECT 4.400 416.480 1767.255 417.880 ;
        RECT 1.445 413.800 1767.255 416.480 ;
        RECT 4.400 412.400 1762.995 413.800 ;
        RECT 1.445 410.400 1767.255 412.400 ;
        RECT 4.400 409.000 1767.255 410.400 ;
        RECT 1.445 407.000 1767.255 409.000 ;
        RECT 4.400 405.600 1767.255 407.000 ;
        RECT 1.445 404.960 1767.255 405.600 ;
        RECT 1.445 403.600 1762.995 404.960 ;
        RECT 4.400 403.560 1762.995 403.600 ;
        RECT 4.400 402.200 1767.255 403.560 ;
        RECT 1.445 400.200 1767.255 402.200 ;
        RECT 4.400 398.800 1767.255 400.200 ;
        RECT 1.445 396.120 1767.255 398.800 ;
        RECT 4.400 394.720 1762.995 396.120 ;
        RECT 1.445 392.720 1767.255 394.720 ;
        RECT 4.400 391.320 1767.255 392.720 ;
        RECT 1.445 389.320 1767.255 391.320 ;
        RECT 4.400 387.920 1767.255 389.320 ;
        RECT 1.445 387.280 1767.255 387.920 ;
        RECT 1.445 385.920 1762.995 387.280 ;
        RECT 4.400 385.880 1762.995 385.920 ;
        RECT 4.400 384.520 1767.255 385.880 ;
        RECT 1.445 382.520 1767.255 384.520 ;
        RECT 4.400 381.120 1767.255 382.520 ;
        RECT 1.445 379.120 1767.255 381.120 ;
        RECT 4.400 378.440 1767.255 379.120 ;
        RECT 4.400 377.720 1762.995 378.440 ;
        RECT 1.445 377.040 1762.995 377.720 ;
        RECT 1.445 375.040 1767.255 377.040 ;
        RECT 4.400 373.640 1767.255 375.040 ;
        RECT 1.445 371.640 1767.255 373.640 ;
        RECT 4.400 370.240 1767.255 371.640 ;
        RECT 1.445 369.600 1767.255 370.240 ;
        RECT 1.445 368.240 1762.995 369.600 ;
        RECT 4.400 368.200 1762.995 368.240 ;
        RECT 4.400 366.840 1767.255 368.200 ;
        RECT 1.445 364.840 1767.255 366.840 ;
        RECT 4.400 363.440 1767.255 364.840 ;
        RECT 1.445 361.440 1767.255 363.440 ;
        RECT 4.400 360.760 1767.255 361.440 ;
        RECT 4.400 360.040 1762.995 360.760 ;
        RECT 1.445 359.360 1762.995 360.040 ;
        RECT 1.445 358.040 1767.255 359.360 ;
        RECT 4.400 356.640 1767.255 358.040 ;
        RECT 1.445 353.960 1767.255 356.640 ;
        RECT 4.400 352.560 1767.255 353.960 ;
        RECT 1.445 351.240 1767.255 352.560 ;
        RECT 1.445 350.560 1762.995 351.240 ;
        RECT 4.400 349.840 1762.995 350.560 ;
        RECT 4.400 349.160 1767.255 349.840 ;
        RECT 1.445 347.160 1767.255 349.160 ;
        RECT 4.400 345.760 1767.255 347.160 ;
        RECT 1.445 343.760 1767.255 345.760 ;
        RECT 4.400 342.400 1767.255 343.760 ;
        RECT 4.400 342.360 1762.995 342.400 ;
        RECT 1.445 341.000 1762.995 342.360 ;
        RECT 1.445 340.360 1767.255 341.000 ;
        RECT 4.400 338.960 1767.255 340.360 ;
        RECT 1.445 336.280 1767.255 338.960 ;
        RECT 4.400 334.880 1767.255 336.280 ;
        RECT 1.445 333.560 1767.255 334.880 ;
        RECT 1.445 332.880 1762.995 333.560 ;
        RECT 4.400 332.160 1762.995 332.880 ;
        RECT 4.400 331.480 1767.255 332.160 ;
        RECT 1.445 329.480 1767.255 331.480 ;
        RECT 4.400 328.080 1767.255 329.480 ;
        RECT 1.445 326.080 1767.255 328.080 ;
        RECT 4.400 324.720 1767.255 326.080 ;
        RECT 4.400 324.680 1762.995 324.720 ;
        RECT 1.445 323.320 1762.995 324.680 ;
        RECT 1.445 322.680 1767.255 323.320 ;
        RECT 4.400 321.280 1767.255 322.680 ;
        RECT 1.445 319.280 1767.255 321.280 ;
        RECT 4.400 317.880 1767.255 319.280 ;
        RECT 1.445 315.880 1767.255 317.880 ;
        RECT 1.445 315.200 1762.995 315.880 ;
        RECT 4.400 314.480 1762.995 315.200 ;
        RECT 4.400 313.800 1767.255 314.480 ;
        RECT 1.445 311.800 1767.255 313.800 ;
        RECT 4.400 310.400 1767.255 311.800 ;
        RECT 1.445 308.400 1767.255 310.400 ;
        RECT 4.400 307.040 1767.255 308.400 ;
        RECT 4.400 307.000 1762.995 307.040 ;
        RECT 1.445 305.640 1762.995 307.000 ;
        RECT 1.445 305.000 1767.255 305.640 ;
        RECT 4.400 303.600 1767.255 305.000 ;
        RECT 1.445 301.600 1767.255 303.600 ;
        RECT 4.400 300.200 1767.255 301.600 ;
        RECT 1.445 298.200 1767.255 300.200 ;
        RECT 1.445 297.520 1762.995 298.200 ;
        RECT 4.400 296.800 1762.995 297.520 ;
        RECT 4.400 296.120 1767.255 296.800 ;
        RECT 1.445 294.120 1767.255 296.120 ;
        RECT 4.400 292.720 1767.255 294.120 ;
        RECT 1.445 290.720 1767.255 292.720 ;
        RECT 4.400 289.360 1767.255 290.720 ;
        RECT 4.400 289.320 1762.995 289.360 ;
        RECT 1.445 287.960 1762.995 289.320 ;
        RECT 1.445 287.320 1767.255 287.960 ;
        RECT 4.400 285.920 1767.255 287.320 ;
        RECT 1.445 283.920 1767.255 285.920 ;
        RECT 4.400 282.520 1767.255 283.920 ;
        RECT 1.445 280.520 1767.255 282.520 ;
        RECT 4.400 279.120 1762.995 280.520 ;
        RECT 1.445 276.440 1767.255 279.120 ;
        RECT 4.400 275.040 1767.255 276.440 ;
        RECT 1.445 273.040 1767.255 275.040 ;
        RECT 4.400 271.680 1767.255 273.040 ;
        RECT 4.400 271.640 1762.995 271.680 ;
        RECT 1.445 270.280 1762.995 271.640 ;
        RECT 1.445 269.640 1767.255 270.280 ;
        RECT 4.400 268.240 1767.255 269.640 ;
        RECT 1.445 266.240 1767.255 268.240 ;
        RECT 4.400 264.840 1767.255 266.240 ;
        RECT 1.445 262.840 1767.255 264.840 ;
        RECT 4.400 261.440 1762.995 262.840 ;
        RECT 1.445 259.440 1767.255 261.440 ;
        RECT 4.400 258.040 1767.255 259.440 ;
        RECT 1.445 255.360 1767.255 258.040 ;
        RECT 4.400 254.000 1767.255 255.360 ;
        RECT 4.400 253.960 1762.995 254.000 ;
        RECT 1.445 252.600 1762.995 253.960 ;
        RECT 1.445 251.960 1767.255 252.600 ;
        RECT 4.400 250.560 1767.255 251.960 ;
        RECT 1.445 248.560 1767.255 250.560 ;
        RECT 4.400 247.160 1767.255 248.560 ;
        RECT 1.445 245.160 1767.255 247.160 ;
        RECT 4.400 243.760 1762.995 245.160 ;
        RECT 1.445 241.760 1767.255 243.760 ;
        RECT 4.400 240.360 1767.255 241.760 ;
        RECT 1.445 237.680 1767.255 240.360 ;
        RECT 4.400 236.280 1767.255 237.680 ;
        RECT 1.445 235.640 1767.255 236.280 ;
        RECT 1.445 234.280 1762.995 235.640 ;
        RECT 4.400 234.240 1762.995 234.280 ;
        RECT 4.400 232.880 1767.255 234.240 ;
        RECT 1.445 230.880 1767.255 232.880 ;
        RECT 4.400 229.480 1767.255 230.880 ;
        RECT 1.445 227.480 1767.255 229.480 ;
        RECT 4.400 226.800 1767.255 227.480 ;
        RECT 4.400 226.080 1762.995 226.800 ;
        RECT 1.445 225.400 1762.995 226.080 ;
        RECT 1.445 224.080 1767.255 225.400 ;
        RECT 4.400 222.680 1767.255 224.080 ;
        RECT 1.445 220.680 1767.255 222.680 ;
        RECT 4.400 219.280 1767.255 220.680 ;
        RECT 1.445 217.960 1767.255 219.280 ;
        RECT 1.445 216.600 1762.995 217.960 ;
        RECT 4.400 216.560 1762.995 216.600 ;
        RECT 4.400 215.200 1767.255 216.560 ;
        RECT 1.445 213.200 1767.255 215.200 ;
        RECT 4.400 211.800 1767.255 213.200 ;
        RECT 1.445 209.800 1767.255 211.800 ;
        RECT 4.400 209.120 1767.255 209.800 ;
        RECT 4.400 208.400 1762.995 209.120 ;
        RECT 1.445 207.720 1762.995 208.400 ;
        RECT 1.445 206.400 1767.255 207.720 ;
        RECT 4.400 205.000 1767.255 206.400 ;
        RECT 1.445 203.000 1767.255 205.000 ;
        RECT 4.400 201.600 1767.255 203.000 ;
        RECT 1.445 200.280 1767.255 201.600 ;
        RECT 1.445 198.920 1762.995 200.280 ;
        RECT 4.400 198.880 1762.995 198.920 ;
        RECT 4.400 197.520 1767.255 198.880 ;
        RECT 1.445 195.520 1767.255 197.520 ;
        RECT 4.400 194.120 1767.255 195.520 ;
        RECT 1.445 192.120 1767.255 194.120 ;
        RECT 4.400 191.440 1767.255 192.120 ;
        RECT 4.400 190.720 1762.995 191.440 ;
        RECT 1.445 190.040 1762.995 190.720 ;
        RECT 1.445 188.720 1767.255 190.040 ;
        RECT 4.400 187.320 1767.255 188.720 ;
        RECT 1.445 185.320 1767.255 187.320 ;
        RECT 4.400 183.920 1767.255 185.320 ;
        RECT 1.445 182.600 1767.255 183.920 ;
        RECT 1.445 181.920 1762.995 182.600 ;
        RECT 4.400 181.200 1762.995 181.920 ;
        RECT 4.400 180.520 1767.255 181.200 ;
        RECT 1.445 177.840 1767.255 180.520 ;
        RECT 4.400 176.440 1767.255 177.840 ;
        RECT 1.445 174.440 1767.255 176.440 ;
        RECT 4.400 173.760 1767.255 174.440 ;
        RECT 4.400 173.040 1762.995 173.760 ;
        RECT 1.445 172.360 1762.995 173.040 ;
        RECT 1.445 171.040 1767.255 172.360 ;
        RECT 4.400 169.640 1767.255 171.040 ;
        RECT 1.445 167.640 1767.255 169.640 ;
        RECT 4.400 166.240 1767.255 167.640 ;
        RECT 1.445 164.920 1767.255 166.240 ;
        RECT 1.445 164.240 1762.995 164.920 ;
        RECT 4.400 163.520 1762.995 164.240 ;
        RECT 4.400 162.840 1767.255 163.520 ;
        RECT 1.445 160.840 1767.255 162.840 ;
        RECT 4.400 159.440 1767.255 160.840 ;
        RECT 1.445 156.760 1767.255 159.440 ;
        RECT 4.400 156.080 1767.255 156.760 ;
        RECT 4.400 155.360 1762.995 156.080 ;
        RECT 1.445 154.680 1762.995 155.360 ;
        RECT 1.445 153.360 1767.255 154.680 ;
        RECT 4.400 151.960 1767.255 153.360 ;
        RECT 1.445 149.960 1767.255 151.960 ;
        RECT 4.400 148.560 1767.255 149.960 ;
        RECT 1.445 147.240 1767.255 148.560 ;
        RECT 1.445 146.560 1762.995 147.240 ;
        RECT 4.400 145.840 1762.995 146.560 ;
        RECT 4.400 145.160 1767.255 145.840 ;
        RECT 1.445 143.160 1767.255 145.160 ;
        RECT 4.400 141.760 1767.255 143.160 ;
        RECT 1.445 139.080 1767.255 141.760 ;
        RECT 4.400 138.400 1767.255 139.080 ;
        RECT 4.400 137.680 1762.995 138.400 ;
        RECT 1.445 137.000 1762.995 137.680 ;
        RECT 1.445 135.680 1767.255 137.000 ;
        RECT 4.400 134.280 1767.255 135.680 ;
        RECT 1.445 132.280 1767.255 134.280 ;
        RECT 4.400 130.880 1767.255 132.280 ;
        RECT 1.445 129.560 1767.255 130.880 ;
        RECT 1.445 128.880 1762.995 129.560 ;
        RECT 4.400 128.160 1762.995 128.880 ;
        RECT 4.400 127.480 1767.255 128.160 ;
        RECT 1.445 125.480 1767.255 127.480 ;
        RECT 4.400 124.080 1767.255 125.480 ;
        RECT 1.445 122.080 1767.255 124.080 ;
        RECT 4.400 120.680 1767.255 122.080 ;
        RECT 1.445 120.040 1767.255 120.680 ;
        RECT 1.445 118.640 1762.995 120.040 ;
        RECT 1.445 118.000 1767.255 118.640 ;
        RECT 4.400 116.600 1767.255 118.000 ;
        RECT 1.445 114.600 1767.255 116.600 ;
        RECT 4.400 113.200 1767.255 114.600 ;
        RECT 1.445 111.200 1767.255 113.200 ;
        RECT 4.400 109.800 1762.995 111.200 ;
        RECT 1.445 107.800 1767.255 109.800 ;
        RECT 4.400 106.400 1767.255 107.800 ;
        RECT 1.445 104.400 1767.255 106.400 ;
        RECT 4.400 103.000 1767.255 104.400 ;
        RECT 1.445 102.360 1767.255 103.000 ;
        RECT 1.445 100.960 1762.995 102.360 ;
        RECT 1.445 100.320 1767.255 100.960 ;
        RECT 4.400 98.920 1767.255 100.320 ;
        RECT 1.445 96.920 1767.255 98.920 ;
        RECT 4.400 95.520 1767.255 96.920 ;
        RECT 1.445 93.520 1767.255 95.520 ;
        RECT 4.400 92.120 1762.995 93.520 ;
        RECT 1.445 90.120 1767.255 92.120 ;
        RECT 4.400 88.720 1767.255 90.120 ;
        RECT 1.445 86.720 1767.255 88.720 ;
        RECT 4.400 85.320 1767.255 86.720 ;
        RECT 1.445 84.680 1767.255 85.320 ;
        RECT 1.445 83.320 1762.995 84.680 ;
        RECT 4.400 83.280 1762.995 83.320 ;
        RECT 4.400 81.920 1767.255 83.280 ;
        RECT 1.445 79.240 1767.255 81.920 ;
        RECT 4.400 77.840 1767.255 79.240 ;
        RECT 1.445 75.840 1767.255 77.840 ;
        RECT 4.400 74.440 1762.995 75.840 ;
        RECT 1.445 72.440 1767.255 74.440 ;
        RECT 4.400 71.040 1767.255 72.440 ;
        RECT 1.445 69.040 1767.255 71.040 ;
        RECT 4.400 67.640 1767.255 69.040 ;
        RECT 1.445 67.000 1767.255 67.640 ;
        RECT 1.445 65.640 1762.995 67.000 ;
        RECT 4.400 65.600 1762.995 65.640 ;
        RECT 4.400 64.240 1767.255 65.600 ;
        RECT 1.445 62.240 1767.255 64.240 ;
        RECT 4.400 60.840 1767.255 62.240 ;
        RECT 1.445 58.160 1767.255 60.840 ;
        RECT 4.400 56.760 1762.995 58.160 ;
        RECT 1.445 54.760 1767.255 56.760 ;
        RECT 4.400 53.360 1767.255 54.760 ;
        RECT 1.445 51.360 1767.255 53.360 ;
        RECT 4.400 49.960 1767.255 51.360 ;
        RECT 1.445 49.320 1767.255 49.960 ;
        RECT 1.445 47.960 1762.995 49.320 ;
        RECT 4.400 47.920 1762.995 47.960 ;
        RECT 4.400 46.560 1767.255 47.920 ;
        RECT 1.445 44.560 1767.255 46.560 ;
        RECT 4.400 43.160 1767.255 44.560 ;
        RECT 1.445 40.480 1767.255 43.160 ;
        RECT 4.400 39.080 1762.995 40.480 ;
        RECT 1.445 37.080 1767.255 39.080 ;
        RECT 4.400 35.680 1767.255 37.080 ;
        RECT 1.445 33.680 1767.255 35.680 ;
        RECT 4.400 32.280 1767.255 33.680 ;
        RECT 1.445 31.640 1767.255 32.280 ;
        RECT 1.445 30.280 1762.995 31.640 ;
        RECT 4.400 30.240 1762.995 30.280 ;
        RECT 4.400 28.880 1767.255 30.240 ;
        RECT 1.445 26.880 1767.255 28.880 ;
        RECT 4.400 25.480 1767.255 26.880 ;
        RECT 1.445 23.480 1767.255 25.480 ;
        RECT 4.400 22.800 1767.255 23.480 ;
        RECT 4.400 22.080 1762.995 22.800 ;
        RECT 1.445 21.400 1762.995 22.080 ;
        RECT 1.445 19.400 1767.255 21.400 ;
        RECT 4.400 18.000 1767.255 19.400 ;
        RECT 1.445 16.000 1767.255 18.000 ;
        RECT 4.400 14.600 1767.255 16.000 ;
        RECT 1.445 13.960 1767.255 14.600 ;
        RECT 1.445 12.600 1762.995 13.960 ;
        RECT 4.400 12.560 1762.995 12.600 ;
        RECT 4.400 11.200 1767.255 12.560 ;
        RECT 1.445 9.200 1767.255 11.200 ;
        RECT 4.400 7.800 1767.255 9.200 ;
        RECT 1.445 5.800 1767.255 7.800 ;
        RECT 4.400 5.120 1767.255 5.800 ;
        RECT 4.400 4.400 1762.995 5.120 ;
        RECT 1.445 3.720 1762.995 4.400 ;
        RECT 1.445 2.400 1767.255 3.720 ;
        RECT 4.400 1.535 1767.255 2.400 ;
      LAYER met4 ;
        RECT 3.975 1765.920 1765.185 1767.825 ;
        RECT 3.975 10.240 20.640 1765.920 ;
        RECT 23.040 10.240 97.440 1765.920 ;
        RECT 99.840 10.240 174.240 1765.920 ;
        RECT 176.640 10.240 251.040 1765.920 ;
        RECT 253.440 10.240 327.840 1765.920 ;
        RECT 330.240 10.240 404.640 1765.920 ;
        RECT 407.040 10.240 481.440 1765.920 ;
        RECT 483.840 10.240 558.240 1765.920 ;
        RECT 560.640 10.240 635.040 1765.920 ;
        RECT 637.440 10.240 711.840 1765.920 ;
        RECT 714.240 10.240 788.640 1765.920 ;
        RECT 791.040 10.240 865.440 1765.920 ;
        RECT 867.840 10.240 942.240 1765.920 ;
        RECT 944.640 10.240 1019.040 1765.920 ;
        RECT 1021.440 10.240 1095.840 1765.920 ;
        RECT 1098.240 10.240 1172.640 1765.920 ;
        RECT 1175.040 10.240 1249.440 1765.920 ;
        RECT 1251.840 10.240 1326.240 1765.920 ;
        RECT 1328.640 10.240 1403.040 1765.920 ;
        RECT 1405.440 10.240 1479.840 1765.920 ;
        RECT 1482.240 10.240 1556.640 1765.920 ;
        RECT 1559.040 10.240 1633.440 1765.920 ;
        RECT 1635.840 10.240 1710.240 1765.920 ;
        RECT 1712.640 10.240 1765.185 1765.920 ;
        RECT 3.975 9.015 1765.185 10.240 ;
  END
END Marmot
END LIBRARY

