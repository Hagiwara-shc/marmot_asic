magic
tech sky130A
magscale 1 2
timestamp 1647856827
<< obsli1 >>
rect 1104 2159 350152 350897
<< obsm1 >>
rect 290 1232 350966 353456
<< metal2 >>
rect 386 352669 442 353469
rect 1214 352669 1270 353469
rect 2134 352669 2190 353469
rect 3054 352669 3110 353469
rect 3882 352669 3938 353469
rect 4802 352669 4858 353469
rect 5722 352669 5778 353469
rect 6642 352669 6698 353469
rect 7470 352669 7526 353469
rect 8390 352669 8446 353469
rect 9310 352669 9366 353469
rect 10138 352669 10194 353469
rect 11058 352669 11114 353469
rect 11978 352669 12034 353469
rect 12898 352669 12954 353469
rect 13726 352669 13782 353469
rect 14646 352669 14702 353469
rect 15566 352669 15622 353469
rect 16394 352669 16450 353469
rect 17314 352669 17370 353469
rect 18234 352669 18290 353469
rect 19154 352669 19210 353469
rect 19982 352669 20038 353469
rect 20902 352669 20958 353469
rect 21822 352669 21878 353469
rect 22650 352669 22706 353469
rect 23570 352669 23626 353469
rect 24490 352669 24546 353469
rect 25410 352669 25466 353469
rect 26238 352669 26294 353469
rect 27158 352669 27214 353469
rect 28078 352669 28134 353469
rect 28906 352669 28962 353469
rect 29826 352669 29882 353469
rect 30746 352669 30802 353469
rect 31666 352669 31722 353469
rect 32494 352669 32550 353469
rect 33414 352669 33470 353469
rect 34334 352669 34390 353469
rect 35162 352669 35218 353469
rect 36082 352669 36138 353469
rect 37002 352669 37058 353469
rect 37922 352669 37978 353469
rect 38750 352669 38806 353469
rect 39670 352669 39726 353469
rect 40590 352669 40646 353469
rect 41510 352669 41566 353469
rect 42338 352669 42394 353469
rect 43258 352669 43314 353469
rect 44178 352669 44234 353469
rect 45006 352669 45062 353469
rect 45926 352669 45982 353469
rect 46846 352669 46902 353469
rect 47766 352669 47822 353469
rect 48594 352669 48650 353469
rect 49514 352669 49570 353469
rect 50434 352669 50490 353469
rect 51262 352669 51318 353469
rect 52182 352669 52238 353469
rect 53102 352669 53158 353469
rect 54022 352669 54078 353469
rect 54850 352669 54906 353469
rect 55770 352669 55826 353469
rect 56690 352669 56746 353469
rect 57518 352669 57574 353469
rect 58438 352669 58494 353469
rect 59358 352669 59414 353469
rect 60278 352669 60334 353469
rect 61106 352669 61162 353469
rect 62026 352669 62082 353469
rect 62946 352669 63002 353469
rect 63774 352669 63830 353469
rect 64694 352669 64750 353469
rect 65614 352669 65670 353469
rect 66534 352669 66590 353469
rect 67362 352669 67418 353469
rect 68282 352669 68338 353469
rect 69202 352669 69258 353469
rect 70030 352669 70086 353469
rect 70950 352669 71006 353469
rect 71870 352669 71926 353469
rect 72790 352669 72846 353469
rect 73618 352669 73674 353469
rect 74538 352669 74594 353469
rect 75458 352669 75514 353469
rect 76286 352669 76342 353469
rect 77206 352669 77262 353469
rect 78126 352669 78182 353469
rect 79046 352669 79102 353469
rect 79874 352669 79930 353469
rect 80794 352669 80850 353469
rect 81714 352669 81770 353469
rect 82634 352669 82690 353469
rect 83462 352669 83518 353469
rect 84382 352669 84438 353469
rect 85302 352669 85358 353469
rect 86130 352669 86186 353469
rect 87050 352669 87106 353469
rect 87970 352669 88026 353469
rect 88890 352669 88946 353469
rect 89718 352669 89774 353469
rect 90638 352669 90694 353469
rect 91558 352669 91614 353469
rect 92386 352669 92442 353469
rect 93306 352669 93362 353469
rect 94226 352669 94282 353469
rect 95146 352669 95202 353469
rect 95974 352669 96030 353469
rect 96894 352669 96950 353469
rect 97814 352669 97870 353469
rect 98642 352669 98698 353469
rect 99562 352669 99618 353469
rect 100482 352669 100538 353469
rect 101402 352669 101458 353469
rect 102230 352669 102286 353469
rect 103150 352669 103206 353469
rect 104070 352669 104126 353469
rect 104898 352669 104954 353469
rect 105818 352669 105874 353469
rect 106738 352669 106794 353469
rect 107658 352669 107714 353469
rect 108486 352669 108542 353469
rect 109406 352669 109462 353469
rect 110326 352669 110382 353469
rect 111154 352669 111210 353469
rect 112074 352669 112130 353469
rect 112994 352669 113050 353469
rect 113914 352669 113970 353469
rect 114742 352669 114798 353469
rect 115662 352669 115718 353469
rect 116582 352669 116638 353469
rect 117502 352669 117558 353469
rect 118330 352669 118386 353469
rect 119250 352669 119306 353469
rect 120170 352669 120226 353469
rect 120998 352669 121054 353469
rect 121918 352669 121974 353469
rect 122838 352669 122894 353469
rect 123758 352669 123814 353469
rect 124586 352669 124642 353469
rect 125506 352669 125562 353469
rect 126426 352669 126482 353469
rect 127254 352669 127310 353469
rect 128174 352669 128230 353469
rect 129094 352669 129150 353469
rect 130014 352669 130070 353469
rect 130842 352669 130898 353469
rect 131762 352669 131818 353469
rect 132682 352669 132738 353469
rect 133510 352669 133566 353469
rect 134430 352669 134486 353469
rect 135350 352669 135406 353469
rect 136270 352669 136326 353469
rect 137098 352669 137154 353469
rect 138018 352669 138074 353469
rect 138938 352669 138994 353469
rect 139766 352669 139822 353469
rect 140686 352669 140742 353469
rect 141606 352669 141662 353469
rect 142526 352669 142582 353469
rect 143354 352669 143410 353469
rect 144274 352669 144330 353469
rect 145194 352669 145250 353469
rect 146022 352669 146078 353469
rect 146942 352669 146998 353469
rect 147862 352669 147918 353469
rect 148782 352669 148838 353469
rect 149610 352669 149666 353469
rect 150530 352669 150586 353469
rect 151450 352669 151506 353469
rect 152278 352669 152334 353469
rect 153198 352669 153254 353469
rect 154118 352669 154174 353469
rect 155038 352669 155094 353469
rect 155866 352669 155922 353469
rect 156786 352669 156842 353469
rect 157706 352669 157762 353469
rect 158626 352669 158682 353469
rect 159454 352669 159510 353469
rect 160374 352669 160430 353469
rect 161294 352669 161350 353469
rect 162122 352669 162178 353469
rect 163042 352669 163098 353469
rect 163962 352669 164018 353469
rect 164882 352669 164938 353469
rect 165710 352669 165766 353469
rect 166630 352669 166686 353469
rect 167550 352669 167606 353469
rect 168378 352669 168434 353469
rect 169298 352669 169354 353469
rect 170218 352669 170274 353469
rect 171138 352669 171194 353469
rect 171966 352669 172022 353469
rect 172886 352669 172942 353469
rect 173806 352669 173862 353469
rect 174634 352669 174690 353469
rect 175554 352669 175610 353469
rect 176474 352669 176530 353469
rect 177394 352669 177450 353469
rect 178222 352669 178278 353469
rect 179142 352669 179198 353469
rect 180062 352669 180118 353469
rect 180890 352669 180946 353469
rect 181810 352669 181866 353469
rect 182730 352669 182786 353469
rect 183650 352669 183706 353469
rect 184478 352669 184534 353469
rect 185398 352669 185454 353469
rect 186318 352669 186374 353469
rect 187146 352669 187202 353469
rect 188066 352669 188122 353469
rect 188986 352669 189042 353469
rect 189906 352669 189962 353469
rect 190734 352669 190790 353469
rect 191654 352669 191710 353469
rect 192574 352669 192630 353469
rect 193402 352669 193458 353469
rect 194322 352669 194378 353469
rect 195242 352669 195298 353469
rect 196162 352669 196218 353469
rect 196990 352669 197046 353469
rect 197910 352669 197966 353469
rect 198830 352669 198886 353469
rect 199750 352669 199806 353469
rect 200578 352669 200634 353469
rect 201498 352669 201554 353469
rect 202418 352669 202474 353469
rect 203246 352669 203302 353469
rect 204166 352669 204222 353469
rect 205086 352669 205142 353469
rect 206006 352669 206062 353469
rect 206834 352669 206890 353469
rect 207754 352669 207810 353469
rect 208674 352669 208730 353469
rect 209502 352669 209558 353469
rect 210422 352669 210478 353469
rect 211342 352669 211398 353469
rect 212262 352669 212318 353469
rect 213090 352669 213146 353469
rect 214010 352669 214066 353469
rect 214930 352669 214986 353469
rect 215758 352669 215814 353469
rect 216678 352669 216734 353469
rect 217598 352669 217654 353469
rect 218518 352669 218574 353469
rect 219346 352669 219402 353469
rect 220266 352669 220322 353469
rect 221186 352669 221242 353469
rect 222014 352669 222070 353469
rect 222934 352669 222990 353469
rect 223854 352669 223910 353469
rect 224774 352669 224830 353469
rect 225602 352669 225658 353469
rect 226522 352669 226578 353469
rect 227442 352669 227498 353469
rect 228270 352669 228326 353469
rect 229190 352669 229246 353469
rect 230110 352669 230166 353469
rect 231030 352669 231086 353469
rect 231858 352669 231914 353469
rect 232778 352669 232834 353469
rect 233698 352669 233754 353469
rect 234618 352669 234674 353469
rect 235446 352669 235502 353469
rect 236366 352669 236422 353469
rect 237286 352669 237342 353469
rect 238114 352669 238170 353469
rect 239034 352669 239090 353469
rect 239954 352669 240010 353469
rect 240874 352669 240930 353469
rect 241702 352669 241758 353469
rect 242622 352669 242678 353469
rect 243542 352669 243598 353469
rect 244370 352669 244426 353469
rect 245290 352669 245346 353469
rect 246210 352669 246266 353469
rect 247130 352669 247186 353469
rect 247958 352669 248014 353469
rect 248878 352669 248934 353469
rect 249798 352669 249854 353469
rect 250626 352669 250682 353469
rect 251546 352669 251602 353469
rect 252466 352669 252522 353469
rect 253386 352669 253442 353469
rect 254214 352669 254270 353469
rect 255134 352669 255190 353469
rect 256054 352669 256110 353469
rect 256882 352669 256938 353469
rect 257802 352669 257858 353469
rect 258722 352669 258778 353469
rect 259642 352669 259698 353469
rect 260470 352669 260526 353469
rect 261390 352669 261446 353469
rect 262310 352669 262366 353469
rect 263138 352669 263194 353469
rect 264058 352669 264114 353469
rect 264978 352669 265034 353469
rect 265898 352669 265954 353469
rect 266726 352669 266782 353469
rect 267646 352669 267702 353469
rect 268566 352669 268622 353469
rect 269394 352669 269450 353469
rect 270314 352669 270370 353469
rect 271234 352669 271290 353469
rect 272154 352669 272210 353469
rect 272982 352669 273038 353469
rect 273902 352669 273958 353469
rect 274822 352669 274878 353469
rect 275742 352669 275798 353469
rect 276570 352669 276626 353469
rect 277490 352669 277546 353469
rect 278410 352669 278466 353469
rect 279238 352669 279294 353469
rect 280158 352669 280214 353469
rect 281078 352669 281134 353469
rect 281998 352669 282054 353469
rect 282826 352669 282882 353469
rect 283746 352669 283802 353469
rect 284666 352669 284722 353469
rect 285494 352669 285550 353469
rect 286414 352669 286470 353469
rect 287334 352669 287390 353469
rect 288254 352669 288310 353469
rect 289082 352669 289138 353469
rect 290002 352669 290058 353469
rect 290922 352669 290978 353469
rect 291750 352669 291806 353469
rect 292670 352669 292726 353469
rect 293590 352669 293646 353469
rect 294510 352669 294566 353469
rect 295338 352669 295394 353469
rect 296258 352669 296314 353469
rect 297178 352669 297234 353469
rect 298006 352669 298062 353469
rect 298926 352669 298982 353469
rect 299846 352669 299902 353469
rect 300766 352669 300822 353469
rect 301594 352669 301650 353469
rect 302514 352669 302570 353469
rect 303434 352669 303490 353469
rect 304262 352669 304318 353469
rect 305182 352669 305238 353469
rect 306102 352669 306158 353469
rect 307022 352669 307078 353469
rect 307850 352669 307906 353469
rect 308770 352669 308826 353469
rect 309690 352669 309746 353469
rect 310518 352669 310574 353469
rect 311438 352669 311494 353469
rect 312358 352669 312414 353469
rect 313278 352669 313334 353469
rect 314106 352669 314162 353469
rect 315026 352669 315082 353469
rect 315946 352669 316002 353469
rect 316866 352669 316922 353469
rect 317694 352669 317750 353469
rect 318614 352669 318670 353469
rect 319534 352669 319590 353469
rect 320362 352669 320418 353469
rect 321282 352669 321338 353469
rect 322202 352669 322258 353469
rect 323122 352669 323178 353469
rect 323950 352669 324006 353469
rect 324870 352669 324926 353469
rect 325790 352669 325846 353469
rect 326618 352669 326674 353469
rect 327538 352669 327594 353469
rect 328458 352669 328514 353469
rect 329378 352669 329434 353469
rect 330206 352669 330262 353469
rect 331126 352669 331182 353469
rect 332046 352669 332102 353469
rect 332874 352669 332930 353469
rect 333794 352669 333850 353469
rect 334714 352669 334770 353469
rect 335634 352669 335690 353469
rect 336462 352669 336518 353469
rect 337382 352669 337438 353469
rect 338302 352669 338358 353469
rect 339130 352669 339186 353469
rect 340050 352669 340106 353469
rect 340970 352669 341026 353469
rect 341890 352669 341946 353469
rect 342718 352669 342774 353469
rect 343638 352669 343694 353469
rect 344558 352669 344614 353469
rect 345386 352669 345442 353469
rect 346306 352669 346362 353469
rect 347226 352669 347282 353469
rect 348146 352669 348202 353469
rect 348974 352669 349030 353469
rect 349894 352669 349950 353469
rect 350814 352669 350870 353469
rect 294 0 350 800
rect 938 0 994 800
rect 1674 0 1730 800
rect 2410 0 2466 800
rect 3054 0 3110 800
rect 3790 0 3846 800
rect 4526 0 4582 800
rect 5262 0 5318 800
rect 5906 0 5962 800
rect 6642 0 6698 800
rect 7378 0 7434 800
rect 8114 0 8170 800
rect 8758 0 8814 800
rect 9494 0 9550 800
rect 10230 0 10286 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12346 0 12402 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 14462 0 14518 800
rect 15198 0 15254 800
rect 15934 0 15990 800
rect 16670 0 16726 800
rect 17314 0 17370 800
rect 18050 0 18106 800
rect 18786 0 18842 800
rect 19522 0 19578 800
rect 20166 0 20222 800
rect 20902 0 20958 800
rect 21638 0 21694 800
rect 22374 0 22430 800
rect 23018 0 23074 800
rect 23754 0 23810 800
rect 24490 0 24546 800
rect 25226 0 25282 800
rect 25870 0 25926 800
rect 26606 0 26662 800
rect 27342 0 27398 800
rect 28078 0 28134 800
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30194 0 30250 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32310 0 32366 800
rect 33046 0 33102 800
rect 33782 0 33838 800
rect 34426 0 34482 800
rect 35162 0 35218 800
rect 35898 0 35954 800
rect 36634 0 36690 800
rect 37278 0 37334 800
rect 38014 0 38070 800
rect 38750 0 38806 800
rect 39486 0 39542 800
rect 40130 0 40186 800
rect 40866 0 40922 800
rect 41602 0 41658 800
rect 42338 0 42394 800
rect 42982 0 43038 800
rect 43718 0 43774 800
rect 44454 0 44510 800
rect 45190 0 45246 800
rect 45834 0 45890 800
rect 46570 0 46626 800
rect 47306 0 47362 800
rect 48042 0 48098 800
rect 48686 0 48742 800
rect 49422 0 49478 800
rect 50158 0 50214 800
rect 50802 0 50858 800
rect 51538 0 51594 800
rect 52274 0 52330 800
rect 53010 0 53066 800
rect 53654 0 53710 800
rect 54390 0 54446 800
rect 55126 0 55182 800
rect 55862 0 55918 800
rect 56506 0 56562 800
rect 57242 0 57298 800
rect 57978 0 58034 800
rect 58714 0 58770 800
rect 59358 0 59414 800
rect 60094 0 60150 800
rect 60830 0 60886 800
rect 61566 0 61622 800
rect 62210 0 62266 800
rect 62946 0 63002 800
rect 63682 0 63738 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65798 0 65854 800
rect 66534 0 66590 800
rect 67270 0 67326 800
rect 67914 0 67970 800
rect 68650 0 68706 800
rect 69386 0 69442 800
rect 70122 0 70178 800
rect 70766 0 70822 800
rect 71502 0 71558 800
rect 72238 0 72294 800
rect 72974 0 73030 800
rect 73618 0 73674 800
rect 74354 0 74410 800
rect 75090 0 75146 800
rect 75826 0 75882 800
rect 76470 0 76526 800
rect 77206 0 77262 800
rect 77942 0 77998 800
rect 78678 0 78734 800
rect 79322 0 79378 800
rect 80058 0 80114 800
rect 80794 0 80850 800
rect 81530 0 81586 800
rect 82174 0 82230 800
rect 82910 0 82966 800
rect 83646 0 83702 800
rect 84382 0 84438 800
rect 85026 0 85082 800
rect 85762 0 85818 800
rect 86498 0 86554 800
rect 87234 0 87290 800
rect 87878 0 87934 800
rect 88614 0 88670 800
rect 89350 0 89406 800
rect 90086 0 90142 800
rect 90730 0 90786 800
rect 91466 0 91522 800
rect 92202 0 92258 800
rect 92938 0 92994 800
rect 93582 0 93638 800
rect 94318 0 94374 800
rect 95054 0 95110 800
rect 95790 0 95846 800
rect 96434 0 96490 800
rect 97170 0 97226 800
rect 97906 0 97962 800
rect 98642 0 98698 800
rect 99286 0 99342 800
rect 100022 0 100078 800
rect 100758 0 100814 800
rect 101402 0 101458 800
rect 102138 0 102194 800
rect 102874 0 102930 800
rect 103610 0 103666 800
rect 104254 0 104310 800
rect 104990 0 105046 800
rect 105726 0 105782 800
rect 106462 0 106518 800
rect 107106 0 107162 800
rect 107842 0 107898 800
rect 108578 0 108634 800
rect 109314 0 109370 800
rect 109958 0 110014 800
rect 110694 0 110750 800
rect 111430 0 111486 800
rect 112166 0 112222 800
rect 112810 0 112866 800
rect 113546 0 113602 800
rect 114282 0 114338 800
rect 115018 0 115074 800
rect 115662 0 115718 800
rect 116398 0 116454 800
rect 117134 0 117190 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119250 0 119306 800
rect 119986 0 120042 800
rect 120722 0 120778 800
rect 121366 0 121422 800
rect 122102 0 122158 800
rect 122838 0 122894 800
rect 123574 0 123630 800
rect 124218 0 124274 800
rect 124954 0 125010 800
rect 125690 0 125746 800
rect 126426 0 126482 800
rect 127070 0 127126 800
rect 127806 0 127862 800
rect 128542 0 128598 800
rect 129278 0 129334 800
rect 129922 0 129978 800
rect 130658 0 130714 800
rect 131394 0 131450 800
rect 132130 0 132186 800
rect 132774 0 132830 800
rect 133510 0 133566 800
rect 134246 0 134302 800
rect 134982 0 135038 800
rect 135626 0 135682 800
rect 136362 0 136418 800
rect 137098 0 137154 800
rect 137834 0 137890 800
rect 138478 0 138534 800
rect 139214 0 139270 800
rect 139950 0 140006 800
rect 140686 0 140742 800
rect 141330 0 141386 800
rect 142066 0 142122 800
rect 142802 0 142858 800
rect 143538 0 143594 800
rect 144182 0 144238 800
rect 144918 0 144974 800
rect 145654 0 145710 800
rect 146390 0 146446 800
rect 147034 0 147090 800
rect 147770 0 147826 800
rect 148506 0 148562 800
rect 149242 0 149298 800
rect 149886 0 149942 800
rect 150622 0 150678 800
rect 151358 0 151414 800
rect 152002 0 152058 800
rect 152738 0 152794 800
rect 153474 0 153530 800
rect 154210 0 154266 800
rect 154854 0 154910 800
rect 155590 0 155646 800
rect 156326 0 156382 800
rect 157062 0 157118 800
rect 157706 0 157762 800
rect 158442 0 158498 800
rect 159178 0 159234 800
rect 159914 0 159970 800
rect 160558 0 160614 800
rect 161294 0 161350 800
rect 162030 0 162086 800
rect 162766 0 162822 800
rect 163410 0 163466 800
rect 164146 0 164202 800
rect 164882 0 164938 800
rect 165618 0 165674 800
rect 166262 0 166318 800
rect 166998 0 167054 800
rect 167734 0 167790 800
rect 168470 0 168526 800
rect 169114 0 169170 800
rect 169850 0 169906 800
rect 170586 0 170642 800
rect 171322 0 171378 800
rect 171966 0 172022 800
rect 172702 0 172758 800
rect 173438 0 173494 800
rect 174174 0 174230 800
rect 174818 0 174874 800
rect 175554 0 175610 800
rect 176290 0 176346 800
rect 177026 0 177082 800
rect 177670 0 177726 800
rect 178406 0 178462 800
rect 179142 0 179198 800
rect 179878 0 179934 800
rect 180522 0 180578 800
rect 181258 0 181314 800
rect 181994 0 182050 800
rect 182730 0 182786 800
rect 183374 0 183430 800
rect 184110 0 184166 800
rect 184846 0 184902 800
rect 185582 0 185638 800
rect 186226 0 186282 800
rect 186962 0 187018 800
rect 187698 0 187754 800
rect 188434 0 188490 800
rect 189078 0 189134 800
rect 189814 0 189870 800
rect 190550 0 190606 800
rect 191286 0 191342 800
rect 191930 0 191986 800
rect 192666 0 192722 800
rect 193402 0 193458 800
rect 194138 0 194194 800
rect 194782 0 194838 800
rect 195518 0 195574 800
rect 196254 0 196310 800
rect 196990 0 197046 800
rect 197634 0 197690 800
rect 198370 0 198426 800
rect 199106 0 199162 800
rect 199842 0 199898 800
rect 200486 0 200542 800
rect 201222 0 201278 800
rect 201958 0 202014 800
rect 202602 0 202658 800
rect 203338 0 203394 800
rect 204074 0 204130 800
rect 204810 0 204866 800
rect 205454 0 205510 800
rect 206190 0 206246 800
rect 206926 0 206982 800
rect 207662 0 207718 800
rect 208306 0 208362 800
rect 209042 0 209098 800
rect 209778 0 209834 800
rect 210514 0 210570 800
rect 211158 0 211214 800
rect 211894 0 211950 800
rect 212630 0 212686 800
rect 213366 0 213422 800
rect 214010 0 214066 800
rect 214746 0 214802 800
rect 215482 0 215538 800
rect 216218 0 216274 800
rect 216862 0 216918 800
rect 217598 0 217654 800
rect 218334 0 218390 800
rect 219070 0 219126 800
rect 219714 0 219770 800
rect 220450 0 220506 800
rect 221186 0 221242 800
rect 221922 0 221978 800
rect 222566 0 222622 800
rect 223302 0 223358 800
rect 224038 0 224094 800
rect 224774 0 224830 800
rect 225418 0 225474 800
rect 226154 0 226210 800
rect 226890 0 226946 800
rect 227626 0 227682 800
rect 228270 0 228326 800
rect 229006 0 229062 800
rect 229742 0 229798 800
rect 230478 0 230534 800
rect 231122 0 231178 800
rect 231858 0 231914 800
rect 232594 0 232650 800
rect 233330 0 233386 800
rect 233974 0 234030 800
rect 234710 0 234766 800
rect 235446 0 235502 800
rect 236182 0 236238 800
rect 236826 0 236882 800
rect 237562 0 237618 800
rect 238298 0 238354 800
rect 239034 0 239090 800
rect 239678 0 239734 800
rect 240414 0 240470 800
rect 241150 0 241206 800
rect 241886 0 241942 800
rect 242530 0 242586 800
rect 243266 0 243322 800
rect 244002 0 244058 800
rect 244738 0 244794 800
rect 245382 0 245438 800
rect 246118 0 246174 800
rect 246854 0 246910 800
rect 247590 0 247646 800
rect 248234 0 248290 800
rect 248970 0 249026 800
rect 249706 0 249762 800
rect 250442 0 250498 800
rect 251086 0 251142 800
rect 251822 0 251878 800
rect 252558 0 252614 800
rect 253202 0 253258 800
rect 253938 0 253994 800
rect 254674 0 254730 800
rect 255410 0 255466 800
rect 256054 0 256110 800
rect 256790 0 256846 800
rect 257526 0 257582 800
rect 258262 0 258318 800
rect 258906 0 258962 800
rect 259642 0 259698 800
rect 260378 0 260434 800
rect 261114 0 261170 800
rect 261758 0 261814 800
rect 262494 0 262550 800
rect 263230 0 263286 800
rect 263966 0 264022 800
rect 264610 0 264666 800
rect 265346 0 265402 800
rect 266082 0 266138 800
rect 266818 0 266874 800
rect 267462 0 267518 800
rect 268198 0 268254 800
rect 268934 0 268990 800
rect 269670 0 269726 800
rect 270314 0 270370 800
rect 271050 0 271106 800
rect 271786 0 271842 800
rect 272522 0 272578 800
rect 273166 0 273222 800
rect 273902 0 273958 800
rect 274638 0 274694 800
rect 275374 0 275430 800
rect 276018 0 276074 800
rect 276754 0 276810 800
rect 277490 0 277546 800
rect 278226 0 278282 800
rect 278870 0 278926 800
rect 279606 0 279662 800
rect 280342 0 280398 800
rect 281078 0 281134 800
rect 281722 0 281778 800
rect 282458 0 282514 800
rect 283194 0 283250 800
rect 283930 0 283986 800
rect 284574 0 284630 800
rect 285310 0 285366 800
rect 286046 0 286102 800
rect 286782 0 286838 800
rect 287426 0 287482 800
rect 288162 0 288218 800
rect 288898 0 288954 800
rect 289634 0 289690 800
rect 290278 0 290334 800
rect 291014 0 291070 800
rect 291750 0 291806 800
rect 292486 0 292542 800
rect 293130 0 293186 800
rect 293866 0 293922 800
rect 294602 0 294658 800
rect 295338 0 295394 800
rect 295982 0 296038 800
rect 296718 0 296774 800
rect 297454 0 297510 800
rect 298190 0 298246 800
rect 298834 0 298890 800
rect 299570 0 299626 800
rect 300306 0 300362 800
rect 301042 0 301098 800
rect 301686 0 301742 800
rect 302422 0 302478 800
rect 303158 0 303214 800
rect 303802 0 303858 800
rect 304538 0 304594 800
rect 305274 0 305330 800
rect 306010 0 306066 800
rect 306654 0 306710 800
rect 307390 0 307446 800
rect 308126 0 308182 800
rect 308862 0 308918 800
rect 309506 0 309562 800
rect 310242 0 310298 800
rect 310978 0 311034 800
rect 311714 0 311770 800
rect 312358 0 312414 800
rect 313094 0 313150 800
rect 313830 0 313886 800
rect 314566 0 314622 800
rect 315210 0 315266 800
rect 315946 0 316002 800
rect 316682 0 316738 800
rect 317418 0 317474 800
rect 318062 0 318118 800
rect 318798 0 318854 800
rect 319534 0 319590 800
rect 320270 0 320326 800
rect 320914 0 320970 800
rect 321650 0 321706 800
rect 322386 0 322442 800
rect 323122 0 323178 800
rect 323766 0 323822 800
rect 324502 0 324558 800
rect 325238 0 325294 800
rect 325974 0 326030 800
rect 326618 0 326674 800
rect 327354 0 327410 800
rect 328090 0 328146 800
rect 328826 0 328882 800
rect 329470 0 329526 800
rect 330206 0 330262 800
rect 330942 0 330998 800
rect 331678 0 331734 800
rect 332322 0 332378 800
rect 333058 0 333114 800
rect 333794 0 333850 800
rect 334530 0 334586 800
rect 335174 0 335230 800
rect 335910 0 335966 800
rect 336646 0 336702 800
rect 337382 0 337438 800
rect 338026 0 338082 800
rect 338762 0 338818 800
rect 339498 0 339554 800
rect 340234 0 340290 800
rect 340878 0 340934 800
rect 341614 0 341670 800
rect 342350 0 342406 800
rect 343086 0 343142 800
rect 343730 0 343786 800
rect 344466 0 344522 800
rect 345202 0 345258 800
rect 345938 0 345994 800
rect 346582 0 346638 800
rect 347318 0 347374 800
rect 348054 0 348110 800
rect 348790 0 348846 800
rect 349434 0 349490 800
rect 350170 0 350226 800
rect 350906 0 350962 800
<< obsm2 >>
rect 296 352613 330 353462
rect 498 352613 1158 353462
rect 1326 352613 2078 353462
rect 2246 352613 2998 353462
rect 3166 352613 3826 353462
rect 3994 352613 4746 353462
rect 4914 352613 5666 353462
rect 5834 352613 6586 353462
rect 6754 352613 7414 353462
rect 7582 352613 8334 353462
rect 8502 352613 9254 353462
rect 9422 352613 10082 353462
rect 10250 352613 11002 353462
rect 11170 352613 11922 353462
rect 12090 352613 12842 353462
rect 13010 352613 13670 353462
rect 13838 352613 14590 353462
rect 14758 352613 15510 353462
rect 15678 352613 16338 353462
rect 16506 352613 17258 353462
rect 17426 352613 18178 353462
rect 18346 352613 19098 353462
rect 19266 352613 19926 353462
rect 20094 352613 20846 353462
rect 21014 352613 21766 353462
rect 21934 352613 22594 353462
rect 22762 352613 23514 353462
rect 23682 352613 24434 353462
rect 24602 352613 25354 353462
rect 25522 352613 26182 353462
rect 26350 352613 27102 353462
rect 27270 352613 28022 353462
rect 28190 352613 28850 353462
rect 29018 352613 29770 353462
rect 29938 352613 30690 353462
rect 30858 352613 31610 353462
rect 31778 352613 32438 353462
rect 32606 352613 33358 353462
rect 33526 352613 34278 353462
rect 34446 352613 35106 353462
rect 35274 352613 36026 353462
rect 36194 352613 36946 353462
rect 37114 352613 37866 353462
rect 38034 352613 38694 353462
rect 38862 352613 39614 353462
rect 39782 352613 40534 353462
rect 40702 352613 41454 353462
rect 41622 352613 42282 353462
rect 42450 352613 43202 353462
rect 43370 352613 44122 353462
rect 44290 352613 44950 353462
rect 45118 352613 45870 353462
rect 46038 352613 46790 353462
rect 46958 352613 47710 353462
rect 47878 352613 48538 353462
rect 48706 352613 49458 353462
rect 49626 352613 50378 353462
rect 50546 352613 51206 353462
rect 51374 352613 52126 353462
rect 52294 352613 53046 353462
rect 53214 352613 53966 353462
rect 54134 352613 54794 353462
rect 54962 352613 55714 353462
rect 55882 352613 56634 353462
rect 56802 352613 57462 353462
rect 57630 352613 58382 353462
rect 58550 352613 59302 353462
rect 59470 352613 60222 353462
rect 60390 352613 61050 353462
rect 61218 352613 61970 353462
rect 62138 352613 62890 353462
rect 63058 352613 63718 353462
rect 63886 352613 64638 353462
rect 64806 352613 65558 353462
rect 65726 352613 66478 353462
rect 66646 352613 67306 353462
rect 67474 352613 68226 353462
rect 68394 352613 69146 353462
rect 69314 352613 69974 353462
rect 70142 352613 70894 353462
rect 71062 352613 71814 353462
rect 71982 352613 72734 353462
rect 72902 352613 73562 353462
rect 73730 352613 74482 353462
rect 74650 352613 75402 353462
rect 75570 352613 76230 353462
rect 76398 352613 77150 353462
rect 77318 352613 78070 353462
rect 78238 352613 78990 353462
rect 79158 352613 79818 353462
rect 79986 352613 80738 353462
rect 80906 352613 81658 353462
rect 81826 352613 82578 353462
rect 82746 352613 83406 353462
rect 83574 352613 84326 353462
rect 84494 352613 85246 353462
rect 85414 352613 86074 353462
rect 86242 352613 86994 353462
rect 87162 352613 87914 353462
rect 88082 352613 88834 353462
rect 89002 352613 89662 353462
rect 89830 352613 90582 353462
rect 90750 352613 91502 353462
rect 91670 352613 92330 353462
rect 92498 352613 93250 353462
rect 93418 352613 94170 353462
rect 94338 352613 95090 353462
rect 95258 352613 95918 353462
rect 96086 352613 96838 353462
rect 97006 352613 97758 353462
rect 97926 352613 98586 353462
rect 98754 352613 99506 353462
rect 99674 352613 100426 353462
rect 100594 352613 101346 353462
rect 101514 352613 102174 353462
rect 102342 352613 103094 353462
rect 103262 352613 104014 353462
rect 104182 352613 104842 353462
rect 105010 352613 105762 353462
rect 105930 352613 106682 353462
rect 106850 352613 107602 353462
rect 107770 352613 108430 353462
rect 108598 352613 109350 353462
rect 109518 352613 110270 353462
rect 110438 352613 111098 353462
rect 111266 352613 112018 353462
rect 112186 352613 112938 353462
rect 113106 352613 113858 353462
rect 114026 352613 114686 353462
rect 114854 352613 115606 353462
rect 115774 352613 116526 353462
rect 116694 352613 117446 353462
rect 117614 352613 118274 353462
rect 118442 352613 119194 353462
rect 119362 352613 120114 353462
rect 120282 352613 120942 353462
rect 121110 352613 121862 353462
rect 122030 352613 122782 353462
rect 122950 352613 123702 353462
rect 123870 352613 124530 353462
rect 124698 352613 125450 353462
rect 125618 352613 126370 353462
rect 126538 352613 127198 353462
rect 127366 352613 128118 353462
rect 128286 352613 129038 353462
rect 129206 352613 129958 353462
rect 130126 352613 130786 353462
rect 130954 352613 131706 353462
rect 131874 352613 132626 353462
rect 132794 352613 133454 353462
rect 133622 352613 134374 353462
rect 134542 352613 135294 353462
rect 135462 352613 136214 353462
rect 136382 352613 137042 353462
rect 137210 352613 137962 353462
rect 138130 352613 138882 353462
rect 139050 352613 139710 353462
rect 139878 352613 140630 353462
rect 140798 352613 141550 353462
rect 141718 352613 142470 353462
rect 142638 352613 143298 353462
rect 143466 352613 144218 353462
rect 144386 352613 145138 353462
rect 145306 352613 145966 353462
rect 146134 352613 146886 353462
rect 147054 352613 147806 353462
rect 147974 352613 148726 353462
rect 148894 352613 149554 353462
rect 149722 352613 150474 353462
rect 150642 352613 151394 353462
rect 151562 352613 152222 353462
rect 152390 352613 153142 353462
rect 153310 352613 154062 353462
rect 154230 352613 154982 353462
rect 155150 352613 155810 353462
rect 155978 352613 156730 353462
rect 156898 352613 157650 353462
rect 157818 352613 158570 353462
rect 158738 352613 159398 353462
rect 159566 352613 160318 353462
rect 160486 352613 161238 353462
rect 161406 352613 162066 353462
rect 162234 352613 162986 353462
rect 163154 352613 163906 353462
rect 164074 352613 164826 353462
rect 164994 352613 165654 353462
rect 165822 352613 166574 353462
rect 166742 352613 167494 353462
rect 167662 352613 168322 353462
rect 168490 352613 169242 353462
rect 169410 352613 170162 353462
rect 170330 352613 171082 353462
rect 171250 352613 171910 353462
rect 172078 352613 172830 353462
rect 172998 352613 173750 353462
rect 173918 352613 174578 353462
rect 174746 352613 175498 353462
rect 175666 352613 176418 353462
rect 176586 352613 177338 353462
rect 177506 352613 178166 353462
rect 178334 352613 179086 353462
rect 179254 352613 180006 353462
rect 180174 352613 180834 353462
rect 181002 352613 181754 353462
rect 181922 352613 182674 353462
rect 182842 352613 183594 353462
rect 183762 352613 184422 353462
rect 184590 352613 185342 353462
rect 185510 352613 186262 353462
rect 186430 352613 187090 353462
rect 187258 352613 188010 353462
rect 188178 352613 188930 353462
rect 189098 352613 189850 353462
rect 190018 352613 190678 353462
rect 190846 352613 191598 353462
rect 191766 352613 192518 353462
rect 192686 352613 193346 353462
rect 193514 352613 194266 353462
rect 194434 352613 195186 353462
rect 195354 352613 196106 353462
rect 196274 352613 196934 353462
rect 197102 352613 197854 353462
rect 198022 352613 198774 353462
rect 198942 352613 199694 353462
rect 199862 352613 200522 353462
rect 200690 352613 201442 353462
rect 201610 352613 202362 353462
rect 202530 352613 203190 353462
rect 203358 352613 204110 353462
rect 204278 352613 205030 353462
rect 205198 352613 205950 353462
rect 206118 352613 206778 353462
rect 206946 352613 207698 353462
rect 207866 352613 208618 353462
rect 208786 352613 209446 353462
rect 209614 352613 210366 353462
rect 210534 352613 211286 353462
rect 211454 352613 212206 353462
rect 212374 352613 213034 353462
rect 213202 352613 213954 353462
rect 214122 352613 214874 353462
rect 215042 352613 215702 353462
rect 215870 352613 216622 353462
rect 216790 352613 217542 353462
rect 217710 352613 218462 353462
rect 218630 352613 219290 353462
rect 219458 352613 220210 353462
rect 220378 352613 221130 353462
rect 221298 352613 221958 353462
rect 222126 352613 222878 353462
rect 223046 352613 223798 353462
rect 223966 352613 224718 353462
rect 224886 352613 225546 353462
rect 225714 352613 226466 353462
rect 226634 352613 227386 353462
rect 227554 352613 228214 353462
rect 228382 352613 229134 353462
rect 229302 352613 230054 353462
rect 230222 352613 230974 353462
rect 231142 352613 231802 353462
rect 231970 352613 232722 353462
rect 232890 352613 233642 353462
rect 233810 352613 234562 353462
rect 234730 352613 235390 353462
rect 235558 352613 236310 353462
rect 236478 352613 237230 353462
rect 237398 352613 238058 353462
rect 238226 352613 238978 353462
rect 239146 352613 239898 353462
rect 240066 352613 240818 353462
rect 240986 352613 241646 353462
rect 241814 352613 242566 353462
rect 242734 352613 243486 353462
rect 243654 352613 244314 353462
rect 244482 352613 245234 353462
rect 245402 352613 246154 353462
rect 246322 352613 247074 353462
rect 247242 352613 247902 353462
rect 248070 352613 248822 353462
rect 248990 352613 249742 353462
rect 249910 352613 250570 353462
rect 250738 352613 251490 353462
rect 251658 352613 252410 353462
rect 252578 352613 253330 353462
rect 253498 352613 254158 353462
rect 254326 352613 255078 353462
rect 255246 352613 255998 353462
rect 256166 352613 256826 353462
rect 256994 352613 257746 353462
rect 257914 352613 258666 353462
rect 258834 352613 259586 353462
rect 259754 352613 260414 353462
rect 260582 352613 261334 353462
rect 261502 352613 262254 353462
rect 262422 352613 263082 353462
rect 263250 352613 264002 353462
rect 264170 352613 264922 353462
rect 265090 352613 265842 353462
rect 266010 352613 266670 353462
rect 266838 352613 267590 353462
rect 267758 352613 268510 353462
rect 268678 352613 269338 353462
rect 269506 352613 270258 353462
rect 270426 352613 271178 353462
rect 271346 352613 272098 353462
rect 272266 352613 272926 353462
rect 273094 352613 273846 353462
rect 274014 352613 274766 353462
rect 274934 352613 275686 353462
rect 275854 352613 276514 353462
rect 276682 352613 277434 353462
rect 277602 352613 278354 353462
rect 278522 352613 279182 353462
rect 279350 352613 280102 353462
rect 280270 352613 281022 353462
rect 281190 352613 281942 353462
rect 282110 352613 282770 353462
rect 282938 352613 283690 353462
rect 283858 352613 284610 353462
rect 284778 352613 285438 353462
rect 285606 352613 286358 353462
rect 286526 352613 287278 353462
rect 287446 352613 288198 353462
rect 288366 352613 289026 353462
rect 289194 352613 289946 353462
rect 290114 352613 290866 353462
rect 291034 352613 291694 353462
rect 291862 352613 292614 353462
rect 292782 352613 293534 353462
rect 293702 352613 294454 353462
rect 294622 352613 295282 353462
rect 295450 352613 296202 353462
rect 296370 352613 297122 353462
rect 297290 352613 297950 353462
rect 298118 352613 298870 353462
rect 299038 352613 299790 353462
rect 299958 352613 300710 353462
rect 300878 352613 301538 353462
rect 301706 352613 302458 353462
rect 302626 352613 303378 353462
rect 303546 352613 304206 353462
rect 304374 352613 305126 353462
rect 305294 352613 306046 353462
rect 306214 352613 306966 353462
rect 307134 352613 307794 353462
rect 307962 352613 308714 353462
rect 308882 352613 309634 353462
rect 309802 352613 310462 353462
rect 310630 352613 311382 353462
rect 311550 352613 312302 353462
rect 312470 352613 313222 353462
rect 313390 352613 314050 353462
rect 314218 352613 314970 353462
rect 315138 352613 315890 353462
rect 316058 352613 316810 353462
rect 316978 352613 317638 353462
rect 317806 352613 318558 353462
rect 318726 352613 319478 353462
rect 319646 352613 320306 353462
rect 320474 352613 321226 353462
rect 321394 352613 322146 353462
rect 322314 352613 323066 353462
rect 323234 352613 323894 353462
rect 324062 352613 324814 353462
rect 324982 352613 325734 353462
rect 325902 352613 326562 353462
rect 326730 352613 327482 353462
rect 327650 352613 328402 353462
rect 328570 352613 329322 353462
rect 329490 352613 330150 353462
rect 330318 352613 331070 353462
rect 331238 352613 331990 353462
rect 332158 352613 332818 353462
rect 332986 352613 333738 353462
rect 333906 352613 334658 353462
rect 334826 352613 335578 353462
rect 335746 352613 336406 353462
rect 336574 352613 337326 353462
rect 337494 352613 338246 353462
rect 338414 352613 339074 353462
rect 339242 352613 339994 353462
rect 340162 352613 340914 353462
rect 341082 352613 341834 353462
rect 342002 352613 342662 353462
rect 342830 352613 343582 353462
rect 343750 352613 344502 353462
rect 344670 352613 345330 353462
rect 345498 352613 346250 353462
rect 346418 352613 347170 353462
rect 347338 352613 348090 353462
rect 348258 352613 348918 353462
rect 349086 352613 349838 353462
rect 350006 352613 350758 353462
rect 350926 352613 350960 353462
rect 296 856 350960 352613
rect 406 734 882 856
rect 1050 734 1618 856
rect 1786 734 2354 856
rect 2522 734 2998 856
rect 3166 734 3734 856
rect 3902 734 4470 856
rect 4638 734 5206 856
rect 5374 734 5850 856
rect 6018 734 6586 856
rect 6754 734 7322 856
rect 7490 734 8058 856
rect 8226 734 8702 856
rect 8870 734 9438 856
rect 9606 734 10174 856
rect 10342 734 10910 856
rect 11078 734 11554 856
rect 11722 734 12290 856
rect 12458 734 13026 856
rect 13194 734 13762 856
rect 13930 734 14406 856
rect 14574 734 15142 856
rect 15310 734 15878 856
rect 16046 734 16614 856
rect 16782 734 17258 856
rect 17426 734 17994 856
rect 18162 734 18730 856
rect 18898 734 19466 856
rect 19634 734 20110 856
rect 20278 734 20846 856
rect 21014 734 21582 856
rect 21750 734 22318 856
rect 22486 734 22962 856
rect 23130 734 23698 856
rect 23866 734 24434 856
rect 24602 734 25170 856
rect 25338 734 25814 856
rect 25982 734 26550 856
rect 26718 734 27286 856
rect 27454 734 28022 856
rect 28190 734 28666 856
rect 28834 734 29402 856
rect 29570 734 30138 856
rect 30306 734 30874 856
rect 31042 734 31518 856
rect 31686 734 32254 856
rect 32422 734 32990 856
rect 33158 734 33726 856
rect 33894 734 34370 856
rect 34538 734 35106 856
rect 35274 734 35842 856
rect 36010 734 36578 856
rect 36746 734 37222 856
rect 37390 734 37958 856
rect 38126 734 38694 856
rect 38862 734 39430 856
rect 39598 734 40074 856
rect 40242 734 40810 856
rect 40978 734 41546 856
rect 41714 734 42282 856
rect 42450 734 42926 856
rect 43094 734 43662 856
rect 43830 734 44398 856
rect 44566 734 45134 856
rect 45302 734 45778 856
rect 45946 734 46514 856
rect 46682 734 47250 856
rect 47418 734 47986 856
rect 48154 734 48630 856
rect 48798 734 49366 856
rect 49534 734 50102 856
rect 50270 734 50746 856
rect 50914 734 51482 856
rect 51650 734 52218 856
rect 52386 734 52954 856
rect 53122 734 53598 856
rect 53766 734 54334 856
rect 54502 734 55070 856
rect 55238 734 55806 856
rect 55974 734 56450 856
rect 56618 734 57186 856
rect 57354 734 57922 856
rect 58090 734 58658 856
rect 58826 734 59302 856
rect 59470 734 60038 856
rect 60206 734 60774 856
rect 60942 734 61510 856
rect 61678 734 62154 856
rect 62322 734 62890 856
rect 63058 734 63626 856
rect 63794 734 64362 856
rect 64530 734 65006 856
rect 65174 734 65742 856
rect 65910 734 66478 856
rect 66646 734 67214 856
rect 67382 734 67858 856
rect 68026 734 68594 856
rect 68762 734 69330 856
rect 69498 734 70066 856
rect 70234 734 70710 856
rect 70878 734 71446 856
rect 71614 734 72182 856
rect 72350 734 72918 856
rect 73086 734 73562 856
rect 73730 734 74298 856
rect 74466 734 75034 856
rect 75202 734 75770 856
rect 75938 734 76414 856
rect 76582 734 77150 856
rect 77318 734 77886 856
rect 78054 734 78622 856
rect 78790 734 79266 856
rect 79434 734 80002 856
rect 80170 734 80738 856
rect 80906 734 81474 856
rect 81642 734 82118 856
rect 82286 734 82854 856
rect 83022 734 83590 856
rect 83758 734 84326 856
rect 84494 734 84970 856
rect 85138 734 85706 856
rect 85874 734 86442 856
rect 86610 734 87178 856
rect 87346 734 87822 856
rect 87990 734 88558 856
rect 88726 734 89294 856
rect 89462 734 90030 856
rect 90198 734 90674 856
rect 90842 734 91410 856
rect 91578 734 92146 856
rect 92314 734 92882 856
rect 93050 734 93526 856
rect 93694 734 94262 856
rect 94430 734 94998 856
rect 95166 734 95734 856
rect 95902 734 96378 856
rect 96546 734 97114 856
rect 97282 734 97850 856
rect 98018 734 98586 856
rect 98754 734 99230 856
rect 99398 734 99966 856
rect 100134 734 100702 856
rect 100870 734 101346 856
rect 101514 734 102082 856
rect 102250 734 102818 856
rect 102986 734 103554 856
rect 103722 734 104198 856
rect 104366 734 104934 856
rect 105102 734 105670 856
rect 105838 734 106406 856
rect 106574 734 107050 856
rect 107218 734 107786 856
rect 107954 734 108522 856
rect 108690 734 109258 856
rect 109426 734 109902 856
rect 110070 734 110638 856
rect 110806 734 111374 856
rect 111542 734 112110 856
rect 112278 734 112754 856
rect 112922 734 113490 856
rect 113658 734 114226 856
rect 114394 734 114962 856
rect 115130 734 115606 856
rect 115774 734 116342 856
rect 116510 734 117078 856
rect 117246 734 117814 856
rect 117982 734 118458 856
rect 118626 734 119194 856
rect 119362 734 119930 856
rect 120098 734 120666 856
rect 120834 734 121310 856
rect 121478 734 122046 856
rect 122214 734 122782 856
rect 122950 734 123518 856
rect 123686 734 124162 856
rect 124330 734 124898 856
rect 125066 734 125634 856
rect 125802 734 126370 856
rect 126538 734 127014 856
rect 127182 734 127750 856
rect 127918 734 128486 856
rect 128654 734 129222 856
rect 129390 734 129866 856
rect 130034 734 130602 856
rect 130770 734 131338 856
rect 131506 734 132074 856
rect 132242 734 132718 856
rect 132886 734 133454 856
rect 133622 734 134190 856
rect 134358 734 134926 856
rect 135094 734 135570 856
rect 135738 734 136306 856
rect 136474 734 137042 856
rect 137210 734 137778 856
rect 137946 734 138422 856
rect 138590 734 139158 856
rect 139326 734 139894 856
rect 140062 734 140630 856
rect 140798 734 141274 856
rect 141442 734 142010 856
rect 142178 734 142746 856
rect 142914 734 143482 856
rect 143650 734 144126 856
rect 144294 734 144862 856
rect 145030 734 145598 856
rect 145766 734 146334 856
rect 146502 734 146978 856
rect 147146 734 147714 856
rect 147882 734 148450 856
rect 148618 734 149186 856
rect 149354 734 149830 856
rect 149998 734 150566 856
rect 150734 734 151302 856
rect 151470 734 151946 856
rect 152114 734 152682 856
rect 152850 734 153418 856
rect 153586 734 154154 856
rect 154322 734 154798 856
rect 154966 734 155534 856
rect 155702 734 156270 856
rect 156438 734 157006 856
rect 157174 734 157650 856
rect 157818 734 158386 856
rect 158554 734 159122 856
rect 159290 734 159858 856
rect 160026 734 160502 856
rect 160670 734 161238 856
rect 161406 734 161974 856
rect 162142 734 162710 856
rect 162878 734 163354 856
rect 163522 734 164090 856
rect 164258 734 164826 856
rect 164994 734 165562 856
rect 165730 734 166206 856
rect 166374 734 166942 856
rect 167110 734 167678 856
rect 167846 734 168414 856
rect 168582 734 169058 856
rect 169226 734 169794 856
rect 169962 734 170530 856
rect 170698 734 171266 856
rect 171434 734 171910 856
rect 172078 734 172646 856
rect 172814 734 173382 856
rect 173550 734 174118 856
rect 174286 734 174762 856
rect 174930 734 175498 856
rect 175666 734 176234 856
rect 176402 734 176970 856
rect 177138 734 177614 856
rect 177782 734 178350 856
rect 178518 734 179086 856
rect 179254 734 179822 856
rect 179990 734 180466 856
rect 180634 734 181202 856
rect 181370 734 181938 856
rect 182106 734 182674 856
rect 182842 734 183318 856
rect 183486 734 184054 856
rect 184222 734 184790 856
rect 184958 734 185526 856
rect 185694 734 186170 856
rect 186338 734 186906 856
rect 187074 734 187642 856
rect 187810 734 188378 856
rect 188546 734 189022 856
rect 189190 734 189758 856
rect 189926 734 190494 856
rect 190662 734 191230 856
rect 191398 734 191874 856
rect 192042 734 192610 856
rect 192778 734 193346 856
rect 193514 734 194082 856
rect 194250 734 194726 856
rect 194894 734 195462 856
rect 195630 734 196198 856
rect 196366 734 196934 856
rect 197102 734 197578 856
rect 197746 734 198314 856
rect 198482 734 199050 856
rect 199218 734 199786 856
rect 199954 734 200430 856
rect 200598 734 201166 856
rect 201334 734 201902 856
rect 202070 734 202546 856
rect 202714 734 203282 856
rect 203450 734 204018 856
rect 204186 734 204754 856
rect 204922 734 205398 856
rect 205566 734 206134 856
rect 206302 734 206870 856
rect 207038 734 207606 856
rect 207774 734 208250 856
rect 208418 734 208986 856
rect 209154 734 209722 856
rect 209890 734 210458 856
rect 210626 734 211102 856
rect 211270 734 211838 856
rect 212006 734 212574 856
rect 212742 734 213310 856
rect 213478 734 213954 856
rect 214122 734 214690 856
rect 214858 734 215426 856
rect 215594 734 216162 856
rect 216330 734 216806 856
rect 216974 734 217542 856
rect 217710 734 218278 856
rect 218446 734 219014 856
rect 219182 734 219658 856
rect 219826 734 220394 856
rect 220562 734 221130 856
rect 221298 734 221866 856
rect 222034 734 222510 856
rect 222678 734 223246 856
rect 223414 734 223982 856
rect 224150 734 224718 856
rect 224886 734 225362 856
rect 225530 734 226098 856
rect 226266 734 226834 856
rect 227002 734 227570 856
rect 227738 734 228214 856
rect 228382 734 228950 856
rect 229118 734 229686 856
rect 229854 734 230422 856
rect 230590 734 231066 856
rect 231234 734 231802 856
rect 231970 734 232538 856
rect 232706 734 233274 856
rect 233442 734 233918 856
rect 234086 734 234654 856
rect 234822 734 235390 856
rect 235558 734 236126 856
rect 236294 734 236770 856
rect 236938 734 237506 856
rect 237674 734 238242 856
rect 238410 734 238978 856
rect 239146 734 239622 856
rect 239790 734 240358 856
rect 240526 734 241094 856
rect 241262 734 241830 856
rect 241998 734 242474 856
rect 242642 734 243210 856
rect 243378 734 243946 856
rect 244114 734 244682 856
rect 244850 734 245326 856
rect 245494 734 246062 856
rect 246230 734 246798 856
rect 246966 734 247534 856
rect 247702 734 248178 856
rect 248346 734 248914 856
rect 249082 734 249650 856
rect 249818 734 250386 856
rect 250554 734 251030 856
rect 251198 734 251766 856
rect 251934 734 252502 856
rect 252670 734 253146 856
rect 253314 734 253882 856
rect 254050 734 254618 856
rect 254786 734 255354 856
rect 255522 734 255998 856
rect 256166 734 256734 856
rect 256902 734 257470 856
rect 257638 734 258206 856
rect 258374 734 258850 856
rect 259018 734 259586 856
rect 259754 734 260322 856
rect 260490 734 261058 856
rect 261226 734 261702 856
rect 261870 734 262438 856
rect 262606 734 263174 856
rect 263342 734 263910 856
rect 264078 734 264554 856
rect 264722 734 265290 856
rect 265458 734 266026 856
rect 266194 734 266762 856
rect 266930 734 267406 856
rect 267574 734 268142 856
rect 268310 734 268878 856
rect 269046 734 269614 856
rect 269782 734 270258 856
rect 270426 734 270994 856
rect 271162 734 271730 856
rect 271898 734 272466 856
rect 272634 734 273110 856
rect 273278 734 273846 856
rect 274014 734 274582 856
rect 274750 734 275318 856
rect 275486 734 275962 856
rect 276130 734 276698 856
rect 276866 734 277434 856
rect 277602 734 278170 856
rect 278338 734 278814 856
rect 278982 734 279550 856
rect 279718 734 280286 856
rect 280454 734 281022 856
rect 281190 734 281666 856
rect 281834 734 282402 856
rect 282570 734 283138 856
rect 283306 734 283874 856
rect 284042 734 284518 856
rect 284686 734 285254 856
rect 285422 734 285990 856
rect 286158 734 286726 856
rect 286894 734 287370 856
rect 287538 734 288106 856
rect 288274 734 288842 856
rect 289010 734 289578 856
rect 289746 734 290222 856
rect 290390 734 290958 856
rect 291126 734 291694 856
rect 291862 734 292430 856
rect 292598 734 293074 856
rect 293242 734 293810 856
rect 293978 734 294546 856
rect 294714 734 295282 856
rect 295450 734 295926 856
rect 296094 734 296662 856
rect 296830 734 297398 856
rect 297566 734 298134 856
rect 298302 734 298778 856
rect 298946 734 299514 856
rect 299682 734 300250 856
rect 300418 734 300986 856
rect 301154 734 301630 856
rect 301798 734 302366 856
rect 302534 734 303102 856
rect 303270 734 303746 856
rect 303914 734 304482 856
rect 304650 734 305218 856
rect 305386 734 305954 856
rect 306122 734 306598 856
rect 306766 734 307334 856
rect 307502 734 308070 856
rect 308238 734 308806 856
rect 308974 734 309450 856
rect 309618 734 310186 856
rect 310354 734 310922 856
rect 311090 734 311658 856
rect 311826 734 312302 856
rect 312470 734 313038 856
rect 313206 734 313774 856
rect 313942 734 314510 856
rect 314678 734 315154 856
rect 315322 734 315890 856
rect 316058 734 316626 856
rect 316794 734 317362 856
rect 317530 734 318006 856
rect 318174 734 318742 856
rect 318910 734 319478 856
rect 319646 734 320214 856
rect 320382 734 320858 856
rect 321026 734 321594 856
rect 321762 734 322330 856
rect 322498 734 323066 856
rect 323234 734 323710 856
rect 323878 734 324446 856
rect 324614 734 325182 856
rect 325350 734 325918 856
rect 326086 734 326562 856
rect 326730 734 327298 856
rect 327466 734 328034 856
rect 328202 734 328770 856
rect 328938 734 329414 856
rect 329582 734 330150 856
rect 330318 734 330886 856
rect 331054 734 331622 856
rect 331790 734 332266 856
rect 332434 734 333002 856
rect 333170 734 333738 856
rect 333906 734 334474 856
rect 334642 734 335118 856
rect 335286 734 335854 856
rect 336022 734 336590 856
rect 336758 734 337326 856
rect 337494 734 337970 856
rect 338138 734 338706 856
rect 338874 734 339442 856
rect 339610 734 340178 856
rect 340346 734 340822 856
rect 340990 734 341558 856
rect 341726 734 342294 856
rect 342462 734 343030 856
rect 343198 734 343674 856
rect 343842 734 344410 856
rect 344578 734 345146 856
rect 345314 734 345882 856
rect 346050 734 346526 856
rect 346694 734 347262 856
rect 347430 734 347998 856
rect 348166 734 348734 856
rect 348902 734 349378 856
rect 349546 734 350114 856
rect 350282 734 350850 856
<< metal3 >>
rect 0 352520 800 352640
rect 0 351024 800 351144
rect 0 349392 800 349512
rect 0 347896 800 348016
rect 0 346264 800 346384
rect 0 344768 800 344888
rect 0 343136 800 343256
rect 0 341640 800 341760
rect 0 340008 800 340128
rect 0 338512 800 338632
rect 0 336880 800 337000
rect 0 335384 800 335504
rect 0 333752 800 333872
rect 0 332256 800 332376
rect 0 330624 800 330744
rect 0 329128 800 329248
rect 0 327496 800 327616
rect 0 326000 800 326120
rect 0 324368 800 324488
rect 0 322872 800 322992
rect 0 321240 800 321360
rect 0 319744 800 319864
rect 0 318112 800 318232
rect 0 316616 800 316736
rect 0 314984 800 315104
rect 0 313488 800 313608
rect 0 311856 800 311976
rect 0 310360 800 310480
rect 0 308728 800 308848
rect 0 307232 800 307352
rect 0 305600 800 305720
rect 0 304104 800 304224
rect 0 302472 800 302592
rect 0 300976 800 301096
rect 0 299344 800 299464
rect 0 297848 800 297968
rect 0 296216 800 296336
rect 0 294720 800 294840
rect 0 293088 800 293208
rect 0 291592 800 291712
rect 0 289960 800 290080
rect 0 288464 800 288584
rect 0 286832 800 286952
rect 0 285336 800 285456
rect 0 283704 800 283824
rect 0 282208 800 282328
rect 0 280576 800 280696
rect 0 279080 800 279200
rect 0 277448 800 277568
rect 0 275952 800 276072
rect 0 274320 800 274440
rect 0 272824 800 272944
rect 0 271192 800 271312
rect 0 269696 800 269816
rect 0 268064 800 268184
rect 0 266568 800 266688
rect 0 264936 800 265056
rect 0 263440 800 263560
rect 0 261808 800 261928
rect 0 260312 800 260432
rect 0 258680 800 258800
rect 0 257184 800 257304
rect 0 255552 800 255672
rect 0 254056 800 254176
rect 0 252424 800 252544
rect 0 250928 800 251048
rect 0 249296 800 249416
rect 0 247800 800 247920
rect 0 246168 800 246288
rect 0 244672 800 244792
rect 0 243040 800 243160
rect 0 241544 800 241664
rect 0 239912 800 240032
rect 0 238416 800 238536
rect 0 236784 800 236904
rect 0 235288 800 235408
rect 0 233656 800 233776
rect 0 232160 800 232280
rect 0 230528 800 230648
rect 0 229032 800 229152
rect 0 227400 800 227520
rect 0 225904 800 226024
rect 0 224272 800 224392
rect 0 222776 800 222896
rect 0 221144 800 221264
rect 0 219648 800 219768
rect 0 218016 800 218136
rect 0 216520 800 216640
rect 0 214888 800 215008
rect 0 213392 800 213512
rect 0 211760 800 211880
rect 0 210264 800 210384
rect 0 208632 800 208752
rect 0 207136 800 207256
rect 0 205504 800 205624
rect 0 204008 800 204128
rect 0 202376 800 202496
rect 0 200880 800 201000
rect 0 199248 800 199368
rect 0 197752 800 197872
rect 0 196120 800 196240
rect 0 194624 800 194744
rect 0 192992 800 193112
rect 0 191496 800 191616
rect 0 189864 800 189984
rect 0 188368 800 188488
rect 0 186736 800 186856
rect 0 185240 800 185360
rect 0 183608 800 183728
rect 0 182112 800 182232
rect 0 180480 800 180600
rect 0 178984 800 179104
rect 0 177352 800 177472
rect 0 175856 800 175976
rect 0 174224 800 174344
rect 0 172728 800 172848
rect 0 171096 800 171216
rect 0 169600 800 169720
rect 0 167968 800 168088
rect 0 166472 800 166592
rect 0 164840 800 164960
rect 0 163344 800 163464
rect 0 161712 800 161832
rect 0 160216 800 160336
rect 0 158584 800 158704
rect 0 157088 800 157208
rect 0 155456 800 155576
rect 0 153960 800 154080
rect 0 152328 800 152448
rect 0 150832 800 150952
rect 0 149200 800 149320
rect 0 147704 800 147824
rect 0 146072 800 146192
rect 0 144576 800 144696
rect 0 142944 800 143064
rect 0 141448 800 141568
rect 0 139816 800 139936
rect 0 138320 800 138440
rect 0 136688 800 136808
rect 0 135192 800 135312
rect 0 133560 800 133680
rect 0 132064 800 132184
rect 0 130432 800 130552
rect 0 128936 800 129056
rect 0 127304 800 127424
rect 0 125808 800 125928
rect 0 124176 800 124296
rect 0 122680 800 122800
rect 0 121048 800 121168
rect 0 119552 800 119672
rect 0 117920 800 118040
rect 0 116424 800 116544
rect 0 114792 800 114912
rect 0 113296 800 113416
rect 0 111664 800 111784
rect 0 110168 800 110288
rect 0 108536 800 108656
rect 0 107040 800 107160
rect 0 105408 800 105528
rect 0 103912 800 104032
rect 0 102280 800 102400
rect 0 100784 800 100904
rect 0 99152 800 99272
rect 0 97656 800 97776
rect 0 96024 800 96144
rect 0 94528 800 94648
rect 0 92896 800 93016
rect 0 91400 800 91520
rect 0 89768 800 89888
rect 0 88272 800 88392
rect 0 86640 800 86760
rect 0 85144 800 85264
rect 0 83512 800 83632
rect 0 82016 800 82136
rect 0 80384 800 80504
rect 0 78888 800 79008
rect 0 77256 800 77376
rect 0 75760 800 75880
rect 0 74128 800 74248
rect 0 72632 800 72752
rect 0 71000 800 71120
rect 0 69504 800 69624
rect 0 67872 800 67992
rect 0 66376 800 66496
rect 0 64744 800 64864
rect 0 63248 800 63368
rect 0 61616 800 61736
rect 0 60120 800 60240
rect 0 58488 800 58608
rect 0 56992 800 57112
rect 0 55360 800 55480
rect 0 53864 800 53984
rect 0 52232 800 52352
rect 0 50736 800 50856
rect 0 49104 800 49224
rect 0 47608 800 47728
rect 0 45976 800 46096
rect 0 44480 800 44600
rect 0 42848 800 42968
rect 0 41352 800 41472
rect 0 39720 800 39840
rect 0 38224 800 38344
rect 0 36592 800 36712
rect 0 35096 800 35216
rect 0 33464 800 33584
rect 0 31968 800 32088
rect 0 30336 800 30456
rect 0 28840 800 28960
rect 0 27208 800 27328
rect 0 25712 800 25832
rect 0 24080 800 24200
rect 0 22584 800 22704
rect 0 20952 800 21072
rect 0 19456 800 19576
rect 0 17824 800 17944
rect 0 16328 800 16448
rect 0 14696 800 14816
rect 0 13200 800 13320
rect 0 11568 800 11688
rect 0 10072 800 10192
rect 0 8440 800 8560
rect 0 6944 800 7064
rect 0 5312 800 5432
rect 0 3816 800 3936
rect 0 2184 800 2304
rect 0 688 800 808
<< obsm3 >>
rect 381 352720 348299 353429
rect 880 352440 348299 352720
rect 381 351224 348299 352440
rect 880 350944 348299 351224
rect 381 349592 348299 350944
rect 880 349312 348299 349592
rect 381 348096 348299 349312
rect 880 347816 348299 348096
rect 381 346464 348299 347816
rect 880 346184 348299 346464
rect 381 344968 348299 346184
rect 880 344688 348299 344968
rect 381 343336 348299 344688
rect 880 343056 348299 343336
rect 381 341840 348299 343056
rect 880 341560 348299 341840
rect 381 340208 348299 341560
rect 880 339928 348299 340208
rect 381 338712 348299 339928
rect 880 338432 348299 338712
rect 381 337080 348299 338432
rect 880 336800 348299 337080
rect 381 335584 348299 336800
rect 880 335304 348299 335584
rect 381 333952 348299 335304
rect 880 333672 348299 333952
rect 381 332456 348299 333672
rect 880 332176 348299 332456
rect 381 330824 348299 332176
rect 880 330544 348299 330824
rect 381 329328 348299 330544
rect 880 329048 348299 329328
rect 381 327696 348299 329048
rect 880 327416 348299 327696
rect 381 326200 348299 327416
rect 880 325920 348299 326200
rect 381 324568 348299 325920
rect 880 324288 348299 324568
rect 381 323072 348299 324288
rect 880 322792 348299 323072
rect 381 321440 348299 322792
rect 880 321160 348299 321440
rect 381 319944 348299 321160
rect 880 319664 348299 319944
rect 381 318312 348299 319664
rect 880 318032 348299 318312
rect 381 316816 348299 318032
rect 880 316536 348299 316816
rect 381 315184 348299 316536
rect 880 314904 348299 315184
rect 381 313688 348299 314904
rect 880 313408 348299 313688
rect 381 312056 348299 313408
rect 880 311776 348299 312056
rect 381 310560 348299 311776
rect 880 310280 348299 310560
rect 381 308928 348299 310280
rect 880 308648 348299 308928
rect 381 307432 348299 308648
rect 880 307152 348299 307432
rect 381 305800 348299 307152
rect 880 305520 348299 305800
rect 381 304304 348299 305520
rect 880 304024 348299 304304
rect 381 302672 348299 304024
rect 880 302392 348299 302672
rect 381 301176 348299 302392
rect 880 300896 348299 301176
rect 381 299544 348299 300896
rect 880 299264 348299 299544
rect 381 298048 348299 299264
rect 880 297768 348299 298048
rect 381 296416 348299 297768
rect 880 296136 348299 296416
rect 381 294920 348299 296136
rect 880 294640 348299 294920
rect 381 293288 348299 294640
rect 880 293008 348299 293288
rect 381 291792 348299 293008
rect 880 291512 348299 291792
rect 381 290160 348299 291512
rect 880 289880 348299 290160
rect 381 288664 348299 289880
rect 880 288384 348299 288664
rect 381 287032 348299 288384
rect 880 286752 348299 287032
rect 381 285536 348299 286752
rect 880 285256 348299 285536
rect 381 283904 348299 285256
rect 880 283624 348299 283904
rect 381 282408 348299 283624
rect 880 282128 348299 282408
rect 381 280776 348299 282128
rect 880 280496 348299 280776
rect 381 279280 348299 280496
rect 880 279000 348299 279280
rect 381 277648 348299 279000
rect 880 277368 348299 277648
rect 381 276152 348299 277368
rect 880 275872 348299 276152
rect 381 274520 348299 275872
rect 880 274240 348299 274520
rect 381 273024 348299 274240
rect 880 272744 348299 273024
rect 381 271392 348299 272744
rect 880 271112 348299 271392
rect 381 269896 348299 271112
rect 880 269616 348299 269896
rect 381 268264 348299 269616
rect 880 267984 348299 268264
rect 381 266768 348299 267984
rect 880 266488 348299 266768
rect 381 265136 348299 266488
rect 880 264856 348299 265136
rect 381 263640 348299 264856
rect 880 263360 348299 263640
rect 381 262008 348299 263360
rect 880 261728 348299 262008
rect 381 260512 348299 261728
rect 880 260232 348299 260512
rect 381 258880 348299 260232
rect 880 258600 348299 258880
rect 381 257384 348299 258600
rect 880 257104 348299 257384
rect 381 255752 348299 257104
rect 880 255472 348299 255752
rect 381 254256 348299 255472
rect 880 253976 348299 254256
rect 381 252624 348299 253976
rect 880 252344 348299 252624
rect 381 251128 348299 252344
rect 880 250848 348299 251128
rect 381 249496 348299 250848
rect 880 249216 348299 249496
rect 381 248000 348299 249216
rect 880 247720 348299 248000
rect 381 246368 348299 247720
rect 880 246088 348299 246368
rect 381 244872 348299 246088
rect 880 244592 348299 244872
rect 381 243240 348299 244592
rect 880 242960 348299 243240
rect 381 241744 348299 242960
rect 880 241464 348299 241744
rect 381 240112 348299 241464
rect 880 239832 348299 240112
rect 381 238616 348299 239832
rect 880 238336 348299 238616
rect 381 236984 348299 238336
rect 880 236704 348299 236984
rect 381 235488 348299 236704
rect 880 235208 348299 235488
rect 381 233856 348299 235208
rect 880 233576 348299 233856
rect 381 232360 348299 233576
rect 880 232080 348299 232360
rect 381 230728 348299 232080
rect 880 230448 348299 230728
rect 381 229232 348299 230448
rect 880 228952 348299 229232
rect 381 227600 348299 228952
rect 880 227320 348299 227600
rect 381 226104 348299 227320
rect 880 225824 348299 226104
rect 381 224472 348299 225824
rect 880 224192 348299 224472
rect 381 222976 348299 224192
rect 880 222696 348299 222976
rect 381 221344 348299 222696
rect 880 221064 348299 221344
rect 381 219848 348299 221064
rect 880 219568 348299 219848
rect 381 218216 348299 219568
rect 880 217936 348299 218216
rect 381 216720 348299 217936
rect 880 216440 348299 216720
rect 381 215088 348299 216440
rect 880 214808 348299 215088
rect 381 213592 348299 214808
rect 880 213312 348299 213592
rect 381 211960 348299 213312
rect 880 211680 348299 211960
rect 381 210464 348299 211680
rect 880 210184 348299 210464
rect 381 208832 348299 210184
rect 880 208552 348299 208832
rect 381 207336 348299 208552
rect 880 207056 348299 207336
rect 381 205704 348299 207056
rect 880 205424 348299 205704
rect 381 204208 348299 205424
rect 880 203928 348299 204208
rect 381 202576 348299 203928
rect 880 202296 348299 202576
rect 381 201080 348299 202296
rect 880 200800 348299 201080
rect 381 199448 348299 200800
rect 880 199168 348299 199448
rect 381 197952 348299 199168
rect 880 197672 348299 197952
rect 381 196320 348299 197672
rect 880 196040 348299 196320
rect 381 194824 348299 196040
rect 880 194544 348299 194824
rect 381 193192 348299 194544
rect 880 192912 348299 193192
rect 381 191696 348299 192912
rect 880 191416 348299 191696
rect 381 190064 348299 191416
rect 880 189784 348299 190064
rect 381 188568 348299 189784
rect 880 188288 348299 188568
rect 381 186936 348299 188288
rect 880 186656 348299 186936
rect 381 185440 348299 186656
rect 880 185160 348299 185440
rect 381 183808 348299 185160
rect 880 183528 348299 183808
rect 381 182312 348299 183528
rect 880 182032 348299 182312
rect 381 180680 348299 182032
rect 880 180400 348299 180680
rect 381 179184 348299 180400
rect 880 178904 348299 179184
rect 381 177552 348299 178904
rect 880 177272 348299 177552
rect 381 176056 348299 177272
rect 880 175776 348299 176056
rect 381 174424 348299 175776
rect 880 174144 348299 174424
rect 381 172928 348299 174144
rect 880 172648 348299 172928
rect 381 171296 348299 172648
rect 880 171016 348299 171296
rect 381 169800 348299 171016
rect 880 169520 348299 169800
rect 381 168168 348299 169520
rect 880 167888 348299 168168
rect 381 166672 348299 167888
rect 880 166392 348299 166672
rect 381 165040 348299 166392
rect 880 164760 348299 165040
rect 381 163544 348299 164760
rect 880 163264 348299 163544
rect 381 161912 348299 163264
rect 880 161632 348299 161912
rect 381 160416 348299 161632
rect 880 160136 348299 160416
rect 381 158784 348299 160136
rect 880 158504 348299 158784
rect 381 157288 348299 158504
rect 880 157008 348299 157288
rect 381 155656 348299 157008
rect 880 155376 348299 155656
rect 381 154160 348299 155376
rect 880 153880 348299 154160
rect 381 152528 348299 153880
rect 880 152248 348299 152528
rect 381 151032 348299 152248
rect 880 150752 348299 151032
rect 381 149400 348299 150752
rect 880 149120 348299 149400
rect 381 147904 348299 149120
rect 880 147624 348299 147904
rect 381 146272 348299 147624
rect 880 145992 348299 146272
rect 381 144776 348299 145992
rect 880 144496 348299 144776
rect 381 143144 348299 144496
rect 880 142864 348299 143144
rect 381 141648 348299 142864
rect 880 141368 348299 141648
rect 381 140016 348299 141368
rect 880 139736 348299 140016
rect 381 138520 348299 139736
rect 880 138240 348299 138520
rect 381 136888 348299 138240
rect 880 136608 348299 136888
rect 381 135392 348299 136608
rect 880 135112 348299 135392
rect 381 133760 348299 135112
rect 880 133480 348299 133760
rect 381 132264 348299 133480
rect 880 131984 348299 132264
rect 381 130632 348299 131984
rect 880 130352 348299 130632
rect 381 129136 348299 130352
rect 880 128856 348299 129136
rect 381 127504 348299 128856
rect 880 127224 348299 127504
rect 381 126008 348299 127224
rect 880 125728 348299 126008
rect 381 124376 348299 125728
rect 880 124096 348299 124376
rect 381 122880 348299 124096
rect 880 122600 348299 122880
rect 381 121248 348299 122600
rect 880 120968 348299 121248
rect 381 119752 348299 120968
rect 880 119472 348299 119752
rect 381 118120 348299 119472
rect 880 117840 348299 118120
rect 381 116624 348299 117840
rect 880 116344 348299 116624
rect 381 114992 348299 116344
rect 880 114712 348299 114992
rect 381 113496 348299 114712
rect 880 113216 348299 113496
rect 381 111864 348299 113216
rect 880 111584 348299 111864
rect 381 110368 348299 111584
rect 880 110088 348299 110368
rect 381 108736 348299 110088
rect 880 108456 348299 108736
rect 381 107240 348299 108456
rect 880 106960 348299 107240
rect 381 105608 348299 106960
rect 880 105328 348299 105608
rect 381 104112 348299 105328
rect 880 103832 348299 104112
rect 381 102480 348299 103832
rect 880 102200 348299 102480
rect 381 100984 348299 102200
rect 880 100704 348299 100984
rect 381 99352 348299 100704
rect 880 99072 348299 99352
rect 381 97856 348299 99072
rect 880 97576 348299 97856
rect 381 96224 348299 97576
rect 880 95944 348299 96224
rect 381 94728 348299 95944
rect 880 94448 348299 94728
rect 381 93096 348299 94448
rect 880 92816 348299 93096
rect 381 91600 348299 92816
rect 880 91320 348299 91600
rect 381 89968 348299 91320
rect 880 89688 348299 89968
rect 381 88472 348299 89688
rect 880 88192 348299 88472
rect 381 86840 348299 88192
rect 880 86560 348299 86840
rect 381 85344 348299 86560
rect 880 85064 348299 85344
rect 381 83712 348299 85064
rect 880 83432 348299 83712
rect 381 82216 348299 83432
rect 880 81936 348299 82216
rect 381 80584 348299 81936
rect 880 80304 348299 80584
rect 381 79088 348299 80304
rect 880 78808 348299 79088
rect 381 77456 348299 78808
rect 880 77176 348299 77456
rect 381 75960 348299 77176
rect 880 75680 348299 75960
rect 381 74328 348299 75680
rect 880 74048 348299 74328
rect 381 72832 348299 74048
rect 880 72552 348299 72832
rect 381 71200 348299 72552
rect 880 70920 348299 71200
rect 381 69704 348299 70920
rect 880 69424 348299 69704
rect 381 68072 348299 69424
rect 880 67792 348299 68072
rect 381 66576 348299 67792
rect 880 66296 348299 66576
rect 381 64944 348299 66296
rect 880 64664 348299 64944
rect 381 63448 348299 64664
rect 880 63168 348299 63448
rect 381 61816 348299 63168
rect 880 61536 348299 61816
rect 381 60320 348299 61536
rect 880 60040 348299 60320
rect 381 58688 348299 60040
rect 880 58408 348299 58688
rect 381 57192 348299 58408
rect 880 56912 348299 57192
rect 381 55560 348299 56912
rect 880 55280 348299 55560
rect 381 54064 348299 55280
rect 880 53784 348299 54064
rect 381 52432 348299 53784
rect 880 52152 348299 52432
rect 381 50936 348299 52152
rect 880 50656 348299 50936
rect 381 49304 348299 50656
rect 880 49024 348299 49304
rect 381 47808 348299 49024
rect 880 47528 348299 47808
rect 381 46176 348299 47528
rect 880 45896 348299 46176
rect 381 44680 348299 45896
rect 880 44400 348299 44680
rect 381 43048 348299 44400
rect 880 42768 348299 43048
rect 381 41552 348299 42768
rect 880 41272 348299 41552
rect 381 39920 348299 41272
rect 880 39640 348299 39920
rect 381 38424 348299 39640
rect 880 38144 348299 38424
rect 381 36792 348299 38144
rect 880 36512 348299 36792
rect 381 35296 348299 36512
rect 880 35016 348299 35296
rect 381 33664 348299 35016
rect 880 33384 348299 33664
rect 381 32168 348299 33384
rect 880 31888 348299 32168
rect 381 30536 348299 31888
rect 880 30256 348299 30536
rect 381 29040 348299 30256
rect 880 28760 348299 29040
rect 381 27408 348299 28760
rect 880 27128 348299 27408
rect 381 25912 348299 27128
rect 880 25632 348299 25912
rect 381 24280 348299 25632
rect 880 24000 348299 24280
rect 381 22784 348299 24000
rect 880 22504 348299 22784
rect 381 21152 348299 22504
rect 880 20872 348299 21152
rect 381 19656 348299 20872
rect 880 19376 348299 19656
rect 381 18024 348299 19376
rect 880 17744 348299 18024
rect 381 16528 348299 17744
rect 880 16248 348299 16528
rect 381 14896 348299 16248
rect 880 14616 348299 14896
rect 381 13400 348299 14616
rect 880 13120 348299 13400
rect 381 11768 348299 13120
rect 880 11488 348299 11768
rect 381 10272 348299 11488
rect 880 9992 348299 10272
rect 381 8640 348299 9992
rect 880 8360 348299 8640
rect 381 7144 348299 8360
rect 880 6864 348299 7144
rect 381 5512 348299 6864
rect 880 5232 348299 5512
rect 381 4016 348299 5232
rect 880 3736 348299 4016
rect 381 2384 348299 3736
rect 880 2104 348299 2384
rect 381 888 348299 2104
rect 880 718 348299 888
<< metal4 >>
rect 4208 2128 4528 350928
rect 19568 2128 19888 350928
rect 34928 2128 35248 350928
rect 50288 2128 50608 350928
rect 65648 2128 65968 350928
rect 81008 2128 81328 350928
rect 96368 2128 96688 350928
rect 111728 2128 112048 350928
rect 127088 2128 127408 350928
rect 142448 2128 142768 350928
rect 157808 2128 158128 350928
rect 173168 2128 173488 350928
rect 188528 2128 188848 350928
rect 203888 2128 204208 350928
rect 219248 2128 219568 350928
rect 234608 2128 234928 350928
rect 249968 2128 250288 350928
rect 265328 2128 265648 350928
rect 280688 2128 281008 350928
rect 296048 2128 296368 350928
rect 311408 2128 311728 350928
rect 326768 2128 327088 350928
rect 342128 2128 342448 350928
<< obsm4 >>
rect 427 351008 346781 353429
rect 427 2347 4128 351008
rect 4608 2347 19488 351008
rect 19968 2347 34848 351008
rect 35328 2347 50208 351008
rect 50688 2347 65568 351008
rect 66048 2347 80928 351008
rect 81408 2347 96288 351008
rect 96768 2347 111648 351008
rect 112128 2347 127008 351008
rect 127488 2347 142368 351008
rect 142848 2347 157728 351008
rect 158208 2347 173088 351008
rect 173568 2347 188448 351008
rect 188928 2347 203808 351008
rect 204288 2347 219168 351008
rect 219648 2347 234528 351008
rect 235008 2347 249888 351008
rect 250368 2347 265248 351008
rect 265728 2347 280608 351008
rect 281088 2347 295968 351008
rect 296448 2347 311328 351008
rect 311808 2347 326688 351008
rect 327168 2347 342048 351008
rect 342528 2347 346781 351008
<< labels >>
rlabel metal3 s 0 340008 800 340128 6 data_arrays_0_0_ext_ram_addr1[0]
port 1 nsew signal output
rlabel metal3 s 0 341640 800 341760 6 data_arrays_0_0_ext_ram_addr1[1]
port 2 nsew signal output
rlabel metal3 s 0 343136 800 343256 6 data_arrays_0_0_ext_ram_addr1[2]
port 3 nsew signal output
rlabel metal3 s 0 344768 800 344888 6 data_arrays_0_0_ext_ram_addr1[3]
port 4 nsew signal output
rlabel metal3 s 0 346264 800 346384 6 data_arrays_0_0_ext_ram_addr1[4]
port 5 nsew signal output
rlabel metal3 s 0 347896 800 348016 6 data_arrays_0_0_ext_ram_addr1[5]
port 6 nsew signal output
rlabel metal3 s 0 349392 800 349512 6 data_arrays_0_0_ext_ram_addr1[6]
port 7 nsew signal output
rlabel metal3 s 0 351024 800 351144 6 data_arrays_0_0_ext_ram_addr1[7]
port 8 nsew signal output
rlabel metal3 s 0 352520 800 352640 6 data_arrays_0_0_ext_ram_addr1[8]
port 9 nsew signal output
rlabel metal3 s 0 200880 800 201000 6 data_arrays_0_0_ext_ram_addr[0]
port 10 nsew signal output
rlabel metal3 s 0 202376 800 202496 6 data_arrays_0_0_ext_ram_addr[1]
port 11 nsew signal output
rlabel metal3 s 0 204008 800 204128 6 data_arrays_0_0_ext_ram_addr[2]
port 12 nsew signal output
rlabel metal3 s 0 205504 800 205624 6 data_arrays_0_0_ext_ram_addr[3]
port 13 nsew signal output
rlabel metal3 s 0 207136 800 207256 6 data_arrays_0_0_ext_ram_addr[4]
port 14 nsew signal output
rlabel metal3 s 0 208632 800 208752 6 data_arrays_0_0_ext_ram_addr[5]
port 15 nsew signal output
rlabel metal3 s 0 210264 800 210384 6 data_arrays_0_0_ext_ram_addr[6]
port 16 nsew signal output
rlabel metal3 s 0 211760 800 211880 6 data_arrays_0_0_ext_ram_addr[7]
port 17 nsew signal output
rlabel metal3 s 0 213392 800 213512 6 data_arrays_0_0_ext_ram_addr[8]
port 18 nsew signal output
rlabel metal3 s 0 214888 800 215008 6 data_arrays_0_0_ext_ram_clk
port 19 nsew signal output
rlabel metal3 s 0 327496 800 327616 6 data_arrays_0_0_ext_ram_csb1[0]
port 20 nsew signal output
rlabel metal3 s 0 329128 800 329248 6 data_arrays_0_0_ext_ram_csb1[1]
port 21 nsew signal output
rlabel metal3 s 0 330624 800 330744 6 data_arrays_0_0_ext_ram_csb1[2]
port 22 nsew signal output
rlabel metal3 s 0 332256 800 332376 6 data_arrays_0_0_ext_ram_csb1[3]
port 23 nsew signal output
rlabel metal3 s 0 333752 800 333872 6 data_arrays_0_0_ext_ram_csb1[4]
port 24 nsew signal output
rlabel metal3 s 0 335384 800 335504 6 data_arrays_0_0_ext_ram_csb1[5]
port 25 nsew signal output
rlabel metal3 s 0 336880 800 337000 6 data_arrays_0_0_ext_ram_csb1[6]
port 26 nsew signal output
rlabel metal3 s 0 338512 800 338632 6 data_arrays_0_0_ext_ram_csb1[7]
port 27 nsew signal output
rlabel metal3 s 0 319744 800 319864 6 data_arrays_0_0_ext_ram_csb[0]
port 28 nsew signal output
rlabel metal3 s 0 321240 800 321360 6 data_arrays_0_0_ext_ram_csb[1]
port 29 nsew signal output
rlabel metal3 s 0 322872 800 322992 6 data_arrays_0_0_ext_ram_csb[2]
port 30 nsew signal output
rlabel metal3 s 0 324368 800 324488 6 data_arrays_0_0_ext_ram_csb[3]
port 31 nsew signal output
rlabel metal3 s 0 688 800 808 6 data_arrays_0_0_ext_ram_rdata0[0]
port 32 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 data_arrays_0_0_ext_ram_rdata0[10]
port 33 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 data_arrays_0_0_ext_ram_rdata0[11]
port 34 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 data_arrays_0_0_ext_ram_rdata0[12]
port 35 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 data_arrays_0_0_ext_ram_rdata0[13]
port 36 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 data_arrays_0_0_ext_ram_rdata0[14]
port 37 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 data_arrays_0_0_ext_ram_rdata0[15]
port 38 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 data_arrays_0_0_ext_ram_rdata0[16]
port 39 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 data_arrays_0_0_ext_ram_rdata0[17]
port 40 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 data_arrays_0_0_ext_ram_rdata0[18]
port 41 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 data_arrays_0_0_ext_ram_rdata0[19]
port 42 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 data_arrays_0_0_ext_ram_rdata0[1]
port 43 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 data_arrays_0_0_ext_ram_rdata0[20]
port 44 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 data_arrays_0_0_ext_ram_rdata0[21]
port 45 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 data_arrays_0_0_ext_ram_rdata0[22]
port 46 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 data_arrays_0_0_ext_ram_rdata0[23]
port 47 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 data_arrays_0_0_ext_ram_rdata0[24]
port 48 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 data_arrays_0_0_ext_ram_rdata0[25]
port 49 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 data_arrays_0_0_ext_ram_rdata0[26]
port 50 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 data_arrays_0_0_ext_ram_rdata0[27]
port 51 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 data_arrays_0_0_ext_ram_rdata0[28]
port 52 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 data_arrays_0_0_ext_ram_rdata0[29]
port 53 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 data_arrays_0_0_ext_ram_rdata0[2]
port 54 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 data_arrays_0_0_ext_ram_rdata0[30]
port 55 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 data_arrays_0_0_ext_ram_rdata0[31]
port 56 nsew signal input
rlabel metal3 s 0 50736 800 50856 6 data_arrays_0_0_ext_ram_rdata0[32]
port 57 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 data_arrays_0_0_ext_ram_rdata0[33]
port 58 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 data_arrays_0_0_ext_ram_rdata0[34]
port 59 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 data_arrays_0_0_ext_ram_rdata0[35]
port 60 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 data_arrays_0_0_ext_ram_rdata0[36]
port 61 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 data_arrays_0_0_ext_ram_rdata0[37]
port 62 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 data_arrays_0_0_ext_ram_rdata0[38]
port 63 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 data_arrays_0_0_ext_ram_rdata0[39]
port 64 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 data_arrays_0_0_ext_ram_rdata0[3]
port 65 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 data_arrays_0_0_ext_ram_rdata0[40]
port 66 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 data_arrays_0_0_ext_ram_rdata0[41]
port 67 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 data_arrays_0_0_ext_ram_rdata0[42]
port 68 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 data_arrays_0_0_ext_ram_rdata0[43]
port 69 nsew signal input
rlabel metal3 s 0 69504 800 69624 6 data_arrays_0_0_ext_ram_rdata0[44]
port 70 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 data_arrays_0_0_ext_ram_rdata0[45]
port 71 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 data_arrays_0_0_ext_ram_rdata0[46]
port 72 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 data_arrays_0_0_ext_ram_rdata0[47]
port 73 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 data_arrays_0_0_ext_ram_rdata0[48]
port 74 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 data_arrays_0_0_ext_ram_rdata0[49]
port 75 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 data_arrays_0_0_ext_ram_rdata0[4]
port 76 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 data_arrays_0_0_ext_ram_rdata0[50]
port 77 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 data_arrays_0_0_ext_ram_rdata0[51]
port 78 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 data_arrays_0_0_ext_ram_rdata0[52]
port 79 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 data_arrays_0_0_ext_ram_rdata0[53]
port 80 nsew signal input
rlabel metal3 s 0 85144 800 85264 6 data_arrays_0_0_ext_ram_rdata0[54]
port 81 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 data_arrays_0_0_ext_ram_rdata0[55]
port 82 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 data_arrays_0_0_ext_ram_rdata0[56]
port 83 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 data_arrays_0_0_ext_ram_rdata0[57]
port 84 nsew signal input
rlabel metal3 s 0 91400 800 91520 6 data_arrays_0_0_ext_ram_rdata0[58]
port 85 nsew signal input
rlabel metal3 s 0 92896 800 93016 6 data_arrays_0_0_ext_ram_rdata0[59]
port 86 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 data_arrays_0_0_ext_ram_rdata0[5]
port 87 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 data_arrays_0_0_ext_ram_rdata0[60]
port 88 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 data_arrays_0_0_ext_ram_rdata0[61]
port 89 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 data_arrays_0_0_ext_ram_rdata0[62]
port 90 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 data_arrays_0_0_ext_ram_rdata0[63]
port 91 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 data_arrays_0_0_ext_ram_rdata0[6]
port 92 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 data_arrays_0_0_ext_ram_rdata0[7]
port 93 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 data_arrays_0_0_ext_ram_rdata0[8]
port 94 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 data_arrays_0_0_ext_ram_rdata0[9]
port 95 nsew signal input
rlabel metal3 s 0 100784 800 100904 6 data_arrays_0_0_ext_ram_rdata1[0]
port 96 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 data_arrays_0_0_ext_ram_rdata1[10]
port 97 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 data_arrays_0_0_ext_ram_rdata1[11]
port 98 nsew signal input
rlabel metal3 s 0 119552 800 119672 6 data_arrays_0_0_ext_ram_rdata1[12]
port 99 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 data_arrays_0_0_ext_ram_rdata1[13]
port 100 nsew signal input
rlabel metal3 s 0 122680 800 122800 6 data_arrays_0_0_ext_ram_rdata1[14]
port 101 nsew signal input
rlabel metal3 s 0 124176 800 124296 6 data_arrays_0_0_ext_ram_rdata1[15]
port 102 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 data_arrays_0_0_ext_ram_rdata1[16]
port 103 nsew signal input
rlabel metal3 s 0 127304 800 127424 6 data_arrays_0_0_ext_ram_rdata1[17]
port 104 nsew signal input
rlabel metal3 s 0 128936 800 129056 6 data_arrays_0_0_ext_ram_rdata1[18]
port 105 nsew signal input
rlabel metal3 s 0 130432 800 130552 6 data_arrays_0_0_ext_ram_rdata1[19]
port 106 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 data_arrays_0_0_ext_ram_rdata1[1]
port 107 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 data_arrays_0_0_ext_ram_rdata1[20]
port 108 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 data_arrays_0_0_ext_ram_rdata1[21]
port 109 nsew signal input
rlabel metal3 s 0 135192 800 135312 6 data_arrays_0_0_ext_ram_rdata1[22]
port 110 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 data_arrays_0_0_ext_ram_rdata1[23]
port 111 nsew signal input
rlabel metal3 s 0 138320 800 138440 6 data_arrays_0_0_ext_ram_rdata1[24]
port 112 nsew signal input
rlabel metal3 s 0 139816 800 139936 6 data_arrays_0_0_ext_ram_rdata1[25]
port 113 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 data_arrays_0_0_ext_ram_rdata1[26]
port 114 nsew signal input
rlabel metal3 s 0 142944 800 143064 6 data_arrays_0_0_ext_ram_rdata1[27]
port 115 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 data_arrays_0_0_ext_ram_rdata1[28]
port 116 nsew signal input
rlabel metal3 s 0 146072 800 146192 6 data_arrays_0_0_ext_ram_rdata1[29]
port 117 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 data_arrays_0_0_ext_ram_rdata1[2]
port 118 nsew signal input
rlabel metal3 s 0 147704 800 147824 6 data_arrays_0_0_ext_ram_rdata1[30]
port 119 nsew signal input
rlabel metal3 s 0 149200 800 149320 6 data_arrays_0_0_ext_ram_rdata1[31]
port 120 nsew signal input
rlabel metal3 s 0 150832 800 150952 6 data_arrays_0_0_ext_ram_rdata1[32]
port 121 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 data_arrays_0_0_ext_ram_rdata1[33]
port 122 nsew signal input
rlabel metal3 s 0 153960 800 154080 6 data_arrays_0_0_ext_ram_rdata1[34]
port 123 nsew signal input
rlabel metal3 s 0 155456 800 155576 6 data_arrays_0_0_ext_ram_rdata1[35]
port 124 nsew signal input
rlabel metal3 s 0 157088 800 157208 6 data_arrays_0_0_ext_ram_rdata1[36]
port 125 nsew signal input
rlabel metal3 s 0 158584 800 158704 6 data_arrays_0_0_ext_ram_rdata1[37]
port 126 nsew signal input
rlabel metal3 s 0 160216 800 160336 6 data_arrays_0_0_ext_ram_rdata1[38]
port 127 nsew signal input
rlabel metal3 s 0 161712 800 161832 6 data_arrays_0_0_ext_ram_rdata1[39]
port 128 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 data_arrays_0_0_ext_ram_rdata1[3]
port 129 nsew signal input
rlabel metal3 s 0 163344 800 163464 6 data_arrays_0_0_ext_ram_rdata1[40]
port 130 nsew signal input
rlabel metal3 s 0 164840 800 164960 6 data_arrays_0_0_ext_ram_rdata1[41]
port 131 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 data_arrays_0_0_ext_ram_rdata1[42]
port 132 nsew signal input
rlabel metal3 s 0 167968 800 168088 6 data_arrays_0_0_ext_ram_rdata1[43]
port 133 nsew signal input
rlabel metal3 s 0 169600 800 169720 6 data_arrays_0_0_ext_ram_rdata1[44]
port 134 nsew signal input
rlabel metal3 s 0 171096 800 171216 6 data_arrays_0_0_ext_ram_rdata1[45]
port 135 nsew signal input
rlabel metal3 s 0 172728 800 172848 6 data_arrays_0_0_ext_ram_rdata1[46]
port 136 nsew signal input
rlabel metal3 s 0 174224 800 174344 6 data_arrays_0_0_ext_ram_rdata1[47]
port 137 nsew signal input
rlabel metal3 s 0 175856 800 175976 6 data_arrays_0_0_ext_ram_rdata1[48]
port 138 nsew signal input
rlabel metal3 s 0 177352 800 177472 6 data_arrays_0_0_ext_ram_rdata1[49]
port 139 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 data_arrays_0_0_ext_ram_rdata1[4]
port 140 nsew signal input
rlabel metal3 s 0 178984 800 179104 6 data_arrays_0_0_ext_ram_rdata1[50]
port 141 nsew signal input
rlabel metal3 s 0 180480 800 180600 6 data_arrays_0_0_ext_ram_rdata1[51]
port 142 nsew signal input
rlabel metal3 s 0 182112 800 182232 6 data_arrays_0_0_ext_ram_rdata1[52]
port 143 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 data_arrays_0_0_ext_ram_rdata1[53]
port 144 nsew signal input
rlabel metal3 s 0 185240 800 185360 6 data_arrays_0_0_ext_ram_rdata1[54]
port 145 nsew signal input
rlabel metal3 s 0 186736 800 186856 6 data_arrays_0_0_ext_ram_rdata1[55]
port 146 nsew signal input
rlabel metal3 s 0 188368 800 188488 6 data_arrays_0_0_ext_ram_rdata1[56]
port 147 nsew signal input
rlabel metal3 s 0 189864 800 189984 6 data_arrays_0_0_ext_ram_rdata1[57]
port 148 nsew signal input
rlabel metal3 s 0 191496 800 191616 6 data_arrays_0_0_ext_ram_rdata1[58]
port 149 nsew signal input
rlabel metal3 s 0 192992 800 193112 6 data_arrays_0_0_ext_ram_rdata1[59]
port 150 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 data_arrays_0_0_ext_ram_rdata1[5]
port 151 nsew signal input
rlabel metal3 s 0 194624 800 194744 6 data_arrays_0_0_ext_ram_rdata1[60]
port 152 nsew signal input
rlabel metal3 s 0 196120 800 196240 6 data_arrays_0_0_ext_ram_rdata1[61]
port 153 nsew signal input
rlabel metal3 s 0 197752 800 197872 6 data_arrays_0_0_ext_ram_rdata1[62]
port 154 nsew signal input
rlabel metal3 s 0 199248 800 199368 6 data_arrays_0_0_ext_ram_rdata1[63]
port 155 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 data_arrays_0_0_ext_ram_rdata1[6]
port 156 nsew signal input
rlabel metal3 s 0 111664 800 111784 6 data_arrays_0_0_ext_ram_rdata1[7]
port 157 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 data_arrays_0_0_ext_ram_rdata1[8]
port 158 nsew signal input
rlabel metal3 s 0 114792 800 114912 6 data_arrays_0_0_ext_ram_rdata1[9]
port 159 nsew signal input
rlabel metal2 s 237286 352669 237342 353469 6 data_arrays_0_0_ext_ram_rdata2[0]
port 160 nsew signal input
rlabel metal2 s 246210 352669 246266 353469 6 data_arrays_0_0_ext_ram_rdata2[10]
port 161 nsew signal input
rlabel metal2 s 247130 352669 247186 353469 6 data_arrays_0_0_ext_ram_rdata2[11]
port 162 nsew signal input
rlabel metal2 s 247958 352669 248014 353469 6 data_arrays_0_0_ext_ram_rdata2[12]
port 163 nsew signal input
rlabel metal2 s 248878 352669 248934 353469 6 data_arrays_0_0_ext_ram_rdata2[13]
port 164 nsew signal input
rlabel metal2 s 249798 352669 249854 353469 6 data_arrays_0_0_ext_ram_rdata2[14]
port 165 nsew signal input
rlabel metal2 s 250626 352669 250682 353469 6 data_arrays_0_0_ext_ram_rdata2[15]
port 166 nsew signal input
rlabel metal2 s 251546 352669 251602 353469 6 data_arrays_0_0_ext_ram_rdata2[16]
port 167 nsew signal input
rlabel metal2 s 252466 352669 252522 353469 6 data_arrays_0_0_ext_ram_rdata2[17]
port 168 nsew signal input
rlabel metal2 s 253386 352669 253442 353469 6 data_arrays_0_0_ext_ram_rdata2[18]
port 169 nsew signal input
rlabel metal2 s 254214 352669 254270 353469 6 data_arrays_0_0_ext_ram_rdata2[19]
port 170 nsew signal input
rlabel metal2 s 238114 352669 238170 353469 6 data_arrays_0_0_ext_ram_rdata2[1]
port 171 nsew signal input
rlabel metal2 s 255134 352669 255190 353469 6 data_arrays_0_0_ext_ram_rdata2[20]
port 172 nsew signal input
rlabel metal2 s 256054 352669 256110 353469 6 data_arrays_0_0_ext_ram_rdata2[21]
port 173 nsew signal input
rlabel metal2 s 256882 352669 256938 353469 6 data_arrays_0_0_ext_ram_rdata2[22]
port 174 nsew signal input
rlabel metal2 s 257802 352669 257858 353469 6 data_arrays_0_0_ext_ram_rdata2[23]
port 175 nsew signal input
rlabel metal2 s 258722 352669 258778 353469 6 data_arrays_0_0_ext_ram_rdata2[24]
port 176 nsew signal input
rlabel metal2 s 259642 352669 259698 353469 6 data_arrays_0_0_ext_ram_rdata2[25]
port 177 nsew signal input
rlabel metal2 s 260470 352669 260526 353469 6 data_arrays_0_0_ext_ram_rdata2[26]
port 178 nsew signal input
rlabel metal2 s 261390 352669 261446 353469 6 data_arrays_0_0_ext_ram_rdata2[27]
port 179 nsew signal input
rlabel metal2 s 262310 352669 262366 353469 6 data_arrays_0_0_ext_ram_rdata2[28]
port 180 nsew signal input
rlabel metal2 s 263138 352669 263194 353469 6 data_arrays_0_0_ext_ram_rdata2[29]
port 181 nsew signal input
rlabel metal2 s 239034 352669 239090 353469 6 data_arrays_0_0_ext_ram_rdata2[2]
port 182 nsew signal input
rlabel metal2 s 264058 352669 264114 353469 6 data_arrays_0_0_ext_ram_rdata2[30]
port 183 nsew signal input
rlabel metal2 s 264978 352669 265034 353469 6 data_arrays_0_0_ext_ram_rdata2[31]
port 184 nsew signal input
rlabel metal2 s 265898 352669 265954 353469 6 data_arrays_0_0_ext_ram_rdata2[32]
port 185 nsew signal input
rlabel metal2 s 266726 352669 266782 353469 6 data_arrays_0_0_ext_ram_rdata2[33]
port 186 nsew signal input
rlabel metal2 s 267646 352669 267702 353469 6 data_arrays_0_0_ext_ram_rdata2[34]
port 187 nsew signal input
rlabel metal2 s 268566 352669 268622 353469 6 data_arrays_0_0_ext_ram_rdata2[35]
port 188 nsew signal input
rlabel metal2 s 269394 352669 269450 353469 6 data_arrays_0_0_ext_ram_rdata2[36]
port 189 nsew signal input
rlabel metal2 s 270314 352669 270370 353469 6 data_arrays_0_0_ext_ram_rdata2[37]
port 190 nsew signal input
rlabel metal2 s 271234 352669 271290 353469 6 data_arrays_0_0_ext_ram_rdata2[38]
port 191 nsew signal input
rlabel metal2 s 272154 352669 272210 353469 6 data_arrays_0_0_ext_ram_rdata2[39]
port 192 nsew signal input
rlabel metal2 s 239954 352669 240010 353469 6 data_arrays_0_0_ext_ram_rdata2[3]
port 193 nsew signal input
rlabel metal2 s 272982 352669 273038 353469 6 data_arrays_0_0_ext_ram_rdata2[40]
port 194 nsew signal input
rlabel metal2 s 273902 352669 273958 353469 6 data_arrays_0_0_ext_ram_rdata2[41]
port 195 nsew signal input
rlabel metal2 s 274822 352669 274878 353469 6 data_arrays_0_0_ext_ram_rdata2[42]
port 196 nsew signal input
rlabel metal2 s 275742 352669 275798 353469 6 data_arrays_0_0_ext_ram_rdata2[43]
port 197 nsew signal input
rlabel metal2 s 276570 352669 276626 353469 6 data_arrays_0_0_ext_ram_rdata2[44]
port 198 nsew signal input
rlabel metal2 s 277490 352669 277546 353469 6 data_arrays_0_0_ext_ram_rdata2[45]
port 199 nsew signal input
rlabel metal2 s 278410 352669 278466 353469 6 data_arrays_0_0_ext_ram_rdata2[46]
port 200 nsew signal input
rlabel metal2 s 279238 352669 279294 353469 6 data_arrays_0_0_ext_ram_rdata2[47]
port 201 nsew signal input
rlabel metal2 s 280158 352669 280214 353469 6 data_arrays_0_0_ext_ram_rdata2[48]
port 202 nsew signal input
rlabel metal2 s 281078 352669 281134 353469 6 data_arrays_0_0_ext_ram_rdata2[49]
port 203 nsew signal input
rlabel metal2 s 240874 352669 240930 353469 6 data_arrays_0_0_ext_ram_rdata2[4]
port 204 nsew signal input
rlabel metal2 s 281998 352669 282054 353469 6 data_arrays_0_0_ext_ram_rdata2[50]
port 205 nsew signal input
rlabel metal2 s 282826 352669 282882 353469 6 data_arrays_0_0_ext_ram_rdata2[51]
port 206 nsew signal input
rlabel metal2 s 283746 352669 283802 353469 6 data_arrays_0_0_ext_ram_rdata2[52]
port 207 nsew signal input
rlabel metal2 s 284666 352669 284722 353469 6 data_arrays_0_0_ext_ram_rdata2[53]
port 208 nsew signal input
rlabel metal2 s 285494 352669 285550 353469 6 data_arrays_0_0_ext_ram_rdata2[54]
port 209 nsew signal input
rlabel metal2 s 286414 352669 286470 353469 6 data_arrays_0_0_ext_ram_rdata2[55]
port 210 nsew signal input
rlabel metal2 s 287334 352669 287390 353469 6 data_arrays_0_0_ext_ram_rdata2[56]
port 211 nsew signal input
rlabel metal2 s 288254 352669 288310 353469 6 data_arrays_0_0_ext_ram_rdata2[57]
port 212 nsew signal input
rlabel metal2 s 289082 352669 289138 353469 6 data_arrays_0_0_ext_ram_rdata2[58]
port 213 nsew signal input
rlabel metal2 s 290002 352669 290058 353469 6 data_arrays_0_0_ext_ram_rdata2[59]
port 214 nsew signal input
rlabel metal2 s 241702 352669 241758 353469 6 data_arrays_0_0_ext_ram_rdata2[5]
port 215 nsew signal input
rlabel metal2 s 290922 352669 290978 353469 6 data_arrays_0_0_ext_ram_rdata2[60]
port 216 nsew signal input
rlabel metal2 s 291750 352669 291806 353469 6 data_arrays_0_0_ext_ram_rdata2[61]
port 217 nsew signal input
rlabel metal2 s 292670 352669 292726 353469 6 data_arrays_0_0_ext_ram_rdata2[62]
port 218 nsew signal input
rlabel metal2 s 293590 352669 293646 353469 6 data_arrays_0_0_ext_ram_rdata2[63]
port 219 nsew signal input
rlabel metal2 s 242622 352669 242678 353469 6 data_arrays_0_0_ext_ram_rdata2[6]
port 220 nsew signal input
rlabel metal2 s 243542 352669 243598 353469 6 data_arrays_0_0_ext_ram_rdata2[7]
port 221 nsew signal input
rlabel metal2 s 244370 352669 244426 353469 6 data_arrays_0_0_ext_ram_rdata2[8]
port 222 nsew signal input
rlabel metal2 s 245290 352669 245346 353469 6 data_arrays_0_0_ext_ram_rdata2[9]
port 223 nsew signal input
rlabel metal2 s 294510 352669 294566 353469 6 data_arrays_0_0_ext_ram_rdata3[0]
port 224 nsew signal input
rlabel metal2 s 303434 352669 303490 353469 6 data_arrays_0_0_ext_ram_rdata3[10]
port 225 nsew signal input
rlabel metal2 s 304262 352669 304318 353469 6 data_arrays_0_0_ext_ram_rdata3[11]
port 226 nsew signal input
rlabel metal2 s 305182 352669 305238 353469 6 data_arrays_0_0_ext_ram_rdata3[12]
port 227 nsew signal input
rlabel metal2 s 306102 352669 306158 353469 6 data_arrays_0_0_ext_ram_rdata3[13]
port 228 nsew signal input
rlabel metal2 s 307022 352669 307078 353469 6 data_arrays_0_0_ext_ram_rdata3[14]
port 229 nsew signal input
rlabel metal2 s 307850 352669 307906 353469 6 data_arrays_0_0_ext_ram_rdata3[15]
port 230 nsew signal input
rlabel metal2 s 308770 352669 308826 353469 6 data_arrays_0_0_ext_ram_rdata3[16]
port 231 nsew signal input
rlabel metal2 s 309690 352669 309746 353469 6 data_arrays_0_0_ext_ram_rdata3[17]
port 232 nsew signal input
rlabel metal2 s 310518 352669 310574 353469 6 data_arrays_0_0_ext_ram_rdata3[18]
port 233 nsew signal input
rlabel metal2 s 311438 352669 311494 353469 6 data_arrays_0_0_ext_ram_rdata3[19]
port 234 nsew signal input
rlabel metal2 s 295338 352669 295394 353469 6 data_arrays_0_0_ext_ram_rdata3[1]
port 235 nsew signal input
rlabel metal2 s 312358 352669 312414 353469 6 data_arrays_0_0_ext_ram_rdata3[20]
port 236 nsew signal input
rlabel metal2 s 313278 352669 313334 353469 6 data_arrays_0_0_ext_ram_rdata3[21]
port 237 nsew signal input
rlabel metal2 s 314106 352669 314162 353469 6 data_arrays_0_0_ext_ram_rdata3[22]
port 238 nsew signal input
rlabel metal2 s 315026 352669 315082 353469 6 data_arrays_0_0_ext_ram_rdata3[23]
port 239 nsew signal input
rlabel metal2 s 315946 352669 316002 353469 6 data_arrays_0_0_ext_ram_rdata3[24]
port 240 nsew signal input
rlabel metal2 s 316866 352669 316922 353469 6 data_arrays_0_0_ext_ram_rdata3[25]
port 241 nsew signal input
rlabel metal2 s 317694 352669 317750 353469 6 data_arrays_0_0_ext_ram_rdata3[26]
port 242 nsew signal input
rlabel metal2 s 318614 352669 318670 353469 6 data_arrays_0_0_ext_ram_rdata3[27]
port 243 nsew signal input
rlabel metal2 s 319534 352669 319590 353469 6 data_arrays_0_0_ext_ram_rdata3[28]
port 244 nsew signal input
rlabel metal2 s 320362 352669 320418 353469 6 data_arrays_0_0_ext_ram_rdata3[29]
port 245 nsew signal input
rlabel metal2 s 296258 352669 296314 353469 6 data_arrays_0_0_ext_ram_rdata3[2]
port 246 nsew signal input
rlabel metal2 s 321282 352669 321338 353469 6 data_arrays_0_0_ext_ram_rdata3[30]
port 247 nsew signal input
rlabel metal2 s 322202 352669 322258 353469 6 data_arrays_0_0_ext_ram_rdata3[31]
port 248 nsew signal input
rlabel metal2 s 323122 352669 323178 353469 6 data_arrays_0_0_ext_ram_rdata3[32]
port 249 nsew signal input
rlabel metal2 s 323950 352669 324006 353469 6 data_arrays_0_0_ext_ram_rdata3[33]
port 250 nsew signal input
rlabel metal2 s 324870 352669 324926 353469 6 data_arrays_0_0_ext_ram_rdata3[34]
port 251 nsew signal input
rlabel metal2 s 325790 352669 325846 353469 6 data_arrays_0_0_ext_ram_rdata3[35]
port 252 nsew signal input
rlabel metal2 s 326618 352669 326674 353469 6 data_arrays_0_0_ext_ram_rdata3[36]
port 253 nsew signal input
rlabel metal2 s 327538 352669 327594 353469 6 data_arrays_0_0_ext_ram_rdata3[37]
port 254 nsew signal input
rlabel metal2 s 328458 352669 328514 353469 6 data_arrays_0_0_ext_ram_rdata3[38]
port 255 nsew signal input
rlabel metal2 s 329378 352669 329434 353469 6 data_arrays_0_0_ext_ram_rdata3[39]
port 256 nsew signal input
rlabel metal2 s 297178 352669 297234 353469 6 data_arrays_0_0_ext_ram_rdata3[3]
port 257 nsew signal input
rlabel metal2 s 330206 352669 330262 353469 6 data_arrays_0_0_ext_ram_rdata3[40]
port 258 nsew signal input
rlabel metal2 s 331126 352669 331182 353469 6 data_arrays_0_0_ext_ram_rdata3[41]
port 259 nsew signal input
rlabel metal2 s 332046 352669 332102 353469 6 data_arrays_0_0_ext_ram_rdata3[42]
port 260 nsew signal input
rlabel metal2 s 332874 352669 332930 353469 6 data_arrays_0_0_ext_ram_rdata3[43]
port 261 nsew signal input
rlabel metal2 s 333794 352669 333850 353469 6 data_arrays_0_0_ext_ram_rdata3[44]
port 262 nsew signal input
rlabel metal2 s 334714 352669 334770 353469 6 data_arrays_0_0_ext_ram_rdata3[45]
port 263 nsew signal input
rlabel metal2 s 335634 352669 335690 353469 6 data_arrays_0_0_ext_ram_rdata3[46]
port 264 nsew signal input
rlabel metal2 s 336462 352669 336518 353469 6 data_arrays_0_0_ext_ram_rdata3[47]
port 265 nsew signal input
rlabel metal2 s 337382 352669 337438 353469 6 data_arrays_0_0_ext_ram_rdata3[48]
port 266 nsew signal input
rlabel metal2 s 338302 352669 338358 353469 6 data_arrays_0_0_ext_ram_rdata3[49]
port 267 nsew signal input
rlabel metal2 s 298006 352669 298062 353469 6 data_arrays_0_0_ext_ram_rdata3[4]
port 268 nsew signal input
rlabel metal2 s 339130 352669 339186 353469 6 data_arrays_0_0_ext_ram_rdata3[50]
port 269 nsew signal input
rlabel metal2 s 340050 352669 340106 353469 6 data_arrays_0_0_ext_ram_rdata3[51]
port 270 nsew signal input
rlabel metal2 s 340970 352669 341026 353469 6 data_arrays_0_0_ext_ram_rdata3[52]
port 271 nsew signal input
rlabel metal2 s 341890 352669 341946 353469 6 data_arrays_0_0_ext_ram_rdata3[53]
port 272 nsew signal input
rlabel metal2 s 342718 352669 342774 353469 6 data_arrays_0_0_ext_ram_rdata3[54]
port 273 nsew signal input
rlabel metal2 s 343638 352669 343694 353469 6 data_arrays_0_0_ext_ram_rdata3[55]
port 274 nsew signal input
rlabel metal2 s 344558 352669 344614 353469 6 data_arrays_0_0_ext_ram_rdata3[56]
port 275 nsew signal input
rlabel metal2 s 345386 352669 345442 353469 6 data_arrays_0_0_ext_ram_rdata3[57]
port 276 nsew signal input
rlabel metal2 s 346306 352669 346362 353469 6 data_arrays_0_0_ext_ram_rdata3[58]
port 277 nsew signal input
rlabel metal2 s 347226 352669 347282 353469 6 data_arrays_0_0_ext_ram_rdata3[59]
port 278 nsew signal input
rlabel metal2 s 298926 352669 298982 353469 6 data_arrays_0_0_ext_ram_rdata3[5]
port 279 nsew signal input
rlabel metal2 s 348146 352669 348202 353469 6 data_arrays_0_0_ext_ram_rdata3[60]
port 280 nsew signal input
rlabel metal2 s 348974 352669 349030 353469 6 data_arrays_0_0_ext_ram_rdata3[61]
port 281 nsew signal input
rlabel metal2 s 349894 352669 349950 353469 6 data_arrays_0_0_ext_ram_rdata3[62]
port 282 nsew signal input
rlabel metal2 s 350814 352669 350870 353469 6 data_arrays_0_0_ext_ram_rdata3[63]
port 283 nsew signal input
rlabel metal2 s 299846 352669 299902 353469 6 data_arrays_0_0_ext_ram_rdata3[6]
port 284 nsew signal input
rlabel metal2 s 300766 352669 300822 353469 6 data_arrays_0_0_ext_ram_rdata3[7]
port 285 nsew signal input
rlabel metal2 s 301594 352669 301650 353469 6 data_arrays_0_0_ext_ram_rdata3[8]
port 286 nsew signal input
rlabel metal2 s 302514 352669 302570 353469 6 data_arrays_0_0_ext_ram_rdata3[9]
port 287 nsew signal input
rlabel metal3 s 0 216520 800 216640 6 data_arrays_0_0_ext_ram_wdata[0]
port 288 nsew signal output
rlabel metal3 s 0 232160 800 232280 6 data_arrays_0_0_ext_ram_wdata[10]
port 289 nsew signal output
rlabel metal3 s 0 233656 800 233776 6 data_arrays_0_0_ext_ram_wdata[11]
port 290 nsew signal output
rlabel metal3 s 0 235288 800 235408 6 data_arrays_0_0_ext_ram_wdata[12]
port 291 nsew signal output
rlabel metal3 s 0 236784 800 236904 6 data_arrays_0_0_ext_ram_wdata[13]
port 292 nsew signal output
rlabel metal3 s 0 238416 800 238536 6 data_arrays_0_0_ext_ram_wdata[14]
port 293 nsew signal output
rlabel metal3 s 0 239912 800 240032 6 data_arrays_0_0_ext_ram_wdata[15]
port 294 nsew signal output
rlabel metal3 s 0 241544 800 241664 6 data_arrays_0_0_ext_ram_wdata[16]
port 295 nsew signal output
rlabel metal3 s 0 243040 800 243160 6 data_arrays_0_0_ext_ram_wdata[17]
port 296 nsew signal output
rlabel metal3 s 0 244672 800 244792 6 data_arrays_0_0_ext_ram_wdata[18]
port 297 nsew signal output
rlabel metal3 s 0 246168 800 246288 6 data_arrays_0_0_ext_ram_wdata[19]
port 298 nsew signal output
rlabel metal3 s 0 218016 800 218136 6 data_arrays_0_0_ext_ram_wdata[1]
port 299 nsew signal output
rlabel metal3 s 0 247800 800 247920 6 data_arrays_0_0_ext_ram_wdata[20]
port 300 nsew signal output
rlabel metal3 s 0 249296 800 249416 6 data_arrays_0_0_ext_ram_wdata[21]
port 301 nsew signal output
rlabel metal3 s 0 250928 800 251048 6 data_arrays_0_0_ext_ram_wdata[22]
port 302 nsew signal output
rlabel metal3 s 0 252424 800 252544 6 data_arrays_0_0_ext_ram_wdata[23]
port 303 nsew signal output
rlabel metal3 s 0 254056 800 254176 6 data_arrays_0_0_ext_ram_wdata[24]
port 304 nsew signal output
rlabel metal3 s 0 255552 800 255672 6 data_arrays_0_0_ext_ram_wdata[25]
port 305 nsew signal output
rlabel metal3 s 0 257184 800 257304 6 data_arrays_0_0_ext_ram_wdata[26]
port 306 nsew signal output
rlabel metal3 s 0 258680 800 258800 6 data_arrays_0_0_ext_ram_wdata[27]
port 307 nsew signal output
rlabel metal3 s 0 260312 800 260432 6 data_arrays_0_0_ext_ram_wdata[28]
port 308 nsew signal output
rlabel metal3 s 0 261808 800 261928 6 data_arrays_0_0_ext_ram_wdata[29]
port 309 nsew signal output
rlabel metal3 s 0 219648 800 219768 6 data_arrays_0_0_ext_ram_wdata[2]
port 310 nsew signal output
rlabel metal3 s 0 263440 800 263560 6 data_arrays_0_0_ext_ram_wdata[30]
port 311 nsew signal output
rlabel metal3 s 0 264936 800 265056 6 data_arrays_0_0_ext_ram_wdata[31]
port 312 nsew signal output
rlabel metal3 s 0 266568 800 266688 6 data_arrays_0_0_ext_ram_wdata[32]
port 313 nsew signal output
rlabel metal3 s 0 268064 800 268184 6 data_arrays_0_0_ext_ram_wdata[33]
port 314 nsew signal output
rlabel metal3 s 0 269696 800 269816 6 data_arrays_0_0_ext_ram_wdata[34]
port 315 nsew signal output
rlabel metal3 s 0 271192 800 271312 6 data_arrays_0_0_ext_ram_wdata[35]
port 316 nsew signal output
rlabel metal3 s 0 272824 800 272944 6 data_arrays_0_0_ext_ram_wdata[36]
port 317 nsew signal output
rlabel metal3 s 0 274320 800 274440 6 data_arrays_0_0_ext_ram_wdata[37]
port 318 nsew signal output
rlabel metal3 s 0 275952 800 276072 6 data_arrays_0_0_ext_ram_wdata[38]
port 319 nsew signal output
rlabel metal3 s 0 277448 800 277568 6 data_arrays_0_0_ext_ram_wdata[39]
port 320 nsew signal output
rlabel metal3 s 0 221144 800 221264 6 data_arrays_0_0_ext_ram_wdata[3]
port 321 nsew signal output
rlabel metal3 s 0 279080 800 279200 6 data_arrays_0_0_ext_ram_wdata[40]
port 322 nsew signal output
rlabel metal3 s 0 280576 800 280696 6 data_arrays_0_0_ext_ram_wdata[41]
port 323 nsew signal output
rlabel metal3 s 0 282208 800 282328 6 data_arrays_0_0_ext_ram_wdata[42]
port 324 nsew signal output
rlabel metal3 s 0 283704 800 283824 6 data_arrays_0_0_ext_ram_wdata[43]
port 325 nsew signal output
rlabel metal3 s 0 285336 800 285456 6 data_arrays_0_0_ext_ram_wdata[44]
port 326 nsew signal output
rlabel metal3 s 0 286832 800 286952 6 data_arrays_0_0_ext_ram_wdata[45]
port 327 nsew signal output
rlabel metal3 s 0 288464 800 288584 6 data_arrays_0_0_ext_ram_wdata[46]
port 328 nsew signal output
rlabel metal3 s 0 289960 800 290080 6 data_arrays_0_0_ext_ram_wdata[47]
port 329 nsew signal output
rlabel metal3 s 0 291592 800 291712 6 data_arrays_0_0_ext_ram_wdata[48]
port 330 nsew signal output
rlabel metal3 s 0 293088 800 293208 6 data_arrays_0_0_ext_ram_wdata[49]
port 331 nsew signal output
rlabel metal3 s 0 222776 800 222896 6 data_arrays_0_0_ext_ram_wdata[4]
port 332 nsew signal output
rlabel metal3 s 0 294720 800 294840 6 data_arrays_0_0_ext_ram_wdata[50]
port 333 nsew signal output
rlabel metal3 s 0 296216 800 296336 6 data_arrays_0_0_ext_ram_wdata[51]
port 334 nsew signal output
rlabel metal3 s 0 297848 800 297968 6 data_arrays_0_0_ext_ram_wdata[52]
port 335 nsew signal output
rlabel metal3 s 0 299344 800 299464 6 data_arrays_0_0_ext_ram_wdata[53]
port 336 nsew signal output
rlabel metal3 s 0 300976 800 301096 6 data_arrays_0_0_ext_ram_wdata[54]
port 337 nsew signal output
rlabel metal3 s 0 302472 800 302592 6 data_arrays_0_0_ext_ram_wdata[55]
port 338 nsew signal output
rlabel metal3 s 0 304104 800 304224 6 data_arrays_0_0_ext_ram_wdata[56]
port 339 nsew signal output
rlabel metal3 s 0 305600 800 305720 6 data_arrays_0_0_ext_ram_wdata[57]
port 340 nsew signal output
rlabel metal3 s 0 307232 800 307352 6 data_arrays_0_0_ext_ram_wdata[58]
port 341 nsew signal output
rlabel metal3 s 0 308728 800 308848 6 data_arrays_0_0_ext_ram_wdata[59]
port 342 nsew signal output
rlabel metal3 s 0 224272 800 224392 6 data_arrays_0_0_ext_ram_wdata[5]
port 343 nsew signal output
rlabel metal3 s 0 310360 800 310480 6 data_arrays_0_0_ext_ram_wdata[60]
port 344 nsew signal output
rlabel metal3 s 0 311856 800 311976 6 data_arrays_0_0_ext_ram_wdata[61]
port 345 nsew signal output
rlabel metal3 s 0 313488 800 313608 6 data_arrays_0_0_ext_ram_wdata[62]
port 346 nsew signal output
rlabel metal3 s 0 314984 800 315104 6 data_arrays_0_0_ext_ram_wdata[63]
port 347 nsew signal output
rlabel metal3 s 0 225904 800 226024 6 data_arrays_0_0_ext_ram_wdata[6]
port 348 nsew signal output
rlabel metal3 s 0 227400 800 227520 6 data_arrays_0_0_ext_ram_wdata[7]
port 349 nsew signal output
rlabel metal3 s 0 229032 800 229152 6 data_arrays_0_0_ext_ram_wdata[8]
port 350 nsew signal output
rlabel metal3 s 0 230528 800 230648 6 data_arrays_0_0_ext_ram_wdata[9]
port 351 nsew signal output
rlabel metal3 s 0 326000 800 326120 6 data_arrays_0_0_ext_ram_web
port 352 nsew signal output
rlabel metal3 s 0 316616 800 316736 6 data_arrays_0_0_ext_ram_wmask[0]
port 353 nsew signal output
rlabel metal3 s 0 318112 800 318232 6 data_arrays_0_0_ext_ram_wmask[1]
port 354 nsew signal output
rlabel metal2 s 135350 352669 135406 353469 6 io_in[0]
port 355 nsew signal input
rlabel metal2 s 162122 352669 162178 353469 6 io_in[10]
port 356 nsew signal input
rlabel metal2 s 164882 352669 164938 353469 6 io_in[11]
port 357 nsew signal input
rlabel metal2 s 167550 352669 167606 353469 6 io_in[12]
port 358 nsew signal input
rlabel metal2 s 170218 352669 170274 353469 6 io_in[13]
port 359 nsew signal input
rlabel metal2 s 172886 352669 172942 353469 6 io_in[14]
port 360 nsew signal input
rlabel metal2 s 175554 352669 175610 353469 6 io_in[15]
port 361 nsew signal input
rlabel metal2 s 178222 352669 178278 353469 6 io_in[16]
port 362 nsew signal input
rlabel metal2 s 180890 352669 180946 353469 6 io_in[17]
port 363 nsew signal input
rlabel metal2 s 183650 352669 183706 353469 6 io_in[18]
port 364 nsew signal input
rlabel metal2 s 186318 352669 186374 353469 6 io_in[19]
port 365 nsew signal input
rlabel metal2 s 138018 352669 138074 353469 6 io_in[1]
port 366 nsew signal input
rlabel metal2 s 188986 352669 189042 353469 6 io_in[20]
port 367 nsew signal input
rlabel metal2 s 191654 352669 191710 353469 6 io_in[21]
port 368 nsew signal input
rlabel metal2 s 194322 352669 194378 353469 6 io_in[22]
port 369 nsew signal input
rlabel metal2 s 196990 352669 197046 353469 6 io_in[23]
port 370 nsew signal input
rlabel metal2 s 199750 352669 199806 353469 6 io_in[24]
port 371 nsew signal input
rlabel metal2 s 202418 352669 202474 353469 6 io_in[25]
port 372 nsew signal input
rlabel metal2 s 205086 352669 205142 353469 6 io_in[26]
port 373 nsew signal input
rlabel metal2 s 207754 352669 207810 353469 6 io_in[27]
port 374 nsew signal input
rlabel metal2 s 210422 352669 210478 353469 6 io_in[28]
port 375 nsew signal input
rlabel metal2 s 213090 352669 213146 353469 6 io_in[29]
port 376 nsew signal input
rlabel metal2 s 140686 352669 140742 353469 6 io_in[2]
port 377 nsew signal input
rlabel metal2 s 215758 352669 215814 353469 6 io_in[30]
port 378 nsew signal input
rlabel metal2 s 218518 352669 218574 353469 6 io_in[31]
port 379 nsew signal input
rlabel metal2 s 221186 352669 221242 353469 6 io_in[32]
port 380 nsew signal input
rlabel metal2 s 223854 352669 223910 353469 6 io_in[33]
port 381 nsew signal input
rlabel metal2 s 226522 352669 226578 353469 6 io_in[34]
port 382 nsew signal input
rlabel metal2 s 229190 352669 229246 353469 6 io_in[35]
port 383 nsew signal input
rlabel metal2 s 231858 352669 231914 353469 6 io_in[36]
port 384 nsew signal input
rlabel metal2 s 234618 352669 234674 353469 6 io_in[37]
port 385 nsew signal input
rlabel metal2 s 143354 352669 143410 353469 6 io_in[3]
port 386 nsew signal input
rlabel metal2 s 146022 352669 146078 353469 6 io_in[4]
port 387 nsew signal input
rlabel metal2 s 148782 352669 148838 353469 6 io_in[5]
port 388 nsew signal input
rlabel metal2 s 151450 352669 151506 353469 6 io_in[6]
port 389 nsew signal input
rlabel metal2 s 154118 352669 154174 353469 6 io_in[7]
port 390 nsew signal input
rlabel metal2 s 156786 352669 156842 353469 6 io_in[8]
port 391 nsew signal input
rlabel metal2 s 159454 352669 159510 353469 6 io_in[9]
port 392 nsew signal input
rlabel metal2 s 136270 352669 136326 353469 6 io_oeb[0]
port 393 nsew signal output
rlabel metal2 s 163042 352669 163098 353469 6 io_oeb[10]
port 394 nsew signal output
rlabel metal2 s 165710 352669 165766 353469 6 io_oeb[11]
port 395 nsew signal output
rlabel metal2 s 168378 352669 168434 353469 6 io_oeb[12]
port 396 nsew signal output
rlabel metal2 s 171138 352669 171194 353469 6 io_oeb[13]
port 397 nsew signal output
rlabel metal2 s 173806 352669 173862 353469 6 io_oeb[14]
port 398 nsew signal output
rlabel metal2 s 176474 352669 176530 353469 6 io_oeb[15]
port 399 nsew signal output
rlabel metal2 s 179142 352669 179198 353469 6 io_oeb[16]
port 400 nsew signal output
rlabel metal2 s 181810 352669 181866 353469 6 io_oeb[17]
port 401 nsew signal output
rlabel metal2 s 184478 352669 184534 353469 6 io_oeb[18]
port 402 nsew signal output
rlabel metal2 s 187146 352669 187202 353469 6 io_oeb[19]
port 403 nsew signal output
rlabel metal2 s 138938 352669 138994 353469 6 io_oeb[1]
port 404 nsew signal output
rlabel metal2 s 189906 352669 189962 353469 6 io_oeb[20]
port 405 nsew signal output
rlabel metal2 s 192574 352669 192630 353469 6 io_oeb[21]
port 406 nsew signal output
rlabel metal2 s 195242 352669 195298 353469 6 io_oeb[22]
port 407 nsew signal output
rlabel metal2 s 197910 352669 197966 353469 6 io_oeb[23]
port 408 nsew signal output
rlabel metal2 s 200578 352669 200634 353469 6 io_oeb[24]
port 409 nsew signal output
rlabel metal2 s 203246 352669 203302 353469 6 io_oeb[25]
port 410 nsew signal output
rlabel metal2 s 206006 352669 206062 353469 6 io_oeb[26]
port 411 nsew signal output
rlabel metal2 s 208674 352669 208730 353469 6 io_oeb[27]
port 412 nsew signal output
rlabel metal2 s 211342 352669 211398 353469 6 io_oeb[28]
port 413 nsew signal output
rlabel metal2 s 214010 352669 214066 353469 6 io_oeb[29]
port 414 nsew signal output
rlabel metal2 s 141606 352669 141662 353469 6 io_oeb[2]
port 415 nsew signal output
rlabel metal2 s 216678 352669 216734 353469 6 io_oeb[30]
port 416 nsew signal output
rlabel metal2 s 219346 352669 219402 353469 6 io_oeb[31]
port 417 nsew signal output
rlabel metal2 s 222014 352669 222070 353469 6 io_oeb[32]
port 418 nsew signal output
rlabel metal2 s 224774 352669 224830 353469 6 io_oeb[33]
port 419 nsew signal output
rlabel metal2 s 227442 352669 227498 353469 6 io_oeb[34]
port 420 nsew signal output
rlabel metal2 s 230110 352669 230166 353469 6 io_oeb[35]
port 421 nsew signal output
rlabel metal2 s 232778 352669 232834 353469 6 io_oeb[36]
port 422 nsew signal output
rlabel metal2 s 235446 352669 235502 353469 6 io_oeb[37]
port 423 nsew signal output
rlabel metal2 s 144274 352669 144330 353469 6 io_oeb[3]
port 424 nsew signal output
rlabel metal2 s 146942 352669 146998 353469 6 io_oeb[4]
port 425 nsew signal output
rlabel metal2 s 149610 352669 149666 353469 6 io_oeb[5]
port 426 nsew signal output
rlabel metal2 s 152278 352669 152334 353469 6 io_oeb[6]
port 427 nsew signal output
rlabel metal2 s 155038 352669 155094 353469 6 io_oeb[7]
port 428 nsew signal output
rlabel metal2 s 157706 352669 157762 353469 6 io_oeb[8]
port 429 nsew signal output
rlabel metal2 s 160374 352669 160430 353469 6 io_oeb[9]
port 430 nsew signal output
rlabel metal2 s 137098 352669 137154 353469 6 io_out[0]
port 431 nsew signal output
rlabel metal2 s 163962 352669 164018 353469 6 io_out[10]
port 432 nsew signal output
rlabel metal2 s 166630 352669 166686 353469 6 io_out[11]
port 433 nsew signal output
rlabel metal2 s 169298 352669 169354 353469 6 io_out[12]
port 434 nsew signal output
rlabel metal2 s 171966 352669 172022 353469 6 io_out[13]
port 435 nsew signal output
rlabel metal2 s 174634 352669 174690 353469 6 io_out[14]
port 436 nsew signal output
rlabel metal2 s 177394 352669 177450 353469 6 io_out[15]
port 437 nsew signal output
rlabel metal2 s 180062 352669 180118 353469 6 io_out[16]
port 438 nsew signal output
rlabel metal2 s 182730 352669 182786 353469 6 io_out[17]
port 439 nsew signal output
rlabel metal2 s 185398 352669 185454 353469 6 io_out[18]
port 440 nsew signal output
rlabel metal2 s 188066 352669 188122 353469 6 io_out[19]
port 441 nsew signal output
rlabel metal2 s 139766 352669 139822 353469 6 io_out[1]
port 442 nsew signal output
rlabel metal2 s 190734 352669 190790 353469 6 io_out[20]
port 443 nsew signal output
rlabel metal2 s 193402 352669 193458 353469 6 io_out[21]
port 444 nsew signal output
rlabel metal2 s 196162 352669 196218 353469 6 io_out[22]
port 445 nsew signal output
rlabel metal2 s 198830 352669 198886 353469 6 io_out[23]
port 446 nsew signal output
rlabel metal2 s 201498 352669 201554 353469 6 io_out[24]
port 447 nsew signal output
rlabel metal2 s 204166 352669 204222 353469 6 io_out[25]
port 448 nsew signal output
rlabel metal2 s 206834 352669 206890 353469 6 io_out[26]
port 449 nsew signal output
rlabel metal2 s 209502 352669 209558 353469 6 io_out[27]
port 450 nsew signal output
rlabel metal2 s 212262 352669 212318 353469 6 io_out[28]
port 451 nsew signal output
rlabel metal2 s 214930 352669 214986 353469 6 io_out[29]
port 452 nsew signal output
rlabel metal2 s 142526 352669 142582 353469 6 io_out[2]
port 453 nsew signal output
rlabel metal2 s 217598 352669 217654 353469 6 io_out[30]
port 454 nsew signal output
rlabel metal2 s 220266 352669 220322 353469 6 io_out[31]
port 455 nsew signal output
rlabel metal2 s 222934 352669 222990 353469 6 io_out[32]
port 456 nsew signal output
rlabel metal2 s 225602 352669 225658 353469 6 io_out[33]
port 457 nsew signal output
rlabel metal2 s 228270 352669 228326 353469 6 io_out[34]
port 458 nsew signal output
rlabel metal2 s 231030 352669 231086 353469 6 io_out[35]
port 459 nsew signal output
rlabel metal2 s 233698 352669 233754 353469 6 io_out[36]
port 460 nsew signal output
rlabel metal2 s 236366 352669 236422 353469 6 io_out[37]
port 461 nsew signal output
rlabel metal2 s 145194 352669 145250 353469 6 io_out[3]
port 462 nsew signal output
rlabel metal2 s 147862 352669 147918 353469 6 io_out[4]
port 463 nsew signal output
rlabel metal2 s 150530 352669 150586 353469 6 io_out[5]
port 464 nsew signal output
rlabel metal2 s 153198 352669 153254 353469 6 io_out[6]
port 465 nsew signal output
rlabel metal2 s 155866 352669 155922 353469 6 io_out[7]
port 466 nsew signal output
rlabel metal2 s 158626 352669 158682 353469 6 io_out[8]
port 467 nsew signal output
rlabel metal2 s 161294 352669 161350 353469 6 io_out[9]
port 468 nsew signal output
rlabel metal2 s 349434 0 349490 800 6 irq[0]
port 469 nsew signal output
rlabel metal2 s 350170 0 350226 800 6 irq[1]
port 470 nsew signal output
rlabel metal2 s 350906 0 350962 800 6 irq[2]
port 471 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 la_data_in[0]
port 472 nsew signal input
rlabel metal2 s 289634 0 289690 800 6 la_data_in[100]
port 473 nsew signal input
rlabel metal2 s 291750 0 291806 800 6 la_data_in[101]
port 474 nsew signal input
rlabel metal2 s 293866 0 293922 800 6 la_data_in[102]
port 475 nsew signal input
rlabel metal2 s 295982 0 296038 800 6 la_data_in[103]
port 476 nsew signal input
rlabel metal2 s 298190 0 298246 800 6 la_data_in[104]
port 477 nsew signal input
rlabel metal2 s 300306 0 300362 800 6 la_data_in[105]
port 478 nsew signal input
rlabel metal2 s 302422 0 302478 800 6 la_data_in[106]
port 479 nsew signal input
rlabel metal2 s 304538 0 304594 800 6 la_data_in[107]
port 480 nsew signal input
rlabel metal2 s 306654 0 306710 800 6 la_data_in[108]
port 481 nsew signal input
rlabel metal2 s 308862 0 308918 800 6 la_data_in[109]
port 482 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_data_in[10]
port 483 nsew signal input
rlabel metal2 s 310978 0 311034 800 6 la_data_in[110]
port 484 nsew signal input
rlabel metal2 s 313094 0 313150 800 6 la_data_in[111]
port 485 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_data_in[112]
port 486 nsew signal input
rlabel metal2 s 317418 0 317474 800 6 la_data_in[113]
port 487 nsew signal input
rlabel metal2 s 319534 0 319590 800 6 la_data_in[114]
port 488 nsew signal input
rlabel metal2 s 321650 0 321706 800 6 la_data_in[115]
port 489 nsew signal input
rlabel metal2 s 323766 0 323822 800 6 la_data_in[116]
port 490 nsew signal input
rlabel metal2 s 325974 0 326030 800 6 la_data_in[117]
port 491 nsew signal input
rlabel metal2 s 328090 0 328146 800 6 la_data_in[118]
port 492 nsew signal input
rlabel metal2 s 330206 0 330262 800 6 la_data_in[119]
port 493 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[11]
port 494 nsew signal input
rlabel metal2 s 332322 0 332378 800 6 la_data_in[120]
port 495 nsew signal input
rlabel metal2 s 334530 0 334586 800 6 la_data_in[121]
port 496 nsew signal input
rlabel metal2 s 336646 0 336702 800 6 la_data_in[122]
port 497 nsew signal input
rlabel metal2 s 338762 0 338818 800 6 la_data_in[123]
port 498 nsew signal input
rlabel metal2 s 340878 0 340934 800 6 la_data_in[124]
port 499 nsew signal input
rlabel metal2 s 343086 0 343142 800 6 la_data_in[125]
port 500 nsew signal input
rlabel metal2 s 345202 0 345258 800 6 la_data_in[126]
port 501 nsew signal input
rlabel metal2 s 347318 0 347374 800 6 la_data_in[127]
port 502 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[12]
port 503 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[13]
port 504 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_data_in[14]
port 505 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[15]
port 506 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[16]
port 507 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_data_in[17]
port 508 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[18]
port 509 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[19]
port 510 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[1]
port 511 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[20]
port 512 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_data_in[21]
port 513 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[22]
port 514 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[23]
port 515 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_data_in[24]
port 516 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[25]
port 517 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[26]
port 518 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[27]
port 519 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_data_in[28]
port 520 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_data_in[29]
port 521 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[2]
port 522 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[30]
port 523 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_data_in[31]
port 524 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[32]
port 525 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[33]
port 526 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_data_in[34]
port 527 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_data_in[35]
port 528 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[36]
port 529 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_data_in[37]
port 530 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_data_in[38]
port 531 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_data_in[39]
port 532 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[3]
port 533 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_data_in[40]
port 534 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[41]
port 535 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_data_in[42]
port 536 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_data_in[43]
port 537 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_data_in[44]
port 538 nsew signal input
rlabel metal2 s 171966 0 172022 800 6 la_data_in[45]
port 539 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_data_in[46]
port 540 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 la_data_in[47]
port 541 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_data_in[48]
port 542 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_data_in[49]
port 543 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[4]
port 544 nsew signal input
rlabel metal2 s 182730 0 182786 800 6 la_data_in[50]
port 545 nsew signal input
rlabel metal2 s 184846 0 184902 800 6 la_data_in[51]
port 546 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_data_in[52]
port 547 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_data_in[53]
port 548 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 la_data_in[54]
port 549 nsew signal input
rlabel metal2 s 193402 0 193458 800 6 la_data_in[55]
port 550 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 la_data_in[56]
port 551 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_data_in[57]
port 552 nsew signal input
rlabel metal2 s 199842 0 199898 800 6 la_data_in[58]
port 553 nsew signal input
rlabel metal2 s 201958 0 202014 800 6 la_data_in[59]
port 554 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_data_in[5]
port 555 nsew signal input
rlabel metal2 s 204074 0 204130 800 6 la_data_in[60]
port 556 nsew signal input
rlabel metal2 s 206190 0 206246 800 6 la_data_in[61]
port 557 nsew signal input
rlabel metal2 s 208306 0 208362 800 6 la_data_in[62]
port 558 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_data_in[63]
port 559 nsew signal input
rlabel metal2 s 212630 0 212686 800 6 la_data_in[64]
port 560 nsew signal input
rlabel metal2 s 214746 0 214802 800 6 la_data_in[65]
port 561 nsew signal input
rlabel metal2 s 216862 0 216918 800 6 la_data_in[66]
port 562 nsew signal input
rlabel metal2 s 219070 0 219126 800 6 la_data_in[67]
port 563 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_data_in[68]
port 564 nsew signal input
rlabel metal2 s 223302 0 223358 800 6 la_data_in[69]
port 565 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[6]
port 566 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_data_in[70]
port 567 nsew signal input
rlabel metal2 s 227626 0 227682 800 6 la_data_in[71]
port 568 nsew signal input
rlabel metal2 s 229742 0 229798 800 6 la_data_in[72]
port 569 nsew signal input
rlabel metal2 s 231858 0 231914 800 6 la_data_in[73]
port 570 nsew signal input
rlabel metal2 s 233974 0 234030 800 6 la_data_in[74]
port 571 nsew signal input
rlabel metal2 s 236182 0 236238 800 6 la_data_in[75]
port 572 nsew signal input
rlabel metal2 s 238298 0 238354 800 6 la_data_in[76]
port 573 nsew signal input
rlabel metal2 s 240414 0 240470 800 6 la_data_in[77]
port 574 nsew signal input
rlabel metal2 s 242530 0 242586 800 6 la_data_in[78]
port 575 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 la_data_in[79]
port 576 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[7]
port 577 nsew signal input
rlabel metal2 s 246854 0 246910 800 6 la_data_in[80]
port 578 nsew signal input
rlabel metal2 s 248970 0 249026 800 6 la_data_in[81]
port 579 nsew signal input
rlabel metal2 s 251086 0 251142 800 6 la_data_in[82]
port 580 nsew signal input
rlabel metal2 s 253202 0 253258 800 6 la_data_in[83]
port 581 nsew signal input
rlabel metal2 s 255410 0 255466 800 6 la_data_in[84]
port 582 nsew signal input
rlabel metal2 s 257526 0 257582 800 6 la_data_in[85]
port 583 nsew signal input
rlabel metal2 s 259642 0 259698 800 6 la_data_in[86]
port 584 nsew signal input
rlabel metal2 s 261758 0 261814 800 6 la_data_in[87]
port 585 nsew signal input
rlabel metal2 s 263966 0 264022 800 6 la_data_in[88]
port 586 nsew signal input
rlabel metal2 s 266082 0 266138 800 6 la_data_in[89]
port 587 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[8]
port 588 nsew signal input
rlabel metal2 s 268198 0 268254 800 6 la_data_in[90]
port 589 nsew signal input
rlabel metal2 s 270314 0 270370 800 6 la_data_in[91]
port 590 nsew signal input
rlabel metal2 s 272522 0 272578 800 6 la_data_in[92]
port 591 nsew signal input
rlabel metal2 s 274638 0 274694 800 6 la_data_in[93]
port 592 nsew signal input
rlabel metal2 s 276754 0 276810 800 6 la_data_in[94]
port 593 nsew signal input
rlabel metal2 s 278870 0 278926 800 6 la_data_in[95]
port 594 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_data_in[96]
port 595 nsew signal input
rlabel metal2 s 283194 0 283250 800 6 la_data_in[97]
port 596 nsew signal input
rlabel metal2 s 285310 0 285366 800 6 la_data_in[98]
port 597 nsew signal input
rlabel metal2 s 287426 0 287482 800 6 la_data_in[99]
port 598 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_data_in[9]
port 599 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_out[0]
port 600 nsew signal output
rlabel metal2 s 290278 0 290334 800 6 la_data_out[100]
port 601 nsew signal output
rlabel metal2 s 292486 0 292542 800 6 la_data_out[101]
port 602 nsew signal output
rlabel metal2 s 294602 0 294658 800 6 la_data_out[102]
port 603 nsew signal output
rlabel metal2 s 296718 0 296774 800 6 la_data_out[103]
port 604 nsew signal output
rlabel metal2 s 298834 0 298890 800 6 la_data_out[104]
port 605 nsew signal output
rlabel metal2 s 301042 0 301098 800 6 la_data_out[105]
port 606 nsew signal output
rlabel metal2 s 303158 0 303214 800 6 la_data_out[106]
port 607 nsew signal output
rlabel metal2 s 305274 0 305330 800 6 la_data_out[107]
port 608 nsew signal output
rlabel metal2 s 307390 0 307446 800 6 la_data_out[108]
port 609 nsew signal output
rlabel metal2 s 309506 0 309562 800 6 la_data_out[109]
port 610 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[10]
port 611 nsew signal output
rlabel metal2 s 311714 0 311770 800 6 la_data_out[110]
port 612 nsew signal output
rlabel metal2 s 313830 0 313886 800 6 la_data_out[111]
port 613 nsew signal output
rlabel metal2 s 315946 0 316002 800 6 la_data_out[112]
port 614 nsew signal output
rlabel metal2 s 318062 0 318118 800 6 la_data_out[113]
port 615 nsew signal output
rlabel metal2 s 320270 0 320326 800 6 la_data_out[114]
port 616 nsew signal output
rlabel metal2 s 322386 0 322442 800 6 la_data_out[115]
port 617 nsew signal output
rlabel metal2 s 324502 0 324558 800 6 la_data_out[116]
port 618 nsew signal output
rlabel metal2 s 326618 0 326674 800 6 la_data_out[117]
port 619 nsew signal output
rlabel metal2 s 328826 0 328882 800 6 la_data_out[118]
port 620 nsew signal output
rlabel metal2 s 330942 0 330998 800 6 la_data_out[119]
port 621 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[11]
port 622 nsew signal output
rlabel metal2 s 333058 0 333114 800 6 la_data_out[120]
port 623 nsew signal output
rlabel metal2 s 335174 0 335230 800 6 la_data_out[121]
port 624 nsew signal output
rlabel metal2 s 337382 0 337438 800 6 la_data_out[122]
port 625 nsew signal output
rlabel metal2 s 339498 0 339554 800 6 la_data_out[123]
port 626 nsew signal output
rlabel metal2 s 341614 0 341670 800 6 la_data_out[124]
port 627 nsew signal output
rlabel metal2 s 343730 0 343786 800 6 la_data_out[125]
port 628 nsew signal output
rlabel metal2 s 345938 0 345994 800 6 la_data_out[126]
port 629 nsew signal output
rlabel metal2 s 348054 0 348110 800 6 la_data_out[127]
port 630 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[12]
port 631 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[13]
port 632 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 la_data_out[14]
port 633 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[15]
port 634 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[16]
port 635 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[17]
port 636 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 la_data_out[18]
port 637 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 la_data_out[19]
port 638 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[1]
port 639 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 la_data_out[20]
port 640 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[21]
port 641 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[22]
port 642 nsew signal output
rlabel metal2 s 125690 0 125746 800 6 la_data_out[23]
port 643 nsew signal output
rlabel metal2 s 127806 0 127862 800 6 la_data_out[24]
port 644 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 la_data_out[25]
port 645 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[26]
port 646 nsew signal output
rlabel metal2 s 134246 0 134302 800 6 la_data_out[27]
port 647 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[28]
port 648 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 la_data_out[29]
port 649 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[2]
port 650 nsew signal output
rlabel metal2 s 140686 0 140742 800 6 la_data_out[30]
port 651 nsew signal output
rlabel metal2 s 142802 0 142858 800 6 la_data_out[31]
port 652 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[32]
port 653 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[33]
port 654 nsew signal output
rlabel metal2 s 149242 0 149298 800 6 la_data_out[34]
port 655 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 la_data_out[35]
port 656 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 la_data_out[36]
port 657 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[37]
port 658 nsew signal output
rlabel metal2 s 157706 0 157762 800 6 la_data_out[38]
port 659 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 la_data_out[39]
port 660 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[3]
port 661 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 la_data_out[40]
port 662 nsew signal output
rlabel metal2 s 164146 0 164202 800 6 la_data_out[41]
port 663 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 la_data_out[42]
port 664 nsew signal output
rlabel metal2 s 168470 0 168526 800 6 la_data_out[43]
port 665 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 la_data_out[44]
port 666 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 la_data_out[45]
port 667 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[46]
port 668 nsew signal output
rlabel metal2 s 177026 0 177082 800 6 la_data_out[47]
port 669 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 la_data_out[48]
port 670 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 la_data_out[49]
port 671 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[4]
port 672 nsew signal output
rlabel metal2 s 183374 0 183430 800 6 la_data_out[50]
port 673 nsew signal output
rlabel metal2 s 185582 0 185638 800 6 la_data_out[51]
port 674 nsew signal output
rlabel metal2 s 187698 0 187754 800 6 la_data_out[52]
port 675 nsew signal output
rlabel metal2 s 189814 0 189870 800 6 la_data_out[53]
port 676 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 la_data_out[54]
port 677 nsew signal output
rlabel metal2 s 194138 0 194194 800 6 la_data_out[55]
port 678 nsew signal output
rlabel metal2 s 196254 0 196310 800 6 la_data_out[56]
port 679 nsew signal output
rlabel metal2 s 198370 0 198426 800 6 la_data_out[57]
port 680 nsew signal output
rlabel metal2 s 200486 0 200542 800 6 la_data_out[58]
port 681 nsew signal output
rlabel metal2 s 202602 0 202658 800 6 la_data_out[59]
port 682 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[5]
port 683 nsew signal output
rlabel metal2 s 204810 0 204866 800 6 la_data_out[60]
port 684 nsew signal output
rlabel metal2 s 206926 0 206982 800 6 la_data_out[61]
port 685 nsew signal output
rlabel metal2 s 209042 0 209098 800 6 la_data_out[62]
port 686 nsew signal output
rlabel metal2 s 211158 0 211214 800 6 la_data_out[63]
port 687 nsew signal output
rlabel metal2 s 213366 0 213422 800 6 la_data_out[64]
port 688 nsew signal output
rlabel metal2 s 215482 0 215538 800 6 la_data_out[65]
port 689 nsew signal output
rlabel metal2 s 217598 0 217654 800 6 la_data_out[66]
port 690 nsew signal output
rlabel metal2 s 219714 0 219770 800 6 la_data_out[67]
port 691 nsew signal output
rlabel metal2 s 221922 0 221978 800 6 la_data_out[68]
port 692 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 la_data_out[69]
port 693 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[6]
port 694 nsew signal output
rlabel metal2 s 226154 0 226210 800 6 la_data_out[70]
port 695 nsew signal output
rlabel metal2 s 228270 0 228326 800 6 la_data_out[71]
port 696 nsew signal output
rlabel metal2 s 230478 0 230534 800 6 la_data_out[72]
port 697 nsew signal output
rlabel metal2 s 232594 0 232650 800 6 la_data_out[73]
port 698 nsew signal output
rlabel metal2 s 234710 0 234766 800 6 la_data_out[74]
port 699 nsew signal output
rlabel metal2 s 236826 0 236882 800 6 la_data_out[75]
port 700 nsew signal output
rlabel metal2 s 239034 0 239090 800 6 la_data_out[76]
port 701 nsew signal output
rlabel metal2 s 241150 0 241206 800 6 la_data_out[77]
port 702 nsew signal output
rlabel metal2 s 243266 0 243322 800 6 la_data_out[78]
port 703 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 la_data_out[79]
port 704 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[7]
port 705 nsew signal output
rlabel metal2 s 247590 0 247646 800 6 la_data_out[80]
port 706 nsew signal output
rlabel metal2 s 249706 0 249762 800 6 la_data_out[81]
port 707 nsew signal output
rlabel metal2 s 251822 0 251878 800 6 la_data_out[82]
port 708 nsew signal output
rlabel metal2 s 253938 0 253994 800 6 la_data_out[83]
port 709 nsew signal output
rlabel metal2 s 256054 0 256110 800 6 la_data_out[84]
port 710 nsew signal output
rlabel metal2 s 258262 0 258318 800 6 la_data_out[85]
port 711 nsew signal output
rlabel metal2 s 260378 0 260434 800 6 la_data_out[86]
port 712 nsew signal output
rlabel metal2 s 262494 0 262550 800 6 la_data_out[87]
port 713 nsew signal output
rlabel metal2 s 264610 0 264666 800 6 la_data_out[88]
port 714 nsew signal output
rlabel metal2 s 266818 0 266874 800 6 la_data_out[89]
port 715 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[8]
port 716 nsew signal output
rlabel metal2 s 268934 0 268990 800 6 la_data_out[90]
port 717 nsew signal output
rlabel metal2 s 271050 0 271106 800 6 la_data_out[91]
port 718 nsew signal output
rlabel metal2 s 273166 0 273222 800 6 la_data_out[92]
port 719 nsew signal output
rlabel metal2 s 275374 0 275430 800 6 la_data_out[93]
port 720 nsew signal output
rlabel metal2 s 277490 0 277546 800 6 la_data_out[94]
port 721 nsew signal output
rlabel metal2 s 279606 0 279662 800 6 la_data_out[95]
port 722 nsew signal output
rlabel metal2 s 281722 0 281778 800 6 la_data_out[96]
port 723 nsew signal output
rlabel metal2 s 283930 0 283986 800 6 la_data_out[97]
port 724 nsew signal output
rlabel metal2 s 286046 0 286102 800 6 la_data_out[98]
port 725 nsew signal output
rlabel metal2 s 288162 0 288218 800 6 la_data_out[99]
port 726 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[9]
port 727 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 la_oenb[0]
port 728 nsew signal input
rlabel metal2 s 291014 0 291070 800 6 la_oenb[100]
port 729 nsew signal input
rlabel metal2 s 293130 0 293186 800 6 la_oenb[101]
port 730 nsew signal input
rlabel metal2 s 295338 0 295394 800 6 la_oenb[102]
port 731 nsew signal input
rlabel metal2 s 297454 0 297510 800 6 la_oenb[103]
port 732 nsew signal input
rlabel metal2 s 299570 0 299626 800 6 la_oenb[104]
port 733 nsew signal input
rlabel metal2 s 301686 0 301742 800 6 la_oenb[105]
port 734 nsew signal input
rlabel metal2 s 303802 0 303858 800 6 la_oenb[106]
port 735 nsew signal input
rlabel metal2 s 306010 0 306066 800 6 la_oenb[107]
port 736 nsew signal input
rlabel metal2 s 308126 0 308182 800 6 la_oenb[108]
port 737 nsew signal input
rlabel metal2 s 310242 0 310298 800 6 la_oenb[109]
port 738 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[10]
port 739 nsew signal input
rlabel metal2 s 312358 0 312414 800 6 la_oenb[110]
port 740 nsew signal input
rlabel metal2 s 314566 0 314622 800 6 la_oenb[111]
port 741 nsew signal input
rlabel metal2 s 316682 0 316738 800 6 la_oenb[112]
port 742 nsew signal input
rlabel metal2 s 318798 0 318854 800 6 la_oenb[113]
port 743 nsew signal input
rlabel metal2 s 320914 0 320970 800 6 la_oenb[114]
port 744 nsew signal input
rlabel metal2 s 323122 0 323178 800 6 la_oenb[115]
port 745 nsew signal input
rlabel metal2 s 325238 0 325294 800 6 la_oenb[116]
port 746 nsew signal input
rlabel metal2 s 327354 0 327410 800 6 la_oenb[117]
port 747 nsew signal input
rlabel metal2 s 329470 0 329526 800 6 la_oenb[118]
port 748 nsew signal input
rlabel metal2 s 331678 0 331734 800 6 la_oenb[119]
port 749 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[11]
port 750 nsew signal input
rlabel metal2 s 333794 0 333850 800 6 la_oenb[120]
port 751 nsew signal input
rlabel metal2 s 335910 0 335966 800 6 la_oenb[121]
port 752 nsew signal input
rlabel metal2 s 338026 0 338082 800 6 la_oenb[122]
port 753 nsew signal input
rlabel metal2 s 340234 0 340290 800 6 la_oenb[123]
port 754 nsew signal input
rlabel metal2 s 342350 0 342406 800 6 la_oenb[124]
port 755 nsew signal input
rlabel metal2 s 344466 0 344522 800 6 la_oenb[125]
port 756 nsew signal input
rlabel metal2 s 346582 0 346638 800 6 la_oenb[126]
port 757 nsew signal input
rlabel metal2 s 348790 0 348846 800 6 la_oenb[127]
port 758 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[12]
port 759 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[13]
port 760 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_oenb[14]
port 761 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_oenb[15]
port 762 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[16]
port 763 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_oenb[17]
port 764 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[18]
port 765 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[19]
port 766 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[1]
port 767 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_oenb[20]
port 768 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_oenb[21]
port 769 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_oenb[22]
port 770 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_oenb[23]
port 771 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oenb[24]
port 772 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_oenb[25]
port 773 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_oenb[26]
port 774 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 la_oenb[27]
port 775 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oenb[28]
port 776 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oenb[29]
port 777 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_oenb[2]
port 778 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[30]
port 779 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_oenb[31]
port 780 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_oenb[32]
port 781 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oenb[33]
port 782 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_oenb[34]
port 783 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_oenb[35]
port 784 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_oenb[36]
port 785 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_oenb[37]
port 786 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oenb[38]
port 787 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oenb[39]
port 788 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[3]
port 789 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[40]
port 790 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_oenb[41]
port 791 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_oenb[42]
port 792 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_oenb[43]
port 793 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_oenb[44]
port 794 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 la_oenb[45]
port 795 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_oenb[46]
port 796 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oenb[47]
port 797 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 la_oenb[48]
port 798 nsew signal input
rlabel metal2 s 181994 0 182050 800 6 la_oenb[49]
port 799 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[4]
port 800 nsew signal input
rlabel metal2 s 184110 0 184166 800 6 la_oenb[50]
port 801 nsew signal input
rlabel metal2 s 186226 0 186282 800 6 la_oenb[51]
port 802 nsew signal input
rlabel metal2 s 188434 0 188490 800 6 la_oenb[52]
port 803 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_oenb[53]
port 804 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 la_oenb[54]
port 805 nsew signal input
rlabel metal2 s 194782 0 194838 800 6 la_oenb[55]
port 806 nsew signal input
rlabel metal2 s 196990 0 197046 800 6 la_oenb[56]
port 807 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_oenb[57]
port 808 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_oenb[58]
port 809 nsew signal input
rlabel metal2 s 203338 0 203394 800 6 la_oenb[59]
port 810 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[5]
port 811 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_oenb[60]
port 812 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_oenb[61]
port 813 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_oenb[62]
port 814 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 la_oenb[63]
port 815 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 la_oenb[64]
port 816 nsew signal input
rlabel metal2 s 216218 0 216274 800 6 la_oenb[65]
port 817 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 la_oenb[66]
port 818 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_oenb[67]
port 819 nsew signal input
rlabel metal2 s 222566 0 222622 800 6 la_oenb[68]
port 820 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_oenb[69]
port 821 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[6]
port 822 nsew signal input
rlabel metal2 s 226890 0 226946 800 6 la_oenb[70]
port 823 nsew signal input
rlabel metal2 s 229006 0 229062 800 6 la_oenb[71]
port 824 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_oenb[72]
port 825 nsew signal input
rlabel metal2 s 233330 0 233386 800 6 la_oenb[73]
port 826 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_oenb[74]
port 827 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_oenb[75]
port 828 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_oenb[76]
port 829 nsew signal input
rlabel metal2 s 241886 0 241942 800 6 la_oenb[77]
port 830 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 la_oenb[78]
port 831 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 la_oenb[79]
port 832 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[7]
port 833 nsew signal input
rlabel metal2 s 248234 0 248290 800 6 la_oenb[80]
port 834 nsew signal input
rlabel metal2 s 250442 0 250498 800 6 la_oenb[81]
port 835 nsew signal input
rlabel metal2 s 252558 0 252614 800 6 la_oenb[82]
port 836 nsew signal input
rlabel metal2 s 254674 0 254730 800 6 la_oenb[83]
port 837 nsew signal input
rlabel metal2 s 256790 0 256846 800 6 la_oenb[84]
port 838 nsew signal input
rlabel metal2 s 258906 0 258962 800 6 la_oenb[85]
port 839 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_oenb[86]
port 840 nsew signal input
rlabel metal2 s 263230 0 263286 800 6 la_oenb[87]
port 841 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 la_oenb[88]
port 842 nsew signal input
rlabel metal2 s 267462 0 267518 800 6 la_oenb[89]
port 843 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_oenb[8]
port 844 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 la_oenb[90]
port 845 nsew signal input
rlabel metal2 s 271786 0 271842 800 6 la_oenb[91]
port 846 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 la_oenb[92]
port 847 nsew signal input
rlabel metal2 s 276018 0 276074 800 6 la_oenb[93]
port 848 nsew signal input
rlabel metal2 s 278226 0 278282 800 6 la_oenb[94]
port 849 nsew signal input
rlabel metal2 s 280342 0 280398 800 6 la_oenb[95]
port 850 nsew signal input
rlabel metal2 s 282458 0 282514 800 6 la_oenb[96]
port 851 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 la_oenb[97]
port 852 nsew signal input
rlabel metal2 s 286782 0 286838 800 6 la_oenb[98]
port 853 nsew signal input
rlabel metal2 s 288898 0 288954 800 6 la_oenb[99]
port 854 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[9]
port 855 nsew signal input
rlabel metal2 s 99562 352669 99618 353469 6 tag_array_ext_ram_addr1[0]
port 856 nsew signal output
rlabel metal2 s 100482 352669 100538 353469 6 tag_array_ext_ram_addr1[1]
port 857 nsew signal output
rlabel metal2 s 101402 352669 101458 353469 6 tag_array_ext_ram_addr1[2]
port 858 nsew signal output
rlabel metal2 s 102230 352669 102286 353469 6 tag_array_ext_ram_addr1[3]
port 859 nsew signal output
rlabel metal2 s 103150 352669 103206 353469 6 tag_array_ext_ram_addr1[4]
port 860 nsew signal output
rlabel metal2 s 104070 352669 104126 353469 6 tag_array_ext_ram_addr1[5]
port 861 nsew signal output
rlabel metal2 s 104898 352669 104954 353469 6 tag_array_ext_ram_addr1[6]
port 862 nsew signal output
rlabel metal2 s 105818 352669 105874 353469 6 tag_array_ext_ram_addr1[7]
port 863 nsew signal output
rlabel metal2 s 28906 352669 28962 353469 6 tag_array_ext_ram_addr[0]
port 864 nsew signal output
rlabel metal2 s 29826 352669 29882 353469 6 tag_array_ext_ram_addr[1]
port 865 nsew signal output
rlabel metal2 s 30746 352669 30802 353469 6 tag_array_ext_ram_addr[2]
port 866 nsew signal output
rlabel metal2 s 31666 352669 31722 353469 6 tag_array_ext_ram_addr[3]
port 867 nsew signal output
rlabel metal2 s 32494 352669 32550 353469 6 tag_array_ext_ram_addr[4]
port 868 nsew signal output
rlabel metal2 s 33414 352669 33470 353469 6 tag_array_ext_ram_addr[5]
port 869 nsew signal output
rlabel metal2 s 34334 352669 34390 353469 6 tag_array_ext_ram_addr[6]
port 870 nsew signal output
rlabel metal2 s 35162 352669 35218 353469 6 tag_array_ext_ram_addr[7]
port 871 nsew signal output
rlabel metal2 s 36082 352669 36138 353469 6 tag_array_ext_ram_clk
port 872 nsew signal output
rlabel metal2 s 95974 352669 96030 353469 6 tag_array_ext_ram_csb
port 873 nsew signal output
rlabel metal2 s 97814 352669 97870 353469 6 tag_array_ext_ram_csb1[0]
port 874 nsew signal output
rlabel metal2 s 98642 352669 98698 353469 6 tag_array_ext_ram_csb1[1]
port 875 nsew signal output
rlabel metal2 s 386 352669 442 353469 6 tag_array_ext_ram_rdata0[0]
port 876 nsew signal input
rlabel metal2 s 9310 352669 9366 353469 6 tag_array_ext_ram_rdata0[10]
port 877 nsew signal input
rlabel metal2 s 10138 352669 10194 353469 6 tag_array_ext_ram_rdata0[11]
port 878 nsew signal input
rlabel metal2 s 11058 352669 11114 353469 6 tag_array_ext_ram_rdata0[12]
port 879 nsew signal input
rlabel metal2 s 11978 352669 12034 353469 6 tag_array_ext_ram_rdata0[13]
port 880 nsew signal input
rlabel metal2 s 12898 352669 12954 353469 6 tag_array_ext_ram_rdata0[14]
port 881 nsew signal input
rlabel metal2 s 13726 352669 13782 353469 6 tag_array_ext_ram_rdata0[15]
port 882 nsew signal input
rlabel metal2 s 14646 352669 14702 353469 6 tag_array_ext_ram_rdata0[16]
port 883 nsew signal input
rlabel metal2 s 15566 352669 15622 353469 6 tag_array_ext_ram_rdata0[17]
port 884 nsew signal input
rlabel metal2 s 16394 352669 16450 353469 6 tag_array_ext_ram_rdata0[18]
port 885 nsew signal input
rlabel metal2 s 17314 352669 17370 353469 6 tag_array_ext_ram_rdata0[19]
port 886 nsew signal input
rlabel metal2 s 1214 352669 1270 353469 6 tag_array_ext_ram_rdata0[1]
port 887 nsew signal input
rlabel metal2 s 18234 352669 18290 353469 6 tag_array_ext_ram_rdata0[20]
port 888 nsew signal input
rlabel metal2 s 19154 352669 19210 353469 6 tag_array_ext_ram_rdata0[21]
port 889 nsew signal input
rlabel metal2 s 19982 352669 20038 353469 6 tag_array_ext_ram_rdata0[22]
port 890 nsew signal input
rlabel metal2 s 20902 352669 20958 353469 6 tag_array_ext_ram_rdata0[23]
port 891 nsew signal input
rlabel metal2 s 21822 352669 21878 353469 6 tag_array_ext_ram_rdata0[24]
port 892 nsew signal input
rlabel metal2 s 22650 352669 22706 353469 6 tag_array_ext_ram_rdata0[25]
port 893 nsew signal input
rlabel metal2 s 23570 352669 23626 353469 6 tag_array_ext_ram_rdata0[26]
port 894 nsew signal input
rlabel metal2 s 24490 352669 24546 353469 6 tag_array_ext_ram_rdata0[27]
port 895 nsew signal input
rlabel metal2 s 25410 352669 25466 353469 6 tag_array_ext_ram_rdata0[28]
port 896 nsew signal input
rlabel metal2 s 26238 352669 26294 353469 6 tag_array_ext_ram_rdata0[29]
port 897 nsew signal input
rlabel metal2 s 2134 352669 2190 353469 6 tag_array_ext_ram_rdata0[2]
port 898 nsew signal input
rlabel metal2 s 27158 352669 27214 353469 6 tag_array_ext_ram_rdata0[30]
port 899 nsew signal input
rlabel metal2 s 28078 352669 28134 353469 6 tag_array_ext_ram_rdata0[31]
port 900 nsew signal input
rlabel metal2 s 3054 352669 3110 353469 6 tag_array_ext_ram_rdata0[3]
port 901 nsew signal input
rlabel metal2 s 3882 352669 3938 353469 6 tag_array_ext_ram_rdata0[4]
port 902 nsew signal input
rlabel metal2 s 4802 352669 4858 353469 6 tag_array_ext_ram_rdata0[5]
port 903 nsew signal input
rlabel metal2 s 5722 352669 5778 353469 6 tag_array_ext_ram_rdata0[6]
port 904 nsew signal input
rlabel metal2 s 6642 352669 6698 353469 6 tag_array_ext_ram_rdata0[7]
port 905 nsew signal input
rlabel metal2 s 7470 352669 7526 353469 6 tag_array_ext_ram_rdata0[8]
port 906 nsew signal input
rlabel metal2 s 8390 352669 8446 353469 6 tag_array_ext_ram_rdata0[9]
port 907 nsew signal input
rlabel metal2 s 106738 352669 106794 353469 6 tag_array_ext_ram_rdata1[0]
port 908 nsew signal input
rlabel metal2 s 115662 352669 115718 353469 6 tag_array_ext_ram_rdata1[10]
port 909 nsew signal input
rlabel metal2 s 116582 352669 116638 353469 6 tag_array_ext_ram_rdata1[11]
port 910 nsew signal input
rlabel metal2 s 117502 352669 117558 353469 6 tag_array_ext_ram_rdata1[12]
port 911 nsew signal input
rlabel metal2 s 118330 352669 118386 353469 6 tag_array_ext_ram_rdata1[13]
port 912 nsew signal input
rlabel metal2 s 119250 352669 119306 353469 6 tag_array_ext_ram_rdata1[14]
port 913 nsew signal input
rlabel metal2 s 120170 352669 120226 353469 6 tag_array_ext_ram_rdata1[15]
port 914 nsew signal input
rlabel metal2 s 120998 352669 121054 353469 6 tag_array_ext_ram_rdata1[16]
port 915 nsew signal input
rlabel metal2 s 121918 352669 121974 353469 6 tag_array_ext_ram_rdata1[17]
port 916 nsew signal input
rlabel metal2 s 122838 352669 122894 353469 6 tag_array_ext_ram_rdata1[18]
port 917 nsew signal input
rlabel metal2 s 123758 352669 123814 353469 6 tag_array_ext_ram_rdata1[19]
port 918 nsew signal input
rlabel metal2 s 107658 352669 107714 353469 6 tag_array_ext_ram_rdata1[1]
port 919 nsew signal input
rlabel metal2 s 124586 352669 124642 353469 6 tag_array_ext_ram_rdata1[20]
port 920 nsew signal input
rlabel metal2 s 125506 352669 125562 353469 6 tag_array_ext_ram_rdata1[21]
port 921 nsew signal input
rlabel metal2 s 126426 352669 126482 353469 6 tag_array_ext_ram_rdata1[22]
port 922 nsew signal input
rlabel metal2 s 127254 352669 127310 353469 6 tag_array_ext_ram_rdata1[23]
port 923 nsew signal input
rlabel metal2 s 128174 352669 128230 353469 6 tag_array_ext_ram_rdata1[24]
port 924 nsew signal input
rlabel metal2 s 129094 352669 129150 353469 6 tag_array_ext_ram_rdata1[25]
port 925 nsew signal input
rlabel metal2 s 130014 352669 130070 353469 6 tag_array_ext_ram_rdata1[26]
port 926 nsew signal input
rlabel metal2 s 130842 352669 130898 353469 6 tag_array_ext_ram_rdata1[27]
port 927 nsew signal input
rlabel metal2 s 131762 352669 131818 353469 6 tag_array_ext_ram_rdata1[28]
port 928 nsew signal input
rlabel metal2 s 132682 352669 132738 353469 6 tag_array_ext_ram_rdata1[29]
port 929 nsew signal input
rlabel metal2 s 108486 352669 108542 353469 6 tag_array_ext_ram_rdata1[2]
port 930 nsew signal input
rlabel metal2 s 133510 352669 133566 353469 6 tag_array_ext_ram_rdata1[30]
port 931 nsew signal input
rlabel metal2 s 134430 352669 134486 353469 6 tag_array_ext_ram_rdata1[31]
port 932 nsew signal input
rlabel metal2 s 109406 352669 109462 353469 6 tag_array_ext_ram_rdata1[3]
port 933 nsew signal input
rlabel metal2 s 110326 352669 110382 353469 6 tag_array_ext_ram_rdata1[4]
port 934 nsew signal input
rlabel metal2 s 111154 352669 111210 353469 6 tag_array_ext_ram_rdata1[5]
port 935 nsew signal input
rlabel metal2 s 112074 352669 112130 353469 6 tag_array_ext_ram_rdata1[6]
port 936 nsew signal input
rlabel metal2 s 112994 352669 113050 353469 6 tag_array_ext_ram_rdata1[7]
port 937 nsew signal input
rlabel metal2 s 113914 352669 113970 353469 6 tag_array_ext_ram_rdata1[8]
port 938 nsew signal input
rlabel metal2 s 114742 352669 114798 353469 6 tag_array_ext_ram_rdata1[9]
port 939 nsew signal input
rlabel metal2 s 37002 352669 37058 353469 6 tag_array_ext_ram_wdata[0]
port 940 nsew signal output
rlabel metal2 s 45926 352669 45982 353469 6 tag_array_ext_ram_wdata[10]
port 941 nsew signal output
rlabel metal2 s 46846 352669 46902 353469 6 tag_array_ext_ram_wdata[11]
port 942 nsew signal output
rlabel metal2 s 47766 352669 47822 353469 6 tag_array_ext_ram_wdata[12]
port 943 nsew signal output
rlabel metal2 s 48594 352669 48650 353469 6 tag_array_ext_ram_wdata[13]
port 944 nsew signal output
rlabel metal2 s 49514 352669 49570 353469 6 tag_array_ext_ram_wdata[14]
port 945 nsew signal output
rlabel metal2 s 50434 352669 50490 353469 6 tag_array_ext_ram_wdata[15]
port 946 nsew signal output
rlabel metal2 s 51262 352669 51318 353469 6 tag_array_ext_ram_wdata[16]
port 947 nsew signal output
rlabel metal2 s 52182 352669 52238 353469 6 tag_array_ext_ram_wdata[17]
port 948 nsew signal output
rlabel metal2 s 53102 352669 53158 353469 6 tag_array_ext_ram_wdata[18]
port 949 nsew signal output
rlabel metal2 s 54022 352669 54078 353469 6 tag_array_ext_ram_wdata[19]
port 950 nsew signal output
rlabel metal2 s 37922 352669 37978 353469 6 tag_array_ext_ram_wdata[1]
port 951 nsew signal output
rlabel metal2 s 54850 352669 54906 353469 6 tag_array_ext_ram_wdata[20]
port 952 nsew signal output
rlabel metal2 s 55770 352669 55826 353469 6 tag_array_ext_ram_wdata[21]
port 953 nsew signal output
rlabel metal2 s 56690 352669 56746 353469 6 tag_array_ext_ram_wdata[22]
port 954 nsew signal output
rlabel metal2 s 57518 352669 57574 353469 6 tag_array_ext_ram_wdata[23]
port 955 nsew signal output
rlabel metal2 s 58438 352669 58494 353469 6 tag_array_ext_ram_wdata[24]
port 956 nsew signal output
rlabel metal2 s 59358 352669 59414 353469 6 tag_array_ext_ram_wdata[25]
port 957 nsew signal output
rlabel metal2 s 60278 352669 60334 353469 6 tag_array_ext_ram_wdata[26]
port 958 nsew signal output
rlabel metal2 s 61106 352669 61162 353469 6 tag_array_ext_ram_wdata[27]
port 959 nsew signal output
rlabel metal2 s 62026 352669 62082 353469 6 tag_array_ext_ram_wdata[28]
port 960 nsew signal output
rlabel metal2 s 62946 352669 63002 353469 6 tag_array_ext_ram_wdata[29]
port 961 nsew signal output
rlabel metal2 s 38750 352669 38806 353469 6 tag_array_ext_ram_wdata[2]
port 962 nsew signal output
rlabel metal2 s 63774 352669 63830 353469 6 tag_array_ext_ram_wdata[30]
port 963 nsew signal output
rlabel metal2 s 64694 352669 64750 353469 6 tag_array_ext_ram_wdata[31]
port 964 nsew signal output
rlabel metal2 s 65614 352669 65670 353469 6 tag_array_ext_ram_wdata[32]
port 965 nsew signal output
rlabel metal2 s 66534 352669 66590 353469 6 tag_array_ext_ram_wdata[33]
port 966 nsew signal output
rlabel metal2 s 67362 352669 67418 353469 6 tag_array_ext_ram_wdata[34]
port 967 nsew signal output
rlabel metal2 s 68282 352669 68338 353469 6 tag_array_ext_ram_wdata[35]
port 968 nsew signal output
rlabel metal2 s 69202 352669 69258 353469 6 tag_array_ext_ram_wdata[36]
port 969 nsew signal output
rlabel metal2 s 70030 352669 70086 353469 6 tag_array_ext_ram_wdata[37]
port 970 nsew signal output
rlabel metal2 s 70950 352669 71006 353469 6 tag_array_ext_ram_wdata[38]
port 971 nsew signal output
rlabel metal2 s 71870 352669 71926 353469 6 tag_array_ext_ram_wdata[39]
port 972 nsew signal output
rlabel metal2 s 39670 352669 39726 353469 6 tag_array_ext_ram_wdata[3]
port 973 nsew signal output
rlabel metal2 s 72790 352669 72846 353469 6 tag_array_ext_ram_wdata[40]
port 974 nsew signal output
rlabel metal2 s 73618 352669 73674 353469 6 tag_array_ext_ram_wdata[41]
port 975 nsew signal output
rlabel metal2 s 74538 352669 74594 353469 6 tag_array_ext_ram_wdata[42]
port 976 nsew signal output
rlabel metal2 s 75458 352669 75514 353469 6 tag_array_ext_ram_wdata[43]
port 977 nsew signal output
rlabel metal2 s 76286 352669 76342 353469 6 tag_array_ext_ram_wdata[44]
port 978 nsew signal output
rlabel metal2 s 77206 352669 77262 353469 6 tag_array_ext_ram_wdata[45]
port 979 nsew signal output
rlabel metal2 s 78126 352669 78182 353469 6 tag_array_ext_ram_wdata[46]
port 980 nsew signal output
rlabel metal2 s 79046 352669 79102 353469 6 tag_array_ext_ram_wdata[47]
port 981 nsew signal output
rlabel metal2 s 79874 352669 79930 353469 6 tag_array_ext_ram_wdata[48]
port 982 nsew signal output
rlabel metal2 s 80794 352669 80850 353469 6 tag_array_ext_ram_wdata[49]
port 983 nsew signal output
rlabel metal2 s 40590 352669 40646 353469 6 tag_array_ext_ram_wdata[4]
port 984 nsew signal output
rlabel metal2 s 81714 352669 81770 353469 6 tag_array_ext_ram_wdata[50]
port 985 nsew signal output
rlabel metal2 s 82634 352669 82690 353469 6 tag_array_ext_ram_wdata[51]
port 986 nsew signal output
rlabel metal2 s 83462 352669 83518 353469 6 tag_array_ext_ram_wdata[52]
port 987 nsew signal output
rlabel metal2 s 84382 352669 84438 353469 6 tag_array_ext_ram_wdata[53]
port 988 nsew signal output
rlabel metal2 s 85302 352669 85358 353469 6 tag_array_ext_ram_wdata[54]
port 989 nsew signal output
rlabel metal2 s 86130 352669 86186 353469 6 tag_array_ext_ram_wdata[55]
port 990 nsew signal output
rlabel metal2 s 87050 352669 87106 353469 6 tag_array_ext_ram_wdata[56]
port 991 nsew signal output
rlabel metal2 s 87970 352669 88026 353469 6 tag_array_ext_ram_wdata[57]
port 992 nsew signal output
rlabel metal2 s 88890 352669 88946 353469 6 tag_array_ext_ram_wdata[58]
port 993 nsew signal output
rlabel metal2 s 89718 352669 89774 353469 6 tag_array_ext_ram_wdata[59]
port 994 nsew signal output
rlabel metal2 s 41510 352669 41566 353469 6 tag_array_ext_ram_wdata[5]
port 995 nsew signal output
rlabel metal2 s 90638 352669 90694 353469 6 tag_array_ext_ram_wdata[60]
port 996 nsew signal output
rlabel metal2 s 91558 352669 91614 353469 6 tag_array_ext_ram_wdata[61]
port 997 nsew signal output
rlabel metal2 s 92386 352669 92442 353469 6 tag_array_ext_ram_wdata[62]
port 998 nsew signal output
rlabel metal2 s 93306 352669 93362 353469 6 tag_array_ext_ram_wdata[63]
port 999 nsew signal output
rlabel metal2 s 42338 352669 42394 353469 6 tag_array_ext_ram_wdata[6]
port 1000 nsew signal output
rlabel metal2 s 43258 352669 43314 353469 6 tag_array_ext_ram_wdata[7]
port 1001 nsew signal output
rlabel metal2 s 44178 352669 44234 353469 6 tag_array_ext_ram_wdata[8]
port 1002 nsew signal output
rlabel metal2 s 45006 352669 45062 353469 6 tag_array_ext_ram_wdata[9]
port 1003 nsew signal output
rlabel metal2 s 96894 352669 96950 353469 6 tag_array_ext_ram_web
port 1004 nsew signal output
rlabel metal2 s 94226 352669 94282 353469 6 tag_array_ext_ram_wmask[0]
port 1005 nsew signal output
rlabel metal2 s 95146 352669 95202 353469 6 tag_array_ext_ram_wmask[1]
port 1006 nsew signal output
rlabel metal4 s 4208 2128 4528 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 34928 2128 35248 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 65648 2128 65968 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 96368 2128 96688 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 127088 2128 127408 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 157808 2128 158128 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 188528 2128 188848 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 219248 2128 219568 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 249968 2128 250288 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 280688 2128 281008 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 311408 2128 311728 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 342128 2128 342448 350928 6 vccd1
port 1007 nsew power input
rlabel metal4 s 19568 2128 19888 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 50288 2128 50608 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 81008 2128 81328 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 111728 2128 112048 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 142448 2128 142768 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 173168 2128 173488 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 203888 2128 204208 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 234608 2128 234928 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 265328 2128 265648 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 296048 2128 296368 350928 6 vssd1
port 1008 nsew ground input
rlabel metal4 s 326768 2128 327088 350928 6 vssd1
port 1008 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 1009 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 1010 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_ack_o
port 1011 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[0]
port 1012 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[10]
port 1013 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[11]
port 1014 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[12]
port 1015 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_adr_i[13]
port 1016 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[14]
port 1017 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[15]
port 1018 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_adr_i[16]
port 1019 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[17]
port 1020 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_adr_i[18]
port 1021 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_adr_i[19]
port 1022 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[1]
port 1023 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[20]
port 1024 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 wbs_adr_i[21]
port 1025 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_adr_i[22]
port 1026 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_adr_i[23]
port 1027 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_adr_i[24]
port 1028 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_adr_i[25]
port 1029 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 wbs_adr_i[26]
port 1030 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_adr_i[27]
port 1031 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 wbs_adr_i[28]
port 1032 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 wbs_adr_i[29]
port 1033 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[2]
port 1034 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 wbs_adr_i[30]
port 1035 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 wbs_adr_i[31]
port 1036 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[3]
port 1037 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[4]
port 1038 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[5]
port 1039 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[6]
port 1040 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_adr_i[7]
port 1041 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[8]
port 1042 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_adr_i[9]
port 1043 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_cyc_i
port 1044 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_i[0]
port 1045 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[10]
port 1046 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[11]
port 1047 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[12]
port 1048 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_i[13]
port 1049 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[14]
port 1050 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[15]
port 1051 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 wbs_dat_i[16]
port 1052 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_dat_i[17]
port 1053 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_i[18]
port 1054 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_dat_i[19]
port 1055 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[1]
port 1056 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[20]
port 1057 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_i[21]
port 1058 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[22]
port 1059 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_i[23]
port 1060 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 wbs_dat_i[24]
port 1061 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_dat_i[25]
port 1062 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 wbs_dat_i[26]
port 1063 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_i[27]
port 1064 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 wbs_dat_i[28]
port 1065 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 wbs_dat_i[29]
port 1066 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[2]
port 1067 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 wbs_dat_i[30]
port 1068 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 wbs_dat_i[31]
port 1069 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[3]
port 1070 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[4]
port 1071 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[5]
port 1072 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_i[6]
port 1073 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[7]
port 1074 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[8]
port 1075 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_i[9]
port 1076 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[0]
port 1077 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_o[10]
port 1078 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[11]
port 1079 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[12]
port 1080 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_o[13]
port 1081 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_o[14]
port 1082 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[15]
port 1083 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[16]
port 1084 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_o[17]
port 1085 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_o[18]
port 1086 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_o[19]
port 1087 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[1]
port 1088 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_o[20]
port 1089 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 wbs_dat_o[21]
port 1090 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 wbs_dat_o[22]
port 1091 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_o[23]
port 1092 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_o[24]
port 1093 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 wbs_dat_o[25]
port 1094 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 wbs_dat_o[26]
port 1095 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 wbs_dat_o[27]
port 1096 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 wbs_dat_o[28]
port 1097 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 wbs_dat_o[29]
port 1098 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[2]
port 1099 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 wbs_dat_o[30]
port 1100 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 wbs_dat_o[31]
port 1101 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[3]
port 1102 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[4]
port 1103 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[5]
port 1104 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[6]
port 1105 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_o[7]
port 1106 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[8]
port 1107 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_o[9]
port 1108 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_sel_i[0]
port 1109 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_sel_i[1]
port 1110 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_sel_i[2]
port 1111 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_sel_i[3]
port 1112 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_stb_i
port 1113 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_we_i
port 1114 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 351325 353469
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 299386342
string GDS_FILE /home/shc/Development/efabless/marmot_asic/openlane/marmot/runs/marmot/results/finishing/Marmot.magic.gds
string GDS_START 1973466
<< end >>

